module fake_netlist_6_3082_n_14691 (n_992, n_2542, n_1671, n_1, n_2817, n_801, n_1613, n_1234, n_1458, n_2576, n_3254, n_1199, n_1674, n_3392, n_741, n_1027, n_1351, n_3266, n_625, n_1189, n_3152, n_223, n_1212, n_226, n_208, n_68, n_726, n_2157, n_3335, n_2332, n_212, n_700, n_50, n_1307, n_3178, n_2003, n_1038, n_578, n_1581, n_1003, n_365, n_168, n_1237, n_1061, n_2353, n_2534, n_3089, n_3301, n_1357, n_1853, n_77, n_783, n_2451, n_1738, n_2243, n_798, n_188, n_1575, n_1854, n_2324, n_3088, n_3443, n_1923, n_3257, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_2260, n_3222, n_677, n_1708, n_805, n_1151, n_396, n_2977, n_1739, n_350, n_78, n_2051, n_2317, n_1380, n_2359, n_442, n_480, n_142, n_2847, n_1402, n_2557, n_1688, n_1691, n_3332, n_3465, n_1975, n_1009, n_1743, n_62, n_1930, n_2405, n_1160, n_883, n_2647, n_1238, n_1991, n_2570, n_2179, n_2386, n_2997, n_1724, n_1032, n_2336, n_1247, n_1547, n_2521, n_3376, n_3046, n_2956, n_1553, n_893, n_1099, n_2491, n_1264, n_1192, n_471, n_1844, n_424, n_1700, n_1555, n_1415, n_2211, n_1370, n_1786, n_369, n_287, n_2382, n_2672, n_3030, n_2291, n_415, n_830, n_2299, n_65, n_230, n_3340, n_461, n_873, n_141, n_383, n_1285, n_1371, n_2886, n_2974, n_200, n_1985, n_2989, n_447, n_2838, n_2184, n_3395, n_2982, n_1803, n_3427, n_1172, n_852, n_2509, n_71, n_229, n_2513, n_3282, n_1590, n_2645, n_1532, n_2313, n_2628, n_3071, n_1393, n_1517, n_1867, n_2926, n_1704, n_1078, n_250, n_544, n_1711, n_2247, n_3106, n_1140, n_2630, n_1444, n_1670, n_1603, n_2344, n_1579, n_3275, n_35, n_2365, n_2470, n_2321, n_1263, n_2019, n_3031, n_836, n_3345, n_375, n_2074, n_2447, n_522, n_2919, n_3440, n_2129, n_2340, n_1261, n_945, n_2286, n_1649, n_2018, n_2094, n_3080, n_1903, n_1511, n_1143, n_2356, n_2399, n_1422, n_1232, n_1772, n_1572, n_616, n_658, n_1874, n_3165, n_1119, n_2865, n_2825, n_3463, n_2013, n_428, n_1433, n_1902, n_1842, n_1620, n_2044, n_1954, n_1735, n_2510, n_1541, n_1300, n_641, n_2480, n_2739, n_3023, n_822, n_3232, n_693, n_1313, n_2791, n_3251, n_1056, n_3316, n_2212, n_758, n_516, n_3048, n_1455, n_2418, n_2864, n_1163, n_2729, n_3063, n_1180, n_2256, n_2582, n_943, n_1798, n_1550, n_2703, n_491, n_2786, n_3371, n_1591, n_42, n_772, n_3122, n_2806, n_1344, n_3261, n_2730, n_2495, n_666, n_371, n_940, n_770, n_567, n_1781, n_1971, n_2058, n_2090, n_2603, n_405, n_213, n_2660, n_538, n_3028, n_2981, n_3076, n_2173, n_2004, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_3077, n_1345, n_1820, n_2873, n_3452, n_494, n_539, n_493, n_3107, n_155, n_2880, n_3225, n_2394, n_2108, n_45, n_454, n_1421, n_2836, n_1936, n_638, n_1404, n_1211, n_2124, n_381, n_2378, n_887, n_1660, n_1961, n_3047, n_112, n_1280, n_713, n_2655, n_1400, n_2625, n_3296, n_2843, n_126, n_1467, n_3297, n_58, n_976, n_3067, n_2155, n_224, n_2686, n_48, n_1445, n_2364, n_2551, n_1526, n_1560, n_734, n_1088, n_1894, n_196, n_1231, n_2996, n_2599, n_2985, n_1978, n_2085, n_3368, n_917, n_574, n_9, n_3347, n_2370, n_2612, n_907, n_6, n_1446, n_14, n_2591, n_659, n_1815, n_2214, n_3351, n_407, n_913, n_1658, n_2593, n_808, n_867, n_3269, n_1230, n_3413, n_473, n_1193, n_1967, n_1054, n_559, n_3412, n_2613, n_1333, n_2496, n_44, n_2708, n_3313, n_1648, n_3189, n_1911, n_1956, n_163, n_1644, n_2011, n_2725, n_2277, n_3164, n_1558, n_1732, n_281, n_551, n_699, n_1986, n_2300, n_564, n_2397, n_451, n_824, n_279, n_686, n_757, n_594, n_1641, n_2113, n_1918, n_2190, n_2907, n_577, n_3438, n_166, n_2735, n_1843, n_619, n_2268, n_1367, n_1336, n_521, n_2778, n_2850, n_572, n_395, n_813, n_1909, n_2080, n_1481, n_323, n_606, n_1441, n_818, n_3373, n_1123, n_1309, n_92, n_2104, n_513, n_645, n_1381, n_2961, n_331, n_1699, n_916, n_2093, n_2633, n_483, n_102, n_2207, n_1970, n_2770, n_608, n_261, n_2101, n_2696, n_630, n_2059, n_32, n_2198, n_3319, n_541, n_512, n_2669, n_2925, n_2073, n_2273, n_121, n_433, n_2546, n_3272, n_3193, n_792, n_2522, n_476, n_2792, n_2, n_1328, n_3396, n_1957, n_2917, n_219, n_2616, n_3118, n_3315, n_1907, n_2529, n_264, n_263, n_1162, n_860, n_1530, n_788, n_939, n_1543, n_821, n_2811, n_938, n_1302, n_1068, n_1599, n_329, n_982, n_2674, n_2832, n_549, n_1762, n_1910, n_1075, n_408, n_932, n_2831, n_2998, n_3446, n_61, n_3317, n_237, n_1876, n_1895, n_2123, n_1697, n_2143, n_243, n_979, n_1873, n_905, n_1866, n_1680, n_117, n_175, n_322, n_993, n_2692, n_689, n_3248, n_2031, n_354, n_2130, n_1330, n_1413, n_1605, n_2228, n_3397, n_134, n_1988, n_2941, n_1278, n_547, n_2455, n_2876, n_558, n_2654, n_3036, n_2469, n_1064, n_3099, n_1396, n_634, n_2355, n_136, n_966, n_2908, n_3168, n_764, n_2751, n_2764, n_3357, n_1663, n_2895, n_2009, n_692, n_3403, n_733, n_1793, n_2922, n_1233, n_1289, n_2714, n_2245, n_487, n_3055, n_3092, n_241, n_30, n_2068, n_1107, n_2866, n_2457, n_3294, n_1014, n_1290, n_1703, n_2580, n_3455, n_882, n_2176, n_2072, n_1354, n_2821, n_586, n_423, n_1865, n_1875, n_1701, n_2459, n_318, n_1111, n_1713, n_2971, n_715, n_2678, n_1251, n_3384, n_1265, n_2711, n_88, n_1726, n_1950, n_530, n_1563, n_1912, n_277, n_2434, n_3369, n_3419, n_1982, n_2878, n_618, n_3012, n_1297, n_1662, n_1312, n_199, n_1167, n_1359, n_2818, n_2428, n_674, n_3247, n_871, n_3069, n_922, n_268, n_1335, n_1760, n_1927, n_210, n_2028, n_1069, n_2664, n_5, n_1664, n_1722, n_612, n_2641, n_3022, n_3052, n_178, n_247, n_1165, n_355, n_702, n_347, n_2008, n_2749, n_3298, n_2192, n_3281, n_2254, n_2345, n_3346, n_1926, n_1175, n_3273, n_328, n_1386, n_2311, n_1896, n_429, n_2965, n_1747, n_3058, n_1012, n_195, n_780, n_675, n_2624, n_903, n_1540, n_1977, n_1802, n_1504, n_2350, n_2804, n_2453, n_286, n_254, n_2193, n_2676, n_1655, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_1801, n_1886, n_2092, n_2347, n_1654, n_816, n_1157, n_3453, n_1750, n_2994, n_1462, n_3410, n_3153, n_3428, n_1188, n_1752, n_877, n_1813, n_2514, n_2206, n_604, n_2810, n_2967, n_2319, n_2519, n_825, n_728, n_2916, n_3415, n_1063, n_1588, n_2963, n_2947, n_2467, n_26, n_2602, n_2468, n_55, n_267, n_3145, n_1124, n_1624, n_515, n_2096, n_2980, n_1965, n_2476, n_3280, n_598, n_3434, n_696, n_1515, n_961, n_437, n_1082, n_1317, n_3227, n_2733, n_2824, n_3289, n_593, n_514, n_687, n_697, n_890, n_637, n_2377, n_295, n_701, n_2178, n_3271, n_950, n_388, n_190, n_2812, n_484, n_2644, n_2036, n_3326, n_2976, n_2152, n_1709, n_3009, n_2652, n_3460, n_2411, n_2525, n_1825, n_2393, n_1757, n_1796, n_170, n_2657, n_1792, n_891, n_2067, n_2136, n_2921, n_2409, n_2082, n_2252, n_1412, n_2497, n_2687, n_3237, n_949, n_1630, n_678, n_2887, n_283, n_2075, n_2194, n_2972, n_2619, n_3139, n_91, n_2763, n_2762, n_1987, n_507, n_968, n_909, n_1369, n_881, n_2271, n_1008, n_3192, n_760, n_1546, n_2583, n_590, n_63, n_2606, n_362, n_148, n_2279, n_161, n_22, n_462, n_1033, n_1052, n_2794, n_1296, n_2663, n_1990, n_3352, n_2391, n_304, n_2431, n_3073, n_2987, n_694, n_2938, n_2150, n_1294, n_2943, n_1420, n_125, n_1634, n_2078, n_3252, n_2932, n_297, n_595, n_627, n_1767, n_1779, n_524, n_1465, n_3253, n_3337, n_3431, n_342, n_3209, n_3450, n_2622, n_1858, n_1044, n_2658, n_2665, n_2165, n_2133, n_1712, n_3021, n_1391, n_449, n_131, n_1523, n_2558, n_2750, n_2775, n_1208, n_2893, n_1164, n_1295, n_1627, n_2954, n_2728, n_2349, n_3128, n_2684, n_2712, n_1072, n_3146, n_1527, n_1495, n_1438, n_495, n_815, n_1100, n_585, n_1487, n_2691, n_3421, n_840, n_2913, n_874, n_1756, n_3183, n_1128, n_2493, n_382, n_673, n_2230, n_2705, n_1969, n_2690, n_1071, n_1067, n_1565, n_1493, n_2145, n_3405, n_1968, n_898, n_255, n_284, n_1952, n_865, n_2573, n_3423, n_2646, n_3436, n_925, n_1932, n_1101, n_15, n_1026, n_1880, n_2535, n_3366, n_3442, n_2631, n_38, n_289, n_1364, n_3078, n_2436, n_615, n_2870, n_1249, n_2706, n_59, n_1293, n_2693, n_1127, n_1512, n_2151, n_3159, n_1451, n_320, n_108, n_639, n_963, n_794, n_2767, n_727, n_894, n_1839, n_2341, n_685, n_1765, n_353, n_2707, n_3240, n_605, n_1514, n_1863, n_826, n_3385, n_3037, n_1646, n_3293, n_872, n_1139, n_1714, n_86, n_3179, n_104, n_718, n_1018, n_3400, n_1521, n_1366, n_542, n_847, n_644, n_682, n_851, n_2537, n_2897, n_305, n_72, n_2554, n_996, n_532, n_173, n_1308, n_2089, n_1376, n_1513, n_2747, n_413, n_3171, n_791, n_1913, n_510, n_837, n_2097, n_79, n_2170, n_3459, n_1488, n_2853, n_1808, n_3053, n_948, n_3358, n_2517, n_2713, n_704, n_2148, n_977, n_2339, n_1005, n_1947, n_2765, n_2861, n_536, n_3158, n_1788, n_3426, n_1999, n_2731, n_622, n_147, n_2590, n_2643, n_3150, n_3018, n_3353, n_1469, n_2060, n_2608, n_1838, n_2638, n_1835, n_1766, n_1776, n_1959, n_3133, n_2002, n_581, n_2650, n_2138, n_765, n_432, n_987, n_1492, n_2414, n_1340, n_3014, n_3166, n_1771, n_2316, n_3104, n_631, n_720, n_3435, n_153, n_842, n_3148, n_2262, n_3229, n_3348, n_1707, n_2239, n_3082, n_1432, n_156, n_145, n_2208, n_843, n_656, n_989, n_2604, n_2407, n_1277, n_2816, n_797, n_2689, n_2933, n_1473, n_2191, n_1723, n_2717, n_1246, n_1878, n_2574, n_899, n_189, n_738, n_2012, n_1304, n_1035, n_294, n_2842, n_499, n_2675, n_1426, n_3418, n_705, n_11, n_1004, n_1176, n_2134, n_1529, n_2335, n_2473, n_1022, n_614, n_529, n_2069, n_2307, n_2362, n_425, n_684, n_2539, n_2667, n_2698, n_1431, n_1615, n_1474, n_3312, n_1571, n_1809, n_3119, n_2948, n_1577, n_2958, n_2297, n_1181, n_2119, n_1822, n_37, n_486, n_947, n_2936, n_3224, n_1117, n_2489, n_1087, n_1448, n_3173, n_1992, n_648, n_657, n_1049, n_3223, n_2771, n_2445, n_3020, n_2057, n_2103, n_3140, n_3185, n_2605, n_1666, n_2772, n_1505, n_803, n_290, n_118, n_1717, n_926, n_1817, n_2449, n_927, n_2610, n_3129, n_1849, n_2848, n_919, n_2868, n_1698, n_478, n_2231, n_929, n_107, n_2520, n_1228, n_417, n_2857, n_446, n_89, n_1568, n_1490, n_2372, n_777, n_1299, n_272, n_2896, n_526, n_2718, n_3019, n_2639, n_1183, n_1436, n_2898, n_2251, n_1384, n_69, n_2494, n_2959, n_2501, n_3203, n_3325, n_2238, n_293, n_2368, n_53, n_458, n_1070, n_2403, n_3342, n_2837, n_998, n_16, n_717, n_3200, n_1665, n_18, n_3259, n_2524, n_154, n_3167, n_1383, n_2460, n_3390, n_1178, n_98, n_2127, n_1424, n_2338, n_3324, n_3341, n_1073, n_1000, n_796, n_252, n_1195, n_3025, n_2137, n_1626, n_3191, n_1507, n_2482, n_184, n_552, n_2532, n_1358, n_1811, n_1388, n_3006, n_216, n_2481, n_912, n_1857, n_1519, n_2144, n_3056, n_745, n_1284, n_1604, n_2296, n_2424, n_3201, n_3447, n_1142, n_2849, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1774, n_2354, n_2682, n_3032, n_3103, n_2589, n_1395, n_2110, n_2199, n_2661, n_731, n_2877, n_1502, n_1659, n_1955, n_755, n_931, n_1021, n_3393, n_474, n_527, n_683, n_811, n_1207, n_2442, n_312, n_1791, n_1368, n_66, n_3451, n_1418, n_958, n_292, n_1250, n_100, n_3331, n_1137, n_1897, n_2064, n_880, n_3072, n_3087, n_2053, n_2259, n_2121, n_2773, n_2545, n_889, n_2432, n_2710, n_150, n_1478, n_589, n_1310, n_3142, n_819, n_2966, n_2294, n_1363, n_2581, n_1334, n_1942, n_1966, n_767, n_1314, n_600, n_964, n_831, n_1837, n_2218, n_2788, n_477, n_3196, n_2435, n_954, n_864, n_2504, n_2797, n_2623, n_1110, n_2213, n_1410, n_399, n_2389, n_1440, n_124, n_2132, n_2892, n_2063, n_1382, n_1534, n_1564, n_1736, n_211, n_2748, n_1483, n_1834, n_2331, n_1372, n_231, n_2292, n_2860, n_3327, n_2330, n_40, n_3441, n_1457, n_505, n_1719, n_319, n_1339, n_1787, n_2701, n_2475, n_537, n_2511, n_1993, n_2281, n_1427, n_311, n_2416, n_2745, n_2617, n_2776, n_1466, n_10, n_403, n_1919, n_1080, n_723, n_1877, n_3144, n_3211, n_3244, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1939, n_2030, n_1769, n_1220, n_2323, n_1893, n_556, n_2784, n_2209, n_2301, n_162, n_3287, n_2387, n_3322, n_1755, n_1602, n_2421, n_1136, n_3270, n_2618, n_2025, n_2357, n_2846, n_2464, n_3265, n_128, n_1125, n_970, n_3306, n_2488, n_2224, n_1980, n_642, n_995, n_276, n_1159, n_2329, n_1092, n_2237, n_3026, n_441, n_221, n_1060, n_1951, n_2250, n_3090, n_444, n_3033, n_146, n_1252, n_1784, n_3311, n_1223, n_303, n_511, n_2990, n_193, n_1286, n_1773, n_1775, n_2115, n_2410, n_2552, n_1053, n_3302, n_2374, n_416, n_1681, n_520, n_418, n_1093, n_113, n_1783, n_1533, n_1597, n_2929, n_2780, n_3226, n_3323, n_3364, n_4, n_266, n_296, n_2596, n_2274, n_3163, n_775, n_651, n_1153, n_439, n_1618, n_3407, n_217, n_518, n_1531, n_2828, n_1185, n_453, n_3425, n_215, n_2384, n_1745, n_914, n_759, n_3127, n_2724, n_1831, n_426, n_317, n_2585, n_2621, n_1653, n_2352, n_1679, n_1625, n_90, n_2601, n_2160, n_3454, n_54, n_1453, n_2146, n_2226, n_2131, n_488, n_2502, n_2801, n_497, n_2920, n_773, n_1901, n_920, n_99, n_1374, n_2556, n_2648, n_3212, n_1315, n_1647, n_13, n_2575, n_2754, n_1224, n_2783, n_2306, n_1614, n_1459, n_1892, n_3188, n_1933, n_2462, n_1135, n_1169, n_1179, n_2889, n_3243, n_401, n_324, n_1617, n_3260, n_3370, n_3386, n_335, n_1470, n_2550, n_463, n_3093, n_3175, n_3214, n_1243, n_848, n_120, n_2732, n_301, n_2928, n_274, n_1096, n_2249, n_1091, n_1917, n_2000, n_1580, n_2227, n_2270, n_2822, n_1425, n_3169, n_36, n_3205, n_1881, n_1267, n_1281, n_1806, n_3284, n_983, n_3109, n_2023, n_3354, n_427, n_2572, n_2204, n_1520, n_496, n_2720, n_3126, n_2159, n_906, n_1390, n_688, n_2289, n_1077, n_1733, n_2315, n_1419, n_2863, n_3299, n_351, n_2955, n_2995, n_259, n_1731, n_177, n_2158, n_2087, n_1855, n_1636, n_3051, n_1437, n_3360, n_2135, n_3367, n_1645, n_1832, n_385, n_1687, n_1439, n_2328, n_1323, n_2859, n_2202, n_858, n_2049, n_1331, n_613, n_736, n_2627, n_501, n_956, n_960, n_2276, n_3234, n_663, n_856, n_2803, n_2100, n_3314, n_379, n_2993, n_778, n_1668, n_2777, n_1134, n_3016, n_3004, n_3202, n_2830, n_2781, n_3220, n_410, n_1129, n_554, n_602, n_1696, n_2829, n_1995, n_1594, n_2181, n_664, n_1869, n_171, n_2911, n_1764, n_169, n_1429, n_2826, n_1610, n_3084, n_3429, n_1889, n_2379, n_435, n_1905, n_2016, n_2343, n_793, n_326, n_587, n_1593, n_580, n_762, n_1030, n_1202, n_1937, n_465, n_1790, n_1778, n_1635, n_2942, n_1079, n_341, n_2515, n_1744, n_828, n_2139, n_2142, n_607, n_316, n_419, n_28, n_1551, n_2448, n_1103, n_2875, n_2555, n_3338, n_144, n_3462, n_2219, n_1203, n_2851, n_3406, n_820, n_2327, n_951, n_106, n_2201, n_725, n_952, n_999, n_358, n_1254, n_160, n_2841, n_3349, n_2420, n_186, n_2984, n_0, n_368, n_575, n_994, n_2263, n_3291, n_2304, n_1508, n_2487, n_732, n_974, n_2983, n_2240, n_392, n_2278, n_2656, n_2538, n_724, n_2597, n_2375, n_3113, n_3194, n_3250, n_1934, n_3276, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_1728, n_557, n_2756, n_1871, n_349, n_3448, n_617, n_845, n_807, n_2924, n_1036, n_140, n_1138, n_3414, n_1661, n_1275, n_2884, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_421, n_3120, n_1468, n_2855, n_1859, n_2102, n_2563, n_238, n_1095, n_2024, n_1595, n_202, n_2156, n_3449, n_1718, n_1749, n_1683, n_1916, n_2598, n_597, n_280, n_1270, n_2549, n_1187, n_610, n_1403, n_1669, n_1852, n_1024, n_1768, n_2153, n_2544, n_2381, n_198, n_1847, n_2052, n_179, n_248, n_2302, n_517, n_1667, n_667, n_1206, n_3230, n_621, n_1037, n_1397, n_3268, n_3236, n_1279, n_1115, n_750, n_901, n_1499, n_468, n_2755, n_3141, n_923, n_504, n_1409, n_1841, n_2637, n_2823, n_1639, n_1623, n_183, n_1015, n_1503, n_3112, n_2819, n_3195, n_466, n_2526, n_3041, n_2423, n_1057, n_3277, n_3108, n_2548, n_603, n_991, n_2785, n_1657, n_235, n_1126, n_2412, n_1997, n_3417, n_2636, n_3131, n_340, n_710, n_1108, n_1818, n_2439, n_2404, n_1182, n_1298, n_2559, n_2177, n_39, n_2595, n_3399, n_2088, n_73, n_1611, n_785, n_2740, n_746, n_609, n_1601, n_3011, n_1960, n_2694, n_2061, n_3416, n_1686, n_2757, n_2337, n_2401, n_101, n_167, n_1356, n_1589, n_3042, n_3213, n_127, n_2309, n_2900, n_2957, n_2607, n_1740, n_2737, n_1497, n_2890, n_1168, n_1216, n_1943, n_3228, n_133, n_1320, n_2716, n_96, n_3249, n_3081, n_2452, n_1430, n_1316, n_1287, n_2722, n_1452, n_2854, n_3010, n_2499, n_3043, n_1622, n_1586, n_2543, n_2264, n_3464, n_302, n_1694, n_380, n_1535, n_3137, n_3382, n_2486, n_3132, n_137, n_2571, n_3138, n_1596, n_3177, n_20, n_1190, n_1734, n_3172, n_397, n_2902, n_3217, n_1983, n_1938, n_2498, n_122, n_2220, n_2577, n_34, n_1262, n_2472, n_218, n_1891, n_2171, n_1213, n_3238, n_70, n_2235, n_3394, n_2988, n_3136, n_1350, n_1673, n_2232, n_1715, n_172, n_1443, n_1272, n_2392, n_2894, n_3424, n_2790, n_239, n_2037, n_97, n_2808, n_2298, n_782, n_2326, n_1539, n_490, n_220, n_809, n_1043, n_3040, n_1797, n_3279, n_1608, n_986, n_2305, n_2120, n_80, n_1472, n_2050, n_2373, n_2164, n_2402, n_2225, n_1081, n_402, n_1870, n_352, n_2964, n_1692, n_800, n_1084, n_1171, n_460, n_2169, n_2371, n_1827, n_1361, n_1864, n_2006, n_3402, n_1491, n_2187, n_662, n_374, n_1152, n_1840, n_1705, n_450, n_3262, n_2904, n_2244, n_3013, n_3356, n_2586, n_1684, n_921, n_2446, n_1346, n_711, n_1642, n_579, n_1352, n_2789, n_3105, n_3210, n_2872, n_937, n_2257, n_1682, n_2017, n_370, n_1695, n_1828, n_2046, n_2272, n_2699, n_2200, n_3029, n_650, n_1046, n_2560, n_1940, n_1979, n_2760, n_2704, n_3329, n_1145, n_330, n_1121, n_1102, n_1963, n_2738, n_972, n_1405, n_2376, n_258, n_1406, n_456, n_2766, n_1332, n_260, n_2670, n_313, n_2700, n_624, n_962, n_1041, n_2346, n_565, n_3134, n_356, n_1569, n_936, n_3045, n_3115, n_1883, n_1288, n_3318, n_1186, n_1062, n_885, n_896, n_83, n_3278, n_2342, n_2167, n_2084, n_2970, n_2882, n_3320, n_2541, n_654, n_2940, n_411, n_2518, n_2458, n_152, n_1222, n_599, n_776, n_321, n_1823, n_2479, n_3050, n_3350, n_105, n_2782, n_227, n_1974, n_2673, n_2456, n_1720, n_2527, n_204, n_482, n_934, n_1637, n_2635, n_3307, n_3439, n_1407, n_1795, n_2768, n_2871, n_420, n_2688, n_1341, n_394, n_1456, n_1845, n_1489, n_164, n_2314, n_23, n_942, n_3003, n_2798, n_2852, n_1524, n_543, n_2229, n_1964, n_2288, n_1920, n_2753, n_2099, n_1496, n_1271, n_3292, n_1545, n_2007, n_3121, n_2039, n_3388, n_1946, n_1355, n_1225, n_3184, n_1544, n_1485, n_2258, n_325, n_1640, n_804, n_464, n_1846, n_3437, n_3245, n_3075, n_2406, n_533, n_2390, n_806, n_879, n_959, n_2310, n_2506, n_584, n_2141, n_2562, n_244, n_2642, n_1343, n_1522, n_76, n_2734, n_548, n_1782, n_94, n_282, n_2383, n_2626, n_1676, n_833, n_1830, n_2351, n_1567, n_523, n_1319, n_707, n_2986, n_345, n_1900, n_3246, n_799, n_1548, n_3381, n_3044, n_2973, n_1155, n_2536, n_139, n_2196, n_41, n_2629, n_273, n_1633, n_2195, n_3208, n_2809, n_3007, n_787, n_2172, n_2835, n_1416, n_1528, n_2820, n_2293, n_1146, n_2021, n_3355, n_2454, n_2114, n_3074, n_3174, n_159, n_1086, n_1066, n_3102, n_1948, n_157, n_2125, n_2026, n_1282, n_2561, n_550, n_3321, n_2567, n_2322, n_275, n_652, n_2154, n_2727, n_2962, n_3377, n_2939, n_560, n_1906, n_1484, n_2992, n_3305, n_1241, n_1321, n_1672, n_569, n_2533, n_3157, n_1758, n_3221, n_3267, n_2283, n_2869, n_2422, n_1925, n_737, n_1318, n_1914, n_1235, n_3457, n_1229, n_2759, n_2945, n_3061, n_2361, n_306, n_1292, n_1373, n_21, n_2266, n_2960, n_3005, n_346, n_3, n_2427, n_3151, n_3411, n_1029, n_1447, n_2388, n_2056, n_790, n_2611, n_2901, n_138, n_3258, n_1706, n_3389, n_1498, n_3143, n_2653, n_2417, n_3000, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_2189, n_2680, n_2246, n_1047, n_3149, n_3375, n_1984, n_3365, n_2236, n_1385, n_431, n_3379, n_3156, n_24, n_459, n_1269, n_1931, n_2083, n_2834, n_3207, n_502, n_2668, n_672, n_2441, n_1257, n_3008, n_1751, n_3401, n_2840, n_3197, n_3242, n_285, n_1375, n_1941, n_85, n_2128, n_655, n_706, n_1045, n_1650, n_786, n_1794, n_1236, n_1962, n_1559, n_1725, n_1928, n_2398, n_1872, n_3091, n_834, n_19, n_29, n_2695, n_75, n_743, n_766, n_3124, n_430, n_1741, n_1325, n_1002, n_1746, n_1949, n_3398, n_545, n_2671, n_489, n_2761, n_2885, n_2793, n_2715, n_2888, n_1804, n_2923, n_1727, n_251, n_2508, n_1019, n_636, n_2054, n_729, n_110, n_151, n_876, n_774, n_2845, n_1337, n_3097, n_660, n_2062, n_2041, n_2975, n_438, n_1477, n_1360, n_2839, n_1860, n_2856, n_1904, n_2874, n_1200, n_2070, n_2588, n_479, n_1607, n_1353, n_1777, n_1908, n_1454, n_2484, n_2348, n_2944, n_2614, n_2126, n_869, n_1154, n_3308, n_1113, n_1600, n_2833, n_2253, n_2758, n_2366, n_646, n_528, n_391, n_1098, n_2937, n_1329, n_2045, n_817, n_2261, n_2216, n_2210, n_262, n_187, n_897, n_846, n_3300, n_2978, n_2066, n_841, n_1476, n_2516, n_3391, n_1001, n_508, n_1800, n_2241, n_1050, n_1411, n_1463, n_2903, n_2827, n_1177, n_3216, n_3458, n_332, n_1150, n_1742, n_3190, n_1562, n_1690, n_398, n_1191, n_1826, n_566, n_1023, n_1882, n_2951, n_1076, n_1118, n_194, n_2949, n_57, n_1007, n_1807, n_1929, n_1378, n_2369, n_855, n_1592, n_1759, n_2719, n_1814, n_1631, n_52, n_591, n_1377, n_1879, n_256, n_853, n_440, n_695, n_1542, n_2587, n_3199, n_2931, n_875, n_209, n_367, n_680, n_3339, n_1678, n_2569, n_661, n_2400, n_1716, n_278, n_1256, n_671, n_1953, n_7, n_933, n_740, n_703, n_3343, n_3303, n_978, n_2752, n_384, n_3135, n_1976, n_2905, n_1291, n_1217, n_751, n_749, n_1824, n_310, n_1628, n_1324, n_1399, n_2122, n_2109, n_1435, n_969, n_988, n_2140, n_3160, n_1065, n_2796, n_3255, n_2507, n_84, n_1401, n_2358, n_1255, n_568, n_1516, n_143, n_1536, n_180, n_2163, n_2186, n_2029, n_2815, n_1204, n_3034, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_2528, n_2814, n_214, n_246, n_2787, n_1338, n_1097, n_2969, n_2395, n_935, n_3027, n_781, n_789, n_1554, n_3231, n_1130, n_3083, n_2979, n_181, n_1810, n_182, n_2953, n_573, n_769, n_2380, n_676, n_327, n_1120, n_832, n_1583, n_3049, n_1730, n_2295, n_555, n_389, n_814, n_2746, n_2946, n_1643, n_2020, n_2500, n_3430, n_2269, n_1729, n_669, n_2290, n_2048, n_176, n_114, n_300, n_222, n_2005, n_747, n_74, n_2565, n_1389, n_1105, n_3117, n_721, n_1461, n_742, n_3432, n_535, n_691, n_372, n_2076, n_2736, n_111, n_2883, n_314, n_1408, n_378, n_1196, n_377, n_1598, n_2935, n_863, n_3015, n_2175, n_601, n_2182, n_338, n_2910, n_1283, n_2385, n_918, n_748, n_506, n_1114, n_1785, n_56, n_763, n_1147, n_1848, n_360, n_1754, n_2149, n_3057, n_3154, n_2396, n_1506, n_119, n_2584, n_1652, n_1812, n_957, n_1994, n_895, n_866, n_1227, n_2450, n_2485, n_2284, n_191, n_2566, n_387, n_2287, n_452, n_744, n_971, n_2702, n_3241, n_946, n_344, n_2906, n_761, n_1303, n_2769, n_1205, n_2492, n_1258, n_2438, n_2914, n_1392, n_174, n_1173, n_1924, n_525, n_2463, n_3363, n_2881, n_1677, n_1116, n_611, n_1570, n_1702, n_1219, n_3064, n_1780, n_3100, n_1689, n_8, n_2180, n_3372, n_2858, n_3062, n_2679, n_1174, n_1944, n_1016, n_1347, n_795, n_1501, n_1221, n_3334, n_1245, n_838, n_3215, n_129, n_3336, n_647, n_197, n_844, n_17, n_448, n_2952, n_1017, n_3068, n_2117, n_2234, n_2779, n_2685, n_1083, n_109, n_445, n_1561, n_2741, n_3114, n_930, n_888, n_2275, n_1112, n_2465, n_2620, n_2081, n_2168, n_2568, n_234, n_2022, n_1945, n_2203, n_910, n_1656, n_1721, n_1460, n_911, n_2112, n_2255, n_82, n_1464, n_27, n_236, n_653, n_1737, n_2430, n_1414, n_752, n_908, n_2649, n_2721, n_944, n_2034, n_576, n_1028, n_2106, n_472, n_2862, n_270, n_2265, n_2615, n_414, n_2683, n_1922, n_563, n_2032, n_2744, n_1011, n_2474, n_1566, n_1215, n_2437, n_25, n_93, n_839, n_2444, n_2743, n_708, n_1973, n_3181, n_2267, n_3456, n_3035, n_668, n_626, n_990, n_1500, n_779, n_1537, n_1821, n_2205, n_3204, n_1104, n_854, n_1058, n_3378, n_2312, n_498, n_3404, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_2242, n_3362, n_1509, n_103, n_3328, n_1693, n_2934, n_3290, n_1109, n_185, n_2222, n_712, n_3256, n_348, n_1276, n_3176, n_376, n_3309, n_2015, n_2118, n_2111, n_2466, n_390, n_2915, n_2530, n_1148, n_31, n_2188, n_2505, n_334, n_1989, n_1161, n_2609, n_1085, n_232, n_2802, n_2999, n_2014, n_2042, n_46, n_1239, n_771, n_1584, n_2425, n_470, n_475, n_924, n_3408, n_3461, n_298, n_1582, n_492, n_2318, n_3286, n_2408, n_1149, n_3170, n_265, n_1184, n_2483, n_2950, n_228, n_719, n_1972, n_3060, n_3304, n_2592, n_1525, n_3098, n_2594, n_455, n_2666, n_1585, n_1851, n_363, n_1799, n_1090, n_2147, n_2564, n_592, n_1816, n_2503, n_2433, n_1518, n_829, n_1156, n_1362, n_3123, n_393, n_984, n_2600, n_3380, n_1829, n_503, n_2035, n_3024, n_1450, n_1638, n_3422, n_132, n_868, n_3038, n_570, n_859, n_2033, n_406, n_3086, n_735, n_1789, n_2531, n_1770, n_878, n_620, n_130, n_3285, n_519, n_2523, n_307, n_469, n_1218, n_2413, n_500, n_1482, n_3361, n_981, n_714, n_1349, n_291, n_1144, n_2071, n_357, n_3219, n_2429, n_3130, n_985, n_2233, n_2440, n_2723, n_481, n_3233, n_997, n_1710, n_2800, n_2161, n_1301, n_2805, n_802, n_561, n_33, n_3310, n_980, n_2681, n_1306, n_3264, n_2010, n_2282, n_1651, n_1198, n_3096, n_2360, n_2047, n_2651, n_2095, n_3239, n_1609, n_2174, n_3161, n_2799, n_436, n_116, n_3344, n_2334, n_3295, n_409, n_1244, n_1685, n_1763, n_1998, n_3066, n_1574, n_2426, n_2490, n_2844, n_3101, n_240, n_756, n_2303, n_1619, n_2478, n_1981, n_2285, n_1606, n_810, n_1133, n_635, n_95, n_1194, n_3374, n_2742, n_2640, n_1051, n_253, n_1552, n_2918, n_583, n_3288, n_1996, n_2367, n_249, n_201, n_2867, n_3198, n_1039, n_1442, n_2726, n_1034, n_2043, n_1480, n_3125, n_1158, n_2909, n_2248, n_754, n_941, n_975, n_3206, n_1031, n_115, n_1305, n_2363, n_2578, n_553, n_43, n_849, n_2662, n_3116, n_3147, n_3383, n_753, n_1753, n_3095, n_3180, n_3359, n_2795, n_2471, n_467, n_3187, n_2540, n_269, n_359, n_973, n_2807, n_1921, n_3218, n_3330, n_1479, n_1055, n_1675, n_2197, n_2217, n_582, n_2065, n_2879, n_861, n_857, n_967, n_571, n_2215, n_2461, n_271, n_404, n_2001, n_158, n_2107, n_1884, n_206, n_2040, n_679, n_2968, n_633, n_1170, n_665, n_1629, n_2221, n_588, n_225, n_1260, n_308, n_309, n_1819, n_2055, n_1010, n_3444, n_2553, n_149, n_1040, n_915, n_632, n_3059, n_1166, n_2038, n_812, n_2891, n_1131, n_2634, n_1761, n_2709, n_3155, n_3445, n_534, n_1578, n_1006, n_1861, n_373, n_3110, n_87, n_1632, n_1890, n_3017, n_1805, n_2477, n_257, n_1557, n_1888, n_2280, n_1833, n_730, n_1311, n_1494, n_2325, n_670, n_203, n_1850, n_1898, n_2443, n_2697, n_3235, n_2308, n_2162, n_1868, n_207, n_2333, n_2079, n_3001, n_1089, n_1887, n_1587, n_2512, n_3433, n_1365, n_1417, n_205, n_1242, n_2086, n_2185, n_2927, n_1836, n_2774, n_3039, n_681, n_1226, n_3162, n_1274, n_1486, n_2166, n_3094, n_412, n_2899, n_3274, n_3333, n_3186, n_640, n_1322, n_81, n_965, n_1899, n_1428, n_1616, n_1576, n_1856, n_1862, n_1958, n_2077, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_3065, n_2632, n_422, n_2579, n_722, n_862, n_2105, n_135, n_3079, n_165, n_2098, n_3085, n_540, n_1423, n_2813, n_1935, n_3387, n_2027, n_457, n_3070, n_2223, n_2091, n_364, n_3263, n_3420, n_2991, n_1915, n_629, n_1621, n_1748, n_2547, n_2415, n_900, n_1449, n_531, n_827, n_2912, n_60, n_361, n_2659, n_2930, n_1025, n_3409, n_2419, n_3111, n_2116, n_336, n_2320, n_12, n_1885, n_2677, n_1013, n_3182, n_1259, n_3054, n_3283, n_192, n_2183, n_3002, n_1538, n_51, n_649, n_1612, n_1240, n_14691);

input n_992;
input n_2542;
input n_1671;
input n_1;
input n_2817;
input n_801;
input n_1613;
input n_1234;
input n_1458;
input n_2576;
input n_3254;
input n_1199;
input n_1674;
input n_3392;
input n_741;
input n_1027;
input n_1351;
input n_3266;
input n_625;
input n_1189;
input n_3152;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_2157;
input n_3335;
input n_2332;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_3178;
input n_2003;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_2353;
input n_2534;
input n_3089;
input n_3301;
input n_1357;
input n_1853;
input n_77;
input n_783;
input n_2451;
input n_1738;
input n_2243;
input n_798;
input n_188;
input n_1575;
input n_1854;
input n_2324;
input n_3088;
input n_3443;
input n_1923;
input n_3257;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_2260;
input n_3222;
input n_677;
input n_1708;
input n_805;
input n_1151;
input n_396;
input n_2977;
input n_1739;
input n_350;
input n_78;
input n_2051;
input n_2317;
input n_1380;
input n_2359;
input n_442;
input n_480;
input n_142;
input n_2847;
input n_1402;
input n_2557;
input n_1688;
input n_1691;
input n_3332;
input n_3465;
input n_1975;
input n_1009;
input n_1743;
input n_62;
input n_1930;
input n_2405;
input n_1160;
input n_883;
input n_2647;
input n_1238;
input n_1991;
input n_2570;
input n_2179;
input n_2386;
input n_2997;
input n_1724;
input n_1032;
input n_2336;
input n_1247;
input n_1547;
input n_2521;
input n_3376;
input n_3046;
input n_2956;
input n_1553;
input n_893;
input n_1099;
input n_2491;
input n_1264;
input n_1192;
input n_471;
input n_1844;
input n_424;
input n_1700;
input n_1555;
input n_1415;
input n_2211;
input n_1370;
input n_1786;
input n_369;
input n_287;
input n_2382;
input n_2672;
input n_3030;
input n_2291;
input n_415;
input n_830;
input n_2299;
input n_65;
input n_230;
input n_3340;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_2886;
input n_2974;
input n_200;
input n_1985;
input n_2989;
input n_447;
input n_2838;
input n_2184;
input n_3395;
input n_2982;
input n_1803;
input n_3427;
input n_1172;
input n_852;
input n_2509;
input n_71;
input n_229;
input n_2513;
input n_3282;
input n_1590;
input n_2645;
input n_1532;
input n_2313;
input n_2628;
input n_3071;
input n_1393;
input n_1517;
input n_1867;
input n_2926;
input n_1704;
input n_1078;
input n_250;
input n_544;
input n_1711;
input n_2247;
input n_3106;
input n_1140;
input n_2630;
input n_1444;
input n_1670;
input n_1603;
input n_2344;
input n_1579;
input n_3275;
input n_35;
input n_2365;
input n_2470;
input n_2321;
input n_1263;
input n_2019;
input n_3031;
input n_836;
input n_3345;
input n_375;
input n_2074;
input n_2447;
input n_522;
input n_2919;
input n_3440;
input n_2129;
input n_2340;
input n_1261;
input n_945;
input n_2286;
input n_1649;
input n_2018;
input n_2094;
input n_3080;
input n_1903;
input n_1511;
input n_1143;
input n_2356;
input n_2399;
input n_1422;
input n_1232;
input n_1772;
input n_1572;
input n_616;
input n_658;
input n_1874;
input n_3165;
input n_1119;
input n_2865;
input n_2825;
input n_3463;
input n_2013;
input n_428;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2044;
input n_1954;
input n_1735;
input n_2510;
input n_1541;
input n_1300;
input n_641;
input n_2480;
input n_2739;
input n_3023;
input n_822;
input n_3232;
input n_693;
input n_1313;
input n_2791;
input n_3251;
input n_1056;
input n_3316;
input n_2212;
input n_758;
input n_516;
input n_3048;
input n_1455;
input n_2418;
input n_2864;
input n_1163;
input n_2729;
input n_3063;
input n_1180;
input n_2256;
input n_2582;
input n_943;
input n_1798;
input n_1550;
input n_2703;
input n_491;
input n_2786;
input n_3371;
input n_1591;
input n_42;
input n_772;
input n_3122;
input n_2806;
input n_1344;
input n_3261;
input n_2730;
input n_2495;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_1781;
input n_1971;
input n_2058;
input n_2090;
input n_2603;
input n_405;
input n_213;
input n_2660;
input n_538;
input n_3028;
input n_2981;
input n_3076;
input n_2173;
input n_2004;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_3077;
input n_1345;
input n_1820;
input n_2873;
input n_3452;
input n_494;
input n_539;
input n_493;
input n_3107;
input n_155;
input n_2880;
input n_3225;
input n_2394;
input n_2108;
input n_45;
input n_454;
input n_1421;
input n_2836;
input n_1936;
input n_638;
input n_1404;
input n_1211;
input n_2124;
input n_381;
input n_2378;
input n_887;
input n_1660;
input n_1961;
input n_3047;
input n_112;
input n_1280;
input n_713;
input n_2655;
input n_1400;
input n_2625;
input n_3296;
input n_2843;
input n_126;
input n_1467;
input n_3297;
input n_58;
input n_976;
input n_3067;
input n_2155;
input n_224;
input n_2686;
input n_48;
input n_1445;
input n_2364;
input n_2551;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_1894;
input n_196;
input n_1231;
input n_2996;
input n_2599;
input n_2985;
input n_1978;
input n_2085;
input n_3368;
input n_917;
input n_574;
input n_9;
input n_3347;
input n_2370;
input n_2612;
input n_907;
input n_6;
input n_1446;
input n_14;
input n_2591;
input n_659;
input n_1815;
input n_2214;
input n_3351;
input n_407;
input n_913;
input n_1658;
input n_2593;
input n_808;
input n_867;
input n_3269;
input n_1230;
input n_3413;
input n_473;
input n_1193;
input n_1967;
input n_1054;
input n_559;
input n_3412;
input n_2613;
input n_1333;
input n_2496;
input n_44;
input n_2708;
input n_3313;
input n_1648;
input n_3189;
input n_1911;
input n_1956;
input n_163;
input n_1644;
input n_2011;
input n_2725;
input n_2277;
input n_3164;
input n_1558;
input n_1732;
input n_281;
input n_551;
input n_699;
input n_1986;
input n_2300;
input n_564;
input n_2397;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_1641;
input n_2113;
input n_1918;
input n_2190;
input n_2907;
input n_577;
input n_3438;
input n_166;
input n_2735;
input n_1843;
input n_619;
input n_2268;
input n_1367;
input n_1336;
input n_521;
input n_2778;
input n_2850;
input n_572;
input n_395;
input n_813;
input n_1909;
input n_2080;
input n_1481;
input n_323;
input n_606;
input n_1441;
input n_818;
input n_3373;
input n_1123;
input n_1309;
input n_92;
input n_2104;
input n_513;
input n_645;
input n_1381;
input n_2961;
input n_331;
input n_1699;
input n_916;
input n_2093;
input n_2633;
input n_483;
input n_102;
input n_2207;
input n_1970;
input n_2770;
input n_608;
input n_261;
input n_2101;
input n_2696;
input n_630;
input n_2059;
input n_32;
input n_2198;
input n_3319;
input n_541;
input n_512;
input n_2669;
input n_2925;
input n_2073;
input n_2273;
input n_121;
input n_433;
input n_2546;
input n_3272;
input n_3193;
input n_792;
input n_2522;
input n_476;
input n_2792;
input n_2;
input n_1328;
input n_3396;
input n_1957;
input n_2917;
input n_219;
input n_2616;
input n_3118;
input n_3315;
input n_1907;
input n_2529;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_1530;
input n_788;
input n_939;
input n_1543;
input n_821;
input n_2811;
input n_938;
input n_1302;
input n_1068;
input n_1599;
input n_329;
input n_982;
input n_2674;
input n_2832;
input n_549;
input n_1762;
input n_1910;
input n_1075;
input n_408;
input n_932;
input n_2831;
input n_2998;
input n_3446;
input n_61;
input n_3317;
input n_237;
input n_1876;
input n_1895;
input n_2123;
input n_1697;
input n_2143;
input n_243;
input n_979;
input n_1873;
input n_905;
input n_1866;
input n_1680;
input n_117;
input n_175;
input n_322;
input n_993;
input n_2692;
input n_689;
input n_3248;
input n_2031;
input n_354;
input n_2130;
input n_1330;
input n_1413;
input n_1605;
input n_2228;
input n_3397;
input n_134;
input n_1988;
input n_2941;
input n_1278;
input n_547;
input n_2455;
input n_2876;
input n_558;
input n_2654;
input n_3036;
input n_2469;
input n_1064;
input n_3099;
input n_1396;
input n_634;
input n_2355;
input n_136;
input n_966;
input n_2908;
input n_3168;
input n_764;
input n_2751;
input n_2764;
input n_3357;
input n_1663;
input n_2895;
input n_2009;
input n_692;
input n_3403;
input n_733;
input n_1793;
input n_2922;
input n_1233;
input n_1289;
input n_2714;
input n_2245;
input n_487;
input n_3055;
input n_3092;
input n_241;
input n_30;
input n_2068;
input n_1107;
input n_2866;
input n_2457;
input n_3294;
input n_1014;
input n_1290;
input n_1703;
input n_2580;
input n_3455;
input n_882;
input n_2176;
input n_2072;
input n_1354;
input n_2821;
input n_586;
input n_423;
input n_1865;
input n_1875;
input n_1701;
input n_2459;
input n_318;
input n_1111;
input n_1713;
input n_2971;
input n_715;
input n_2678;
input n_1251;
input n_3384;
input n_1265;
input n_2711;
input n_88;
input n_1726;
input n_1950;
input n_530;
input n_1563;
input n_1912;
input n_277;
input n_2434;
input n_3369;
input n_3419;
input n_1982;
input n_2878;
input n_618;
input n_3012;
input n_1297;
input n_1662;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_2818;
input n_2428;
input n_674;
input n_3247;
input n_871;
input n_3069;
input n_922;
input n_268;
input n_1335;
input n_1760;
input n_1927;
input n_210;
input n_2028;
input n_1069;
input n_2664;
input n_5;
input n_1664;
input n_1722;
input n_612;
input n_2641;
input n_3022;
input n_3052;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_2008;
input n_2749;
input n_3298;
input n_2192;
input n_3281;
input n_2254;
input n_2345;
input n_3346;
input n_1926;
input n_1175;
input n_3273;
input n_328;
input n_1386;
input n_2311;
input n_1896;
input n_429;
input n_2965;
input n_1747;
input n_3058;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_2624;
input n_903;
input n_1540;
input n_1977;
input n_1802;
input n_1504;
input n_2350;
input n_2804;
input n_2453;
input n_286;
input n_254;
input n_2193;
input n_2676;
input n_1655;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_1801;
input n_1886;
input n_2092;
input n_2347;
input n_1654;
input n_816;
input n_1157;
input n_3453;
input n_1750;
input n_2994;
input n_1462;
input n_3410;
input n_3153;
input n_3428;
input n_1188;
input n_1752;
input n_877;
input n_1813;
input n_2514;
input n_2206;
input n_604;
input n_2810;
input n_2967;
input n_2319;
input n_2519;
input n_825;
input n_728;
input n_2916;
input n_3415;
input n_1063;
input n_1588;
input n_2963;
input n_2947;
input n_2467;
input n_26;
input n_2602;
input n_2468;
input n_55;
input n_267;
input n_3145;
input n_1124;
input n_1624;
input n_515;
input n_2096;
input n_2980;
input n_1965;
input n_2476;
input n_3280;
input n_598;
input n_3434;
input n_696;
input n_1515;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_3227;
input n_2733;
input n_2824;
input n_3289;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_2377;
input n_295;
input n_701;
input n_2178;
input n_3271;
input n_950;
input n_388;
input n_190;
input n_2812;
input n_484;
input n_2644;
input n_2036;
input n_3326;
input n_2976;
input n_2152;
input n_1709;
input n_3009;
input n_2652;
input n_3460;
input n_2411;
input n_2525;
input n_1825;
input n_2393;
input n_1757;
input n_1796;
input n_170;
input n_2657;
input n_1792;
input n_891;
input n_2067;
input n_2136;
input n_2921;
input n_2409;
input n_2082;
input n_2252;
input n_1412;
input n_2497;
input n_2687;
input n_3237;
input n_949;
input n_1630;
input n_678;
input n_2887;
input n_283;
input n_2075;
input n_2194;
input n_2972;
input n_2619;
input n_3139;
input n_91;
input n_2763;
input n_2762;
input n_1987;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_2271;
input n_1008;
input n_3192;
input n_760;
input n_1546;
input n_2583;
input n_590;
input n_63;
input n_2606;
input n_362;
input n_148;
input n_2279;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_2794;
input n_1296;
input n_2663;
input n_1990;
input n_3352;
input n_2391;
input n_304;
input n_2431;
input n_3073;
input n_2987;
input n_694;
input n_2938;
input n_2150;
input n_1294;
input n_2943;
input n_1420;
input n_125;
input n_1634;
input n_2078;
input n_3252;
input n_2932;
input n_297;
input n_595;
input n_627;
input n_1767;
input n_1779;
input n_524;
input n_1465;
input n_3253;
input n_3337;
input n_3431;
input n_342;
input n_3209;
input n_3450;
input n_2622;
input n_1858;
input n_1044;
input n_2658;
input n_2665;
input n_2165;
input n_2133;
input n_1712;
input n_3021;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_2558;
input n_2750;
input n_2775;
input n_1208;
input n_2893;
input n_1164;
input n_1295;
input n_1627;
input n_2954;
input n_2728;
input n_2349;
input n_3128;
input n_2684;
input n_2712;
input n_1072;
input n_3146;
input n_1527;
input n_1495;
input n_1438;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_1487;
input n_2691;
input n_3421;
input n_840;
input n_2913;
input n_874;
input n_1756;
input n_3183;
input n_1128;
input n_2493;
input n_382;
input n_673;
input n_2230;
input n_2705;
input n_1969;
input n_2690;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_2145;
input n_3405;
input n_1968;
input n_898;
input n_255;
input n_284;
input n_1952;
input n_865;
input n_2573;
input n_3423;
input n_2646;
input n_3436;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_1026;
input n_1880;
input n_2535;
input n_3366;
input n_3442;
input n_2631;
input n_38;
input n_289;
input n_1364;
input n_3078;
input n_2436;
input n_615;
input n_2870;
input n_1249;
input n_2706;
input n_59;
input n_1293;
input n_2693;
input n_1127;
input n_1512;
input n_2151;
input n_3159;
input n_1451;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_2767;
input n_727;
input n_894;
input n_1839;
input n_2341;
input n_685;
input n_1765;
input n_353;
input n_2707;
input n_3240;
input n_605;
input n_1514;
input n_1863;
input n_826;
input n_3385;
input n_3037;
input n_1646;
input n_3293;
input n_872;
input n_1139;
input n_1714;
input n_86;
input n_3179;
input n_104;
input n_718;
input n_1018;
input n_3400;
input n_1521;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_2537;
input n_2897;
input n_305;
input n_72;
input n_2554;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_2089;
input n_1376;
input n_1513;
input n_2747;
input n_413;
input n_3171;
input n_791;
input n_1913;
input n_510;
input n_837;
input n_2097;
input n_79;
input n_2170;
input n_3459;
input n_1488;
input n_2853;
input n_1808;
input n_3053;
input n_948;
input n_3358;
input n_2517;
input n_2713;
input n_704;
input n_2148;
input n_977;
input n_2339;
input n_1005;
input n_1947;
input n_2765;
input n_2861;
input n_536;
input n_3158;
input n_1788;
input n_3426;
input n_1999;
input n_2731;
input n_622;
input n_147;
input n_2590;
input n_2643;
input n_3150;
input n_3018;
input n_3353;
input n_1469;
input n_2060;
input n_2608;
input n_1838;
input n_2638;
input n_1835;
input n_1766;
input n_1776;
input n_1959;
input n_3133;
input n_2002;
input n_581;
input n_2650;
input n_2138;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_2414;
input n_1340;
input n_3014;
input n_3166;
input n_1771;
input n_2316;
input n_3104;
input n_631;
input n_720;
input n_3435;
input n_153;
input n_842;
input n_3148;
input n_2262;
input n_3229;
input n_3348;
input n_1707;
input n_2239;
input n_3082;
input n_1432;
input n_156;
input n_145;
input n_2208;
input n_843;
input n_656;
input n_989;
input n_2604;
input n_2407;
input n_1277;
input n_2816;
input n_797;
input n_2689;
input n_2933;
input n_1473;
input n_2191;
input n_1723;
input n_2717;
input n_1246;
input n_1878;
input n_2574;
input n_899;
input n_189;
input n_738;
input n_2012;
input n_1304;
input n_1035;
input n_294;
input n_2842;
input n_499;
input n_2675;
input n_1426;
input n_3418;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_2134;
input n_1529;
input n_2335;
input n_2473;
input n_1022;
input n_614;
input n_529;
input n_2069;
input n_2307;
input n_2362;
input n_425;
input n_684;
input n_2539;
input n_2667;
input n_2698;
input n_1431;
input n_1615;
input n_1474;
input n_3312;
input n_1571;
input n_1809;
input n_3119;
input n_2948;
input n_1577;
input n_2958;
input n_2297;
input n_1181;
input n_2119;
input n_1822;
input n_37;
input n_486;
input n_947;
input n_2936;
input n_3224;
input n_1117;
input n_2489;
input n_1087;
input n_1448;
input n_3173;
input n_1992;
input n_648;
input n_657;
input n_1049;
input n_3223;
input n_2771;
input n_2445;
input n_3020;
input n_2057;
input n_2103;
input n_3140;
input n_3185;
input n_2605;
input n_1666;
input n_2772;
input n_1505;
input n_803;
input n_290;
input n_118;
input n_1717;
input n_926;
input n_1817;
input n_2449;
input n_927;
input n_2610;
input n_3129;
input n_1849;
input n_2848;
input n_919;
input n_2868;
input n_1698;
input n_478;
input n_2231;
input n_929;
input n_107;
input n_2520;
input n_1228;
input n_417;
input n_2857;
input n_446;
input n_89;
input n_1568;
input n_1490;
input n_2372;
input n_777;
input n_1299;
input n_272;
input n_2896;
input n_526;
input n_2718;
input n_3019;
input n_2639;
input n_1183;
input n_1436;
input n_2898;
input n_2251;
input n_1384;
input n_69;
input n_2494;
input n_2959;
input n_2501;
input n_3203;
input n_3325;
input n_2238;
input n_293;
input n_2368;
input n_53;
input n_458;
input n_1070;
input n_2403;
input n_3342;
input n_2837;
input n_998;
input n_16;
input n_717;
input n_3200;
input n_1665;
input n_18;
input n_3259;
input n_2524;
input n_154;
input n_3167;
input n_1383;
input n_2460;
input n_3390;
input n_1178;
input n_98;
input n_2127;
input n_1424;
input n_2338;
input n_3324;
input n_3341;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_3025;
input n_2137;
input n_1626;
input n_3191;
input n_1507;
input n_2482;
input n_184;
input n_552;
input n_2532;
input n_1358;
input n_1811;
input n_1388;
input n_3006;
input n_216;
input n_2481;
input n_912;
input n_1857;
input n_1519;
input n_2144;
input n_3056;
input n_745;
input n_1284;
input n_1604;
input n_2296;
input n_2424;
input n_3201;
input n_3447;
input n_1142;
input n_2849;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1774;
input n_2354;
input n_2682;
input n_3032;
input n_3103;
input n_2589;
input n_1395;
input n_2110;
input n_2199;
input n_2661;
input n_731;
input n_2877;
input n_1502;
input n_1659;
input n_1955;
input n_755;
input n_931;
input n_1021;
input n_3393;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_2442;
input n_312;
input n_1791;
input n_1368;
input n_66;
input n_3451;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_3331;
input n_1137;
input n_1897;
input n_2064;
input n_880;
input n_3072;
input n_3087;
input n_2053;
input n_2259;
input n_2121;
input n_2773;
input n_2545;
input n_889;
input n_2432;
input n_2710;
input n_150;
input n_1478;
input n_589;
input n_1310;
input n_3142;
input n_819;
input n_2966;
input n_2294;
input n_1363;
input n_2581;
input n_1334;
input n_1942;
input n_1966;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_1837;
input n_2218;
input n_2788;
input n_477;
input n_3196;
input n_2435;
input n_954;
input n_864;
input n_2504;
input n_2797;
input n_2623;
input n_1110;
input n_2213;
input n_1410;
input n_399;
input n_2389;
input n_1440;
input n_124;
input n_2132;
input n_2892;
input n_2063;
input n_1382;
input n_1534;
input n_1564;
input n_1736;
input n_211;
input n_2748;
input n_1483;
input n_1834;
input n_2331;
input n_1372;
input n_231;
input n_2292;
input n_2860;
input n_3327;
input n_2330;
input n_40;
input n_3441;
input n_1457;
input n_505;
input n_1719;
input n_319;
input n_1339;
input n_1787;
input n_2701;
input n_2475;
input n_537;
input n_2511;
input n_1993;
input n_2281;
input n_1427;
input n_311;
input n_2416;
input n_2745;
input n_2617;
input n_2776;
input n_1466;
input n_10;
input n_403;
input n_1919;
input n_1080;
input n_723;
input n_1877;
input n_3144;
input n_3211;
input n_3244;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1939;
input n_2030;
input n_1769;
input n_1220;
input n_2323;
input n_1893;
input n_556;
input n_2784;
input n_2209;
input n_2301;
input n_162;
input n_3287;
input n_2387;
input n_3322;
input n_1755;
input n_1602;
input n_2421;
input n_1136;
input n_3270;
input n_2618;
input n_2025;
input n_2357;
input n_2846;
input n_2464;
input n_3265;
input n_128;
input n_1125;
input n_970;
input n_3306;
input n_2488;
input n_2224;
input n_1980;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_2329;
input n_1092;
input n_2237;
input n_3026;
input n_441;
input n_221;
input n_1060;
input n_1951;
input n_2250;
input n_3090;
input n_444;
input n_3033;
input n_146;
input n_1252;
input n_1784;
input n_3311;
input n_1223;
input n_303;
input n_511;
input n_2990;
input n_193;
input n_1286;
input n_1773;
input n_1775;
input n_2115;
input n_2410;
input n_2552;
input n_1053;
input n_3302;
input n_2374;
input n_416;
input n_1681;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1783;
input n_1533;
input n_1597;
input n_2929;
input n_2780;
input n_3226;
input n_3323;
input n_3364;
input n_4;
input n_266;
input n_296;
input n_2596;
input n_2274;
input n_3163;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_1618;
input n_3407;
input n_217;
input n_518;
input n_1531;
input n_2828;
input n_1185;
input n_453;
input n_3425;
input n_215;
input n_2384;
input n_1745;
input n_914;
input n_759;
input n_3127;
input n_2724;
input n_1831;
input n_426;
input n_317;
input n_2585;
input n_2621;
input n_1653;
input n_2352;
input n_1679;
input n_1625;
input n_90;
input n_2601;
input n_2160;
input n_3454;
input n_54;
input n_1453;
input n_2146;
input n_2226;
input n_2131;
input n_488;
input n_2502;
input n_2801;
input n_497;
input n_2920;
input n_773;
input n_1901;
input n_920;
input n_99;
input n_1374;
input n_2556;
input n_2648;
input n_3212;
input n_1315;
input n_1647;
input n_13;
input n_2575;
input n_2754;
input n_1224;
input n_2783;
input n_2306;
input n_1614;
input n_1459;
input n_1892;
input n_3188;
input n_1933;
input n_2462;
input n_1135;
input n_1169;
input n_1179;
input n_2889;
input n_3243;
input n_401;
input n_324;
input n_1617;
input n_3260;
input n_3370;
input n_3386;
input n_335;
input n_1470;
input n_2550;
input n_463;
input n_3093;
input n_3175;
input n_3214;
input n_1243;
input n_848;
input n_120;
input n_2732;
input n_301;
input n_2928;
input n_274;
input n_1096;
input n_2249;
input n_1091;
input n_1917;
input n_2000;
input n_1580;
input n_2227;
input n_2270;
input n_2822;
input n_1425;
input n_3169;
input n_36;
input n_3205;
input n_1881;
input n_1267;
input n_1281;
input n_1806;
input n_3284;
input n_983;
input n_3109;
input n_2023;
input n_3354;
input n_427;
input n_2572;
input n_2204;
input n_1520;
input n_496;
input n_2720;
input n_3126;
input n_2159;
input n_906;
input n_1390;
input n_688;
input n_2289;
input n_1077;
input n_1733;
input n_2315;
input n_1419;
input n_2863;
input n_3299;
input n_351;
input n_2955;
input n_2995;
input n_259;
input n_1731;
input n_177;
input n_2158;
input n_2087;
input n_1855;
input n_1636;
input n_3051;
input n_1437;
input n_3360;
input n_2135;
input n_3367;
input n_1645;
input n_1832;
input n_385;
input n_1687;
input n_1439;
input n_2328;
input n_1323;
input n_2859;
input n_2202;
input n_858;
input n_2049;
input n_1331;
input n_613;
input n_736;
input n_2627;
input n_501;
input n_956;
input n_960;
input n_2276;
input n_3234;
input n_663;
input n_856;
input n_2803;
input n_2100;
input n_3314;
input n_379;
input n_2993;
input n_778;
input n_1668;
input n_2777;
input n_1134;
input n_3016;
input n_3004;
input n_3202;
input n_2830;
input n_2781;
input n_3220;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_1696;
input n_2829;
input n_1995;
input n_1594;
input n_2181;
input n_664;
input n_1869;
input n_171;
input n_2911;
input n_1764;
input n_169;
input n_1429;
input n_2826;
input n_1610;
input n_3084;
input n_3429;
input n_1889;
input n_2379;
input n_435;
input n_1905;
input n_2016;
input n_2343;
input n_793;
input n_326;
input n_587;
input n_1593;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_1937;
input n_465;
input n_1790;
input n_1778;
input n_1635;
input n_2942;
input n_1079;
input n_341;
input n_2515;
input n_1744;
input n_828;
input n_2139;
input n_2142;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_2448;
input n_1103;
input n_2875;
input n_2555;
input n_3338;
input n_144;
input n_3462;
input n_2219;
input n_1203;
input n_2851;
input n_3406;
input n_820;
input n_2327;
input n_951;
input n_106;
input n_2201;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_2841;
input n_3349;
input n_2420;
input n_186;
input n_2984;
input n_0;
input n_368;
input n_575;
input n_994;
input n_2263;
input n_3291;
input n_2304;
input n_1508;
input n_2487;
input n_732;
input n_974;
input n_2983;
input n_2240;
input n_392;
input n_2278;
input n_2656;
input n_2538;
input n_724;
input n_2597;
input n_2375;
input n_3113;
input n_3194;
input n_3250;
input n_1934;
input n_3276;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_1728;
input n_557;
input n_2756;
input n_1871;
input n_349;
input n_3448;
input n_617;
input n_845;
input n_807;
input n_2924;
input n_1036;
input n_140;
input n_1138;
input n_3414;
input n_1661;
input n_1275;
input n_2884;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_421;
input n_3120;
input n_1468;
input n_2855;
input n_1859;
input n_2102;
input n_2563;
input n_238;
input n_1095;
input n_2024;
input n_1595;
input n_202;
input n_2156;
input n_3449;
input n_1718;
input n_1749;
input n_1683;
input n_1916;
input n_2598;
input n_597;
input n_280;
input n_1270;
input n_2549;
input n_1187;
input n_610;
input n_1403;
input n_1669;
input n_1852;
input n_1024;
input n_1768;
input n_2153;
input n_2544;
input n_2381;
input n_198;
input n_1847;
input n_2052;
input n_179;
input n_248;
input n_2302;
input n_517;
input n_1667;
input n_667;
input n_1206;
input n_3230;
input n_621;
input n_1037;
input n_1397;
input n_3268;
input n_3236;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_468;
input n_2755;
input n_3141;
input n_923;
input n_504;
input n_1409;
input n_1841;
input n_2637;
input n_2823;
input n_1639;
input n_1623;
input n_183;
input n_1015;
input n_1503;
input n_3112;
input n_2819;
input n_3195;
input n_466;
input n_2526;
input n_3041;
input n_2423;
input n_1057;
input n_3277;
input n_3108;
input n_2548;
input n_603;
input n_991;
input n_2785;
input n_1657;
input n_235;
input n_1126;
input n_2412;
input n_1997;
input n_3417;
input n_2636;
input n_3131;
input n_340;
input n_710;
input n_1108;
input n_1818;
input n_2439;
input n_2404;
input n_1182;
input n_1298;
input n_2559;
input n_2177;
input n_39;
input n_2595;
input n_3399;
input n_2088;
input n_73;
input n_1611;
input n_785;
input n_2740;
input n_746;
input n_609;
input n_1601;
input n_3011;
input n_1960;
input n_2694;
input n_2061;
input n_3416;
input n_1686;
input n_2757;
input n_2337;
input n_2401;
input n_101;
input n_167;
input n_1356;
input n_1589;
input n_3042;
input n_3213;
input n_127;
input n_2309;
input n_2900;
input n_2957;
input n_2607;
input n_1740;
input n_2737;
input n_1497;
input n_2890;
input n_1168;
input n_1216;
input n_1943;
input n_3228;
input n_133;
input n_1320;
input n_2716;
input n_96;
input n_3249;
input n_3081;
input n_2452;
input n_1430;
input n_1316;
input n_1287;
input n_2722;
input n_1452;
input n_2854;
input n_3010;
input n_2499;
input n_3043;
input n_1622;
input n_1586;
input n_2543;
input n_2264;
input n_3464;
input n_302;
input n_1694;
input n_380;
input n_1535;
input n_3137;
input n_3382;
input n_2486;
input n_3132;
input n_137;
input n_2571;
input n_3138;
input n_1596;
input n_3177;
input n_20;
input n_1190;
input n_1734;
input n_3172;
input n_397;
input n_2902;
input n_3217;
input n_1983;
input n_1938;
input n_2498;
input n_122;
input n_2220;
input n_2577;
input n_34;
input n_1262;
input n_2472;
input n_218;
input n_1891;
input n_2171;
input n_1213;
input n_3238;
input n_70;
input n_2235;
input n_3394;
input n_2988;
input n_3136;
input n_1350;
input n_1673;
input n_2232;
input n_1715;
input n_172;
input n_1443;
input n_1272;
input n_2392;
input n_2894;
input n_3424;
input n_2790;
input n_239;
input n_2037;
input n_97;
input n_2808;
input n_2298;
input n_782;
input n_2326;
input n_1539;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_3040;
input n_1797;
input n_3279;
input n_1608;
input n_986;
input n_2305;
input n_2120;
input n_80;
input n_1472;
input n_2050;
input n_2373;
input n_2164;
input n_2402;
input n_2225;
input n_1081;
input n_402;
input n_1870;
input n_352;
input n_2964;
input n_1692;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_2169;
input n_2371;
input n_1827;
input n_1361;
input n_1864;
input n_2006;
input n_3402;
input n_1491;
input n_2187;
input n_662;
input n_374;
input n_1152;
input n_1840;
input n_1705;
input n_450;
input n_3262;
input n_2904;
input n_2244;
input n_3013;
input n_3356;
input n_2586;
input n_1684;
input n_921;
input n_2446;
input n_1346;
input n_711;
input n_1642;
input n_579;
input n_1352;
input n_2789;
input n_3105;
input n_3210;
input n_2872;
input n_937;
input n_2257;
input n_1682;
input n_2017;
input n_370;
input n_1695;
input n_1828;
input n_2046;
input n_2272;
input n_2699;
input n_2200;
input n_3029;
input n_650;
input n_1046;
input n_2560;
input n_1940;
input n_1979;
input n_2760;
input n_2704;
input n_3329;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_1963;
input n_2738;
input n_972;
input n_1405;
input n_2376;
input n_258;
input n_1406;
input n_456;
input n_2766;
input n_1332;
input n_260;
input n_2670;
input n_313;
input n_2700;
input n_624;
input n_962;
input n_1041;
input n_2346;
input n_565;
input n_3134;
input n_356;
input n_1569;
input n_936;
input n_3045;
input n_3115;
input n_1883;
input n_1288;
input n_3318;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_3278;
input n_2342;
input n_2167;
input n_2084;
input n_2970;
input n_2882;
input n_3320;
input n_2541;
input n_654;
input n_2940;
input n_411;
input n_2518;
input n_2458;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_1823;
input n_2479;
input n_3050;
input n_3350;
input n_105;
input n_2782;
input n_227;
input n_1974;
input n_2673;
input n_2456;
input n_1720;
input n_2527;
input n_204;
input n_482;
input n_934;
input n_1637;
input n_2635;
input n_3307;
input n_3439;
input n_1407;
input n_1795;
input n_2768;
input n_2871;
input n_420;
input n_2688;
input n_1341;
input n_394;
input n_1456;
input n_1845;
input n_1489;
input n_164;
input n_2314;
input n_23;
input n_942;
input n_3003;
input n_2798;
input n_2852;
input n_1524;
input n_543;
input n_2229;
input n_1964;
input n_2288;
input n_1920;
input n_2753;
input n_2099;
input n_1496;
input n_1271;
input n_3292;
input n_1545;
input n_2007;
input n_3121;
input n_2039;
input n_3388;
input n_1946;
input n_1355;
input n_1225;
input n_3184;
input n_1544;
input n_1485;
input n_2258;
input n_325;
input n_1640;
input n_804;
input n_464;
input n_1846;
input n_3437;
input n_3245;
input n_3075;
input n_2406;
input n_533;
input n_2390;
input n_806;
input n_879;
input n_959;
input n_2310;
input n_2506;
input n_584;
input n_2141;
input n_2562;
input n_244;
input n_2642;
input n_1343;
input n_1522;
input n_76;
input n_2734;
input n_548;
input n_1782;
input n_94;
input n_282;
input n_2383;
input n_2626;
input n_1676;
input n_833;
input n_1830;
input n_2351;
input n_1567;
input n_523;
input n_1319;
input n_707;
input n_2986;
input n_345;
input n_1900;
input n_3246;
input n_799;
input n_1548;
input n_3381;
input n_3044;
input n_2973;
input n_1155;
input n_2536;
input n_139;
input n_2196;
input n_41;
input n_2629;
input n_273;
input n_1633;
input n_2195;
input n_3208;
input n_2809;
input n_3007;
input n_787;
input n_2172;
input n_2835;
input n_1416;
input n_1528;
input n_2820;
input n_2293;
input n_1146;
input n_2021;
input n_3355;
input n_2454;
input n_2114;
input n_3074;
input n_3174;
input n_159;
input n_1086;
input n_1066;
input n_3102;
input n_1948;
input n_157;
input n_2125;
input n_2026;
input n_1282;
input n_2561;
input n_550;
input n_3321;
input n_2567;
input n_2322;
input n_275;
input n_652;
input n_2154;
input n_2727;
input n_2962;
input n_3377;
input n_2939;
input n_560;
input n_1906;
input n_1484;
input n_2992;
input n_3305;
input n_1241;
input n_1321;
input n_1672;
input n_569;
input n_2533;
input n_3157;
input n_1758;
input n_3221;
input n_3267;
input n_2283;
input n_2869;
input n_2422;
input n_1925;
input n_737;
input n_1318;
input n_1914;
input n_1235;
input n_3457;
input n_1229;
input n_2759;
input n_2945;
input n_3061;
input n_2361;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_2266;
input n_2960;
input n_3005;
input n_346;
input n_3;
input n_2427;
input n_3151;
input n_3411;
input n_1029;
input n_1447;
input n_2388;
input n_2056;
input n_790;
input n_2611;
input n_2901;
input n_138;
input n_3258;
input n_1706;
input n_3389;
input n_1498;
input n_3143;
input n_2653;
input n_2417;
input n_3000;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_2189;
input n_2680;
input n_2246;
input n_1047;
input n_3149;
input n_3375;
input n_1984;
input n_3365;
input n_2236;
input n_1385;
input n_431;
input n_3379;
input n_3156;
input n_24;
input n_459;
input n_1269;
input n_1931;
input n_2083;
input n_2834;
input n_3207;
input n_502;
input n_2668;
input n_672;
input n_2441;
input n_1257;
input n_3008;
input n_1751;
input n_3401;
input n_2840;
input n_3197;
input n_3242;
input n_285;
input n_1375;
input n_1941;
input n_85;
input n_2128;
input n_655;
input n_706;
input n_1045;
input n_1650;
input n_786;
input n_1794;
input n_1236;
input n_1962;
input n_1559;
input n_1725;
input n_1928;
input n_2398;
input n_1872;
input n_3091;
input n_834;
input n_19;
input n_29;
input n_2695;
input n_75;
input n_743;
input n_766;
input n_3124;
input n_430;
input n_1741;
input n_1325;
input n_1002;
input n_1746;
input n_1949;
input n_3398;
input n_545;
input n_2671;
input n_489;
input n_2761;
input n_2885;
input n_2793;
input n_2715;
input n_2888;
input n_1804;
input n_2923;
input n_1727;
input n_251;
input n_2508;
input n_1019;
input n_636;
input n_2054;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_2845;
input n_1337;
input n_3097;
input n_660;
input n_2062;
input n_2041;
input n_2975;
input n_438;
input n_1477;
input n_1360;
input n_2839;
input n_1860;
input n_2856;
input n_1904;
input n_2874;
input n_1200;
input n_2070;
input n_2588;
input n_479;
input n_1607;
input n_1353;
input n_1777;
input n_1908;
input n_1454;
input n_2484;
input n_2348;
input n_2944;
input n_2614;
input n_2126;
input n_869;
input n_1154;
input n_3308;
input n_1113;
input n_1600;
input n_2833;
input n_2253;
input n_2758;
input n_2366;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_2937;
input n_1329;
input n_2045;
input n_817;
input n_2261;
input n_2216;
input n_2210;
input n_262;
input n_187;
input n_897;
input n_846;
input n_3300;
input n_2978;
input n_2066;
input n_841;
input n_1476;
input n_2516;
input n_3391;
input n_1001;
input n_508;
input n_1800;
input n_2241;
input n_1050;
input n_1411;
input n_1463;
input n_2903;
input n_2827;
input n_1177;
input n_3216;
input n_3458;
input n_332;
input n_1150;
input n_1742;
input n_3190;
input n_1562;
input n_1690;
input n_398;
input n_1191;
input n_1826;
input n_566;
input n_1023;
input n_1882;
input n_2951;
input n_1076;
input n_1118;
input n_194;
input n_2949;
input n_57;
input n_1007;
input n_1807;
input n_1929;
input n_1378;
input n_2369;
input n_855;
input n_1592;
input n_1759;
input n_2719;
input n_1814;
input n_1631;
input n_52;
input n_591;
input n_1377;
input n_1879;
input n_256;
input n_853;
input n_440;
input n_695;
input n_1542;
input n_2587;
input n_3199;
input n_2931;
input n_875;
input n_209;
input n_367;
input n_680;
input n_3339;
input n_1678;
input n_2569;
input n_661;
input n_2400;
input n_1716;
input n_278;
input n_1256;
input n_671;
input n_1953;
input n_7;
input n_933;
input n_740;
input n_703;
input n_3343;
input n_3303;
input n_978;
input n_2752;
input n_384;
input n_3135;
input n_1976;
input n_2905;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_1824;
input n_310;
input n_1628;
input n_1324;
input n_1399;
input n_2122;
input n_2109;
input n_1435;
input n_969;
input n_988;
input n_2140;
input n_3160;
input n_1065;
input n_2796;
input n_3255;
input n_2507;
input n_84;
input n_1401;
input n_2358;
input n_1255;
input n_568;
input n_1516;
input n_143;
input n_1536;
input n_180;
input n_2163;
input n_2186;
input n_2029;
input n_2815;
input n_1204;
input n_3034;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_2528;
input n_2814;
input n_214;
input n_246;
input n_2787;
input n_1338;
input n_1097;
input n_2969;
input n_2395;
input n_935;
input n_3027;
input n_781;
input n_789;
input n_1554;
input n_3231;
input n_1130;
input n_3083;
input n_2979;
input n_181;
input n_1810;
input n_182;
input n_2953;
input n_573;
input n_769;
input n_2380;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_1583;
input n_3049;
input n_1730;
input n_2295;
input n_555;
input n_389;
input n_814;
input n_2746;
input n_2946;
input n_1643;
input n_2020;
input n_2500;
input n_3430;
input n_2269;
input n_1729;
input n_669;
input n_2290;
input n_2048;
input n_176;
input n_114;
input n_300;
input n_222;
input n_2005;
input n_747;
input n_74;
input n_2565;
input n_1389;
input n_1105;
input n_3117;
input n_721;
input n_1461;
input n_742;
input n_3432;
input n_535;
input n_691;
input n_372;
input n_2076;
input n_2736;
input n_111;
input n_2883;
input n_314;
input n_1408;
input n_378;
input n_1196;
input n_377;
input n_1598;
input n_2935;
input n_863;
input n_3015;
input n_2175;
input n_601;
input n_2182;
input n_338;
input n_2910;
input n_1283;
input n_2385;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_1785;
input n_56;
input n_763;
input n_1147;
input n_1848;
input n_360;
input n_1754;
input n_2149;
input n_3057;
input n_3154;
input n_2396;
input n_1506;
input n_119;
input n_2584;
input n_1652;
input n_1812;
input n_957;
input n_1994;
input n_895;
input n_866;
input n_1227;
input n_2450;
input n_2485;
input n_2284;
input n_191;
input n_2566;
input n_387;
input n_2287;
input n_452;
input n_744;
input n_971;
input n_2702;
input n_3241;
input n_946;
input n_344;
input n_2906;
input n_761;
input n_1303;
input n_2769;
input n_1205;
input n_2492;
input n_1258;
input n_2438;
input n_2914;
input n_1392;
input n_174;
input n_1173;
input n_1924;
input n_525;
input n_2463;
input n_3363;
input n_2881;
input n_1677;
input n_1116;
input n_611;
input n_1570;
input n_1702;
input n_1219;
input n_3064;
input n_1780;
input n_3100;
input n_1689;
input n_8;
input n_2180;
input n_3372;
input n_2858;
input n_3062;
input n_2679;
input n_1174;
input n_1944;
input n_1016;
input n_1347;
input n_795;
input n_1501;
input n_1221;
input n_3334;
input n_1245;
input n_838;
input n_3215;
input n_129;
input n_3336;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_2952;
input n_1017;
input n_3068;
input n_2117;
input n_2234;
input n_2779;
input n_2685;
input n_1083;
input n_109;
input n_445;
input n_1561;
input n_2741;
input n_3114;
input n_930;
input n_888;
input n_2275;
input n_1112;
input n_2465;
input n_2620;
input n_2081;
input n_2168;
input n_2568;
input n_234;
input n_2022;
input n_1945;
input n_2203;
input n_910;
input n_1656;
input n_1721;
input n_1460;
input n_911;
input n_2112;
input n_2255;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1737;
input n_2430;
input n_1414;
input n_752;
input n_908;
input n_2649;
input n_2721;
input n_944;
input n_2034;
input n_576;
input n_1028;
input n_2106;
input n_472;
input n_2862;
input n_270;
input n_2265;
input n_2615;
input n_414;
input n_2683;
input n_1922;
input n_563;
input n_2032;
input n_2744;
input n_1011;
input n_2474;
input n_1566;
input n_1215;
input n_2437;
input n_25;
input n_93;
input n_839;
input n_2444;
input n_2743;
input n_708;
input n_1973;
input n_3181;
input n_2267;
input n_3456;
input n_3035;
input n_668;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1821;
input n_2205;
input n_3204;
input n_1104;
input n_854;
input n_1058;
input n_3378;
input n_2312;
input n_498;
input n_3404;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_2242;
input n_3362;
input n_1509;
input n_103;
input n_3328;
input n_1693;
input n_2934;
input n_3290;
input n_1109;
input n_185;
input n_2222;
input n_712;
input n_3256;
input n_348;
input n_1276;
input n_3176;
input n_376;
input n_3309;
input n_2015;
input n_2118;
input n_2111;
input n_2466;
input n_390;
input n_2915;
input n_2530;
input n_1148;
input n_31;
input n_2188;
input n_2505;
input n_334;
input n_1989;
input n_1161;
input n_2609;
input n_1085;
input n_232;
input n_2802;
input n_2999;
input n_2014;
input n_2042;
input n_46;
input n_1239;
input n_771;
input n_1584;
input n_2425;
input n_470;
input n_475;
input n_924;
input n_3408;
input n_3461;
input n_298;
input n_1582;
input n_492;
input n_2318;
input n_3286;
input n_2408;
input n_1149;
input n_3170;
input n_265;
input n_1184;
input n_2483;
input n_2950;
input n_228;
input n_719;
input n_1972;
input n_3060;
input n_3304;
input n_2592;
input n_1525;
input n_3098;
input n_2594;
input n_455;
input n_2666;
input n_1585;
input n_1851;
input n_363;
input n_1799;
input n_1090;
input n_2147;
input n_2564;
input n_592;
input n_1816;
input n_2503;
input n_2433;
input n_1518;
input n_829;
input n_1156;
input n_1362;
input n_3123;
input n_393;
input n_984;
input n_2600;
input n_3380;
input n_1829;
input n_503;
input n_2035;
input n_3024;
input n_1450;
input n_1638;
input n_3422;
input n_132;
input n_868;
input n_3038;
input n_570;
input n_859;
input n_2033;
input n_406;
input n_3086;
input n_735;
input n_1789;
input n_2531;
input n_1770;
input n_878;
input n_620;
input n_130;
input n_3285;
input n_519;
input n_2523;
input n_307;
input n_469;
input n_1218;
input n_2413;
input n_500;
input n_1482;
input n_3361;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_2071;
input n_357;
input n_3219;
input n_2429;
input n_3130;
input n_985;
input n_2233;
input n_2440;
input n_2723;
input n_481;
input n_3233;
input n_997;
input n_1710;
input n_2800;
input n_2161;
input n_1301;
input n_2805;
input n_802;
input n_561;
input n_33;
input n_3310;
input n_980;
input n_2681;
input n_1306;
input n_3264;
input n_2010;
input n_2282;
input n_1651;
input n_1198;
input n_3096;
input n_2360;
input n_2047;
input n_2651;
input n_2095;
input n_3239;
input n_1609;
input n_2174;
input n_3161;
input n_2799;
input n_436;
input n_116;
input n_3344;
input n_2334;
input n_3295;
input n_409;
input n_1244;
input n_1685;
input n_1763;
input n_1998;
input n_3066;
input n_1574;
input n_2426;
input n_2490;
input n_2844;
input n_3101;
input n_240;
input n_756;
input n_2303;
input n_1619;
input n_2478;
input n_1981;
input n_2285;
input n_1606;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_3374;
input n_2742;
input n_2640;
input n_1051;
input n_253;
input n_1552;
input n_2918;
input n_583;
input n_3288;
input n_1996;
input n_2367;
input n_249;
input n_201;
input n_2867;
input n_3198;
input n_1039;
input n_1442;
input n_2726;
input n_1034;
input n_2043;
input n_1480;
input n_3125;
input n_1158;
input n_2909;
input n_2248;
input n_754;
input n_941;
input n_975;
input n_3206;
input n_1031;
input n_115;
input n_1305;
input n_2363;
input n_2578;
input n_553;
input n_43;
input n_849;
input n_2662;
input n_3116;
input n_3147;
input n_3383;
input n_753;
input n_1753;
input n_3095;
input n_3180;
input n_3359;
input n_2795;
input n_2471;
input n_467;
input n_3187;
input n_2540;
input n_269;
input n_359;
input n_973;
input n_2807;
input n_1921;
input n_3218;
input n_3330;
input n_1479;
input n_1055;
input n_1675;
input n_2197;
input n_2217;
input n_582;
input n_2065;
input n_2879;
input n_861;
input n_857;
input n_967;
input n_571;
input n_2215;
input n_2461;
input n_271;
input n_404;
input n_2001;
input n_158;
input n_2107;
input n_1884;
input n_206;
input n_2040;
input n_679;
input n_2968;
input n_633;
input n_1170;
input n_665;
input n_1629;
input n_2221;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1819;
input n_2055;
input n_1010;
input n_3444;
input n_2553;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_3059;
input n_1166;
input n_2038;
input n_812;
input n_2891;
input n_1131;
input n_2634;
input n_1761;
input n_2709;
input n_3155;
input n_3445;
input n_534;
input n_1578;
input n_1006;
input n_1861;
input n_373;
input n_3110;
input n_87;
input n_1632;
input n_1890;
input n_3017;
input n_1805;
input n_2477;
input n_257;
input n_1557;
input n_1888;
input n_2280;
input n_1833;
input n_730;
input n_1311;
input n_1494;
input n_2325;
input n_670;
input n_203;
input n_1850;
input n_1898;
input n_2443;
input n_2697;
input n_3235;
input n_2308;
input n_2162;
input n_1868;
input n_207;
input n_2333;
input n_2079;
input n_3001;
input n_1089;
input n_1887;
input n_1587;
input n_2512;
input n_3433;
input n_1365;
input n_1417;
input n_205;
input n_1242;
input n_2086;
input n_2185;
input n_2927;
input n_1836;
input n_2774;
input n_3039;
input n_681;
input n_1226;
input n_3162;
input n_1274;
input n_1486;
input n_2166;
input n_3094;
input n_412;
input n_2899;
input n_3274;
input n_3333;
input n_3186;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_1899;
input n_1428;
input n_1616;
input n_1576;
input n_1856;
input n_1862;
input n_1958;
input n_2077;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_3065;
input n_2632;
input n_422;
input n_2579;
input n_722;
input n_862;
input n_2105;
input n_135;
input n_3079;
input n_165;
input n_2098;
input n_3085;
input n_540;
input n_1423;
input n_2813;
input n_1935;
input n_3387;
input n_2027;
input n_457;
input n_3070;
input n_2223;
input n_2091;
input n_364;
input n_3263;
input n_3420;
input n_2991;
input n_1915;
input n_629;
input n_1621;
input n_1748;
input n_2547;
input n_2415;
input n_900;
input n_1449;
input n_531;
input n_827;
input n_2912;
input n_60;
input n_361;
input n_2659;
input n_2930;
input n_1025;
input n_3409;
input n_2419;
input n_3111;
input n_2116;
input n_336;
input n_2320;
input n_12;
input n_1885;
input n_2677;
input n_1013;
input n_3182;
input n_1259;
input n_3054;
input n_3283;
input n_192;
input n_2183;
input n_3002;
input n_1538;
input n_51;
input n_649;
input n_1612;
input n_1240;

output n_14691;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_14428;
wire n_13611;
wire n_6566;
wire n_4452;
wire n_13045;
wire n_5172;
wire n_11173;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_6872;
wire n_13998;
wire n_5254;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_13146;
wire n_13235;
wire n_10587;
wire n_5019;
wire n_8713;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_3849;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_5138;
wire n_13522;
wire n_10931;
wire n_4395;
wire n_6960;
wire n_4388;
wire n_8169;
wire n_12265;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_7180;
wire n_5653;
wire n_11574;
wire n_4978;
wire n_13530;
wire n_8604;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_13125;
wire n_8168;
wire n_4829;
wire n_5393;
wire n_7190;
wire n_7504;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_4686;
wire n_12322;
wire n_14318;
wire n_8899;
wire n_14196;
wire n_5524;
wire n_10236;
wire n_5345;
wire n_11205;
wire n_11776;
wire n_11678;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_11650;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_8534;
wire n_5963;
wire n_12179;
wire n_13942;
wire n_5055;
wire n_14439;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_11905;
wire n_4868;
wire n_10020;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_4249;
wire n_11536;
wire n_5950;
wire n_3564;
wire n_9104;
wire n_6999;
wire n_11046;
wire n_11079;
wire n_10283;
wire n_5548;
wire n_5057;
wire n_11065;
wire n_8339;
wire n_8272;
wire n_14215;
wire n_13997;
wire n_14402;
wire n_7161;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_13437;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_11214;
wire n_5101;
wire n_7000;
wire n_8561;
wire n_11954;
wire n_7398;
wire n_14232;
wire n_10392;
wire n_14341;
wire n_12882;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_12617;
wire n_8411;
wire n_8499;
wire n_8236;
wire n_5102;
wire n_13137;
wire n_13221;
wire n_6882;
wire n_10775;
wire n_4501;
wire n_9626;
wire n_11163;
wire n_9526;
wire n_13657;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_14099;
wire n_5598;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_7389;
wire n_4997;
wire n_10719;
wire n_11419;
wire n_9018;
wire n_4843;
wire n_12095;
wire n_8070;
wire n_13663;
wire n_13990;
wire n_4696;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_11740;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_13993;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_7008;
wire n_3877;
wire n_12392;
wire n_3929;
wire n_8366;
wire n_8102;
wire n_9362;
wire n_11979;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_5894;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_9962;
wire n_5908;
wire n_3979;
wire n_4814;
wire n_10373;
wire n_11104;
wire n_8913;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_4956;
wire n_11537;
wire n_13814;
wire n_12707;
wire n_7686;
wire n_3664;
wire n_6914;
wire n_10335;
wire n_5337;
wire n_5129;
wire n_11301;
wire n_12424;
wire n_13681;
wire n_14121;
wire n_5420;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_4414;
wire n_6585;
wire n_11703;
wire n_11699;
wire n_6374;
wire n_4646;
wire n_7651;
wire n_11543;
wire n_10947;
wire n_6628;
wire n_8125;
wire n_13483;
wire n_3760;
wire n_6015;
wire n_14662;
wire n_11261;
wire n_10226;
wire n_13247;
wire n_4262;
wire n_6526;
wire n_13929;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_10767;
wire n_5136;
wire n_8040;
wire n_14646;
wire n_11821;
wire n_14095;
wire n_5638;
wire n_13121;
wire n_13989;
wire n_9100;
wire n_4110;
wire n_6784;
wire n_12107;
wire n_14520;
wire n_10755;
wire n_4950;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_6323;
wire n_9614;
wire n_14431;
wire n_13515;
wire n_10682;
wire n_6110;
wire n_11684;
wire n_3999;
wire n_12652;
wire n_3928;
wire n_6371;
wire n_14410;
wire n_8079;
wire n_10699;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_9400;
wire n_5151;
wire n_8142;
wire n_11627;
wire n_5684;
wire n_8598;
wire n_13139;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_13803;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_14066;
wire n_7856;
wire n_7774;
wire n_5680;
wire n_6674;
wire n_13606;
wire n_6148;
wire n_6951;
wire n_11659;
wire n_7625;
wire n_13501;
wire n_4102;
wire n_3871;
wire n_9106;
wire n_13509;
wire n_12775;
wire n_13729;
wire n_4662;
wire n_8869;
wire n_6989;
wire n_7863;
wire n_4671;
wire n_3959;
wire n_8381;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_9520;
wire n_8958;
wire n_14485;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_14628;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_13687;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_12371;
wire n_4296;
wire n_10114;
wire n_12203;
wire n_10357;
wire n_14540;
wire n_7147;
wire n_8115;
wire n_4507;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_11497;
wire n_3484;
wire n_12359;
wire n_4677;
wire n_12915;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_13149;
wire n_13711;
wire n_13454;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_12742;
wire n_3923;
wire n_14091;
wire n_9042;
wire n_11768;
wire n_3900;
wire n_8412;
wire n_9267;
wire n_3488;
wire n_3732;
wire n_6485;
wire n_8987;
wire n_11805;
wire n_14461;
wire n_14478;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_4226;
wire n_5493;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_13958;
wire n_3980;
wire n_5346;
wire n_5252;
wire n_4366;
wire n_5309;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_12770;
wire n_10012;
wire n_14570;
wire n_4294;
wire n_13754;
wire n_12985;
wire n_4698;
wire n_13797;
wire n_4445;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_7564;
wire n_11635;
wire n_3859;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_14171;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_8119;
wire n_10296;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_9718;
wire n_9128;
wire n_10281;
wire n_13344;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_14380;
wire n_8748;
wire n_3927;
wire n_13984;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_14239;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_8718;
wire n_7110;
wire n_5476;
wire n_12831;
wire n_13920;
wire n_9935;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_14045;
wire n_14288;
wire n_8223;
wire n_3882;
wire n_4856;
wire n_10097;
wire n_3492;
wire n_4369;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_4331;
wire n_7297;
wire n_10018;
wire n_9866;
wire n_4972;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_12427;
wire n_7533;
wire n_14162;
wire n_13771;
wire n_7221;
wire n_4375;
wire n_13977;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_11295;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_11662;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_8246;
wire n_8952;
wire n_4613;
wire n_13014;
wire n_9070;
wire n_11708;
wire n_3875;
wire n_10266;
wire n_14401;
wire n_5609;
wire n_4717;
wire n_10827;
wire n_10897;
wire n_4877;
wire n_5922;
wire n_10449;
wire n_7569;
wire n_7823;
wire n_7734;
wire n_7062;
wire n_7861;
wire n_8955;
wire n_9680;
wire n_5658;
wire n_4731;
wire n_9477;
wire n_12172;
wire n_12147;
wire n_12923;
wire n_7039;
wire n_8577;
wire n_12384;
wire n_11349;
wire n_8594;
wire n_5046;
wire n_13227;
wire n_8428;
wire n_9829;
wire n_11260;
wire n_8848;
wire n_12825;
wire n_13341;
wire n_5058;
wire n_10685;
wire n_11351;
wire n_4467;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_5667;
wire n_8259;
wire n_12540;
wire n_10607;
wire n_14388;
wire n_5865;
wire n_12249;
wire n_8349;
wire n_6836;
wire n_5305;
wire n_5042;
wire n_11998;
wire n_4681;
wire n_8164;
wire n_13239;
wire n_4072;
wire n_10628;
wire n_4752;
wire n_4220;
wire n_13429;
wire n_7905;
wire n_5281;
wire n_8776;
wire n_11775;
wire n_9143;
wire n_8287;
wire n_10256;
wire n_10769;
wire n_7753;
wire n_10368;
wire n_6771;
wire n_7950;
wire n_9947;
wire n_13999;
wire n_9088;
wire n_8607;
wire n_14037;
wire n_10138;
wire n_12117;
wire n_11706;
wire n_6248;
wire n_11800;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_10452;
wire n_11464;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_12960;
wire n_14094;
wire n_13033;
wire n_11642;
wire n_4381;
wire n_11143;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_3968;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_12131;
wire n_6776;
wire n_4510;
wire n_12851;
wire n_5795;
wire n_11934;
wire n_12349;
wire n_6043;
wire n_4473;
wire n_5552;
wire n_7452;
wire n_14282;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_13550;
wire n_14217;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_13348;
wire n_8416;
wire n_10396;
wire n_13919;
wire n_4518;
wire n_10724;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_14062;
wire n_9988;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_14167;
wire n_12740;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_10363;
wire n_13240;
wire n_8949;
wire n_10831;
wire n_3500;
wire n_3834;
wire n_9131;
wire n_11553;
wire n_10517;
wire n_12578;
wire n_12795;
wire n_4589;
wire n_10323;
wire n_12194;
wire n_13623;
wire n_10842;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_10876;
wire n_11511;
wire n_9137;
wire n_11180;
wire n_14043;
wire n_9724;
wire n_11146;
wire n_9281;
wire n_10883;
wire n_8995;
wire n_10101;
wire n_9393;
wire n_4394;
wire n_6581;
wire n_13845;
wire n_12709;
wire n_6010;
wire n_13432;
wire n_8711;
wire n_7013;
wire n_12771;
wire n_14150;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_3696;
wire n_4082;
wire n_7290;
wire n_12278;
wire n_13721;
wire n_10820;
wire n_13514;
wire n_4921;
wire n_9687;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_7315;
wire n_13194;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_4697;
wire n_13244;
wire n_4289;
wire n_4288;
wire n_11866;
wire n_3763;
wire n_6185;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_9102;
wire n_11526;
wire n_13404;
wire n_9578;
wire n_3614;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_7438;
wire n_14355;
wire n_14128;
wire n_7268;
wire n_7337;
wire n_11851;
wire n_4964;
wire n_9489;
wire n_12804;
wire n_14123;
wire n_5957;
wire n_6965;
wire n_12116;
wire n_10728;
wire n_4228;
wire n_6357;
wire n_9144;
wire n_10094;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_14126;
wire n_14105;
wire n_7461;
wire n_8285;
wire n_13870;
wire n_4322;
wire n_10655;
wire n_13791;
wire n_3644;
wire n_9797;
wire n_6955;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_4287;
wire n_4137;
wire n_9521;
wire n_8332;
wire n_9478;
wire n_9932;
wire n_13040;
wire n_7278;
wire n_6509;
wire n_11370;
wire n_13900;
wire n_4576;
wire n_7454;
wire n_11253;
wire n_14652;
wire n_11379;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_11981;
wire n_9895;
wire n_8741;
wire n_12918;
wire n_4000;
wire n_9351;
wire n_11585;
wire n_5445;
wire n_13140;
wire n_13962;
wire n_14556;
wire n_5501;
wire n_5342;
wire n_6839;
wire n_3970;
wire n_7232;
wire n_7377;
wire n_4345;
wire n_4389;
wire n_13753;
wire n_6646;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_9189;
wire n_4664;
wire n_13716;
wire n_4156;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_14391;
wire n_7904;
wire n_11691;
wire n_6033;
wire n_11541;
wire n_13610;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_13332;
wire n_5748;
wire n_14408;
wire n_3782;
wire n_9356;
wire n_12865;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_3700;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_5636;
wire n_7840;
wire n_10972;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_13213;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_8800;
wire n_13385;
wire n_10845;
wire n_7080;
wire n_6636;
wire n_5286;
wire n_8229;
wire n_4528;
wire n_8410;
wire n_5811;
wire n_14156;
wire n_13992;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_7624;
wire n_4914;
wire n_4939;
wire n_7629;
wire n_13790;
wire n_14384;
wire n_9735;
wire n_9186;
wire n_10818;
wire n_5530;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_12552;
wire n_13304;
wire n_14633;
wire n_11069;
wire n_4096;
wire n_5595;
wire n_4123;
wire n_9941;
wire n_12222;
wire n_11951;
wire n_7003;
wire n_11900;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_3735;
wire n_11369;
wire n_4379;
wire n_10563;
wire n_14210;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_5901;
wire n_13362;
wire n_6538;
wire n_14373;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_7010;
wire n_8107;
wire n_11108;
wire n_9728;
wire n_12883;
wire n_11004;
wire n_12992;
wire n_5324;
wire n_6519;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_3770;
wire n_9818;
wire n_6530;
wire n_7219;
wire n_9662;
wire n_14154;
wire n_12896;
wire n_4440;
wire n_8774;
wire n_4402;
wire n_14518;
wire n_10566;
wire n_13397;
wire n_10178;
wire n_5052;
wire n_7299;
wire n_12367;
wire n_4541;
wire n_12104;
wire n_5009;
wire n_4872;
wire n_6402;
wire n_12469;
wire n_13526;
wire n_9936;
wire n_12563;
wire n_4551;
wire n_6195;
wire n_13132;
wire n_7326;
wire n_6609;
wire n_7243;
wire n_9530;
wire n_10115;
wire n_13321;
wire n_5326;
wire n_7471;
wire n_7067;
wire n_10455;
wire n_11778;
wire n_12793;
wire n_13427;
wire n_4627;
wire n_4079;
wire n_5300;
wire n_9909;
wire n_11393;
wire n_8620;
wire n_8691;
wire n_12406;
wire n_6748;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_13270;
wire n_7790;
wire n_11719;
wire n_6149;
wire n_10052;
wire n_10109;
wire n_7484;
wire n_3656;
wire n_7002;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_11963;
wire n_12428;
wire n_14636;
wire n_8424;
wire n_9571;
wire n_8026;
wire n_7528;
wire n_9470;
wire n_9638;
wire n_4798;
wire n_3810;
wire n_10265;
wire n_8174;
wire n_12655;
wire n_7941;
wire n_13524;
wire n_11175;
wire n_13792;
wire n_5010;
wire n_11483;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_14378;
wire n_5089;
wire n_13356;
wire n_11371;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_6264;
wire n_14191;
wire n_8861;
wire n_5359;
wire n_13480;
wire n_8644;
wire n_8907;
wire n_12304;
wire n_13571;
wire n_11080;
wire n_10984;
wire n_5137;
wire n_6902;
wire n_5104;
wire n_14079;
wire n_10100;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7478;
wire n_7913;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_3606;
wire n_12692;
wire n_13600;
wire n_13715;
wire n_3591;
wire n_7939;
wire n_13602;
wire n_14224;
wire n_8503;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_6449;
wire n_6723;
wire n_7458;
wire n_9108;
wire n_9787;
wire n_6440;
wire n_7436;
wire n_10846;
wire n_4746;
wire n_13363;
wire n_14101;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_8446;
wire n_5194;
wire n_9376;
wire n_9786;
wire n_14682;
wire n_9033;
wire n_13810;
wire n_14403;
wire n_12933;
wire n_7435;
wire n_12908;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_3534;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_13893;
wire n_3964;
wire n_12996;
wire n_14201;
wire n_5947;
wire n_8923;
wire n_13625;
wire n_12643;
wire n_13315;
wire n_13473;
wire n_6124;
wire n_6736;
wire n_3944;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_14597;
wire n_5985;
wire n_8197;
wire n_14353;
wire n_3605;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_12827;
wire n_12678;
wire n_13795;
wire n_9115;
wire n_12235;
wire n_14547;
wire n_4584;
wire n_5232;
wire n_11833;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_3847;
wire n_14386;
wire n_5001;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_9938;
wire n_11285;
wire n_8082;
wire n_12098;
wire n_4428;
wire n_8730;
wire n_7917;
wire n_7261;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_9203;
wire n_14415;
wire n_9977;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_5761;
wire n_13982;
wire n_13475;
wire n_9242;
wire n_6773;
wire n_4618;
wire n_12611;
wire n_13859;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_4679;
wire n_13569;
wire n_3479;
wire n_11262;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_12713;
wire n_12880;
wire n_13144;
wire n_4805;
wire n_8651;
wire n_13959;
wire n_9141;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_6531;
wire n_10952;
wire n_10851;
wire n_11027;
wire n_13628;
wire n_11852;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_10221;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_11803;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_13685;
wire n_5100;
wire n_9286;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_8281;
wire n_10819;
wire n_3816;
wire n_4807;
wire n_8842;
wire n_4411;
wire n_14521;
wire n_9184;
wire n_9704;
wire n_13585;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_14486;
wire n_8024;
wire n_7730;
wire n_12562;
wire n_8814;
wire n_8530;
wire n_11428;
wire n_11592;
wire n_4180;
wire n_9193;
wire n_8467;
wire n_11677;
wire n_7281;
wire n_9717;
wire n_13577;
wire n_7711;
wire n_11090;
wire n_8984;
wire n_3663;
wire n_5688;
wire n_6417;
wire n_9290;
wire n_13281;
wire n_5740;
wire n_5820;
wire n_13769;
wire n_5648;
wire n_13266;
wire n_13957;
wire n_14580;
wire n_5745;
wire n_4707;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_13672;
wire n_14028;
wire n_9875;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_8676;
wire n_5534;
wire n_8003;
wire n_4880;
wire n_13827;
wire n_8785;
wire n_9853;
wire n_13192;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_4126;
wire n_14542;
wire n_3845;
wire n_6556;
wire n_8692;
wire n_6889;
wire n_7230;
wire n_9183;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_9778;
wire n_14326;
wire n_5196;
wire n_6199;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_10852;
wire n_4470;
wire n_14665;
wire n_6726;
wire n_12374;
wire n_13200;
wire n_9529;
wire n_4813;
wire n_5542;
wire n_3901;
wire n_7011;
wire n_8998;
wire n_10538;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_4014;
wire n_13342;
wire n_4704;
wire n_11066;
wire n_10315;
wire n_4252;
wire n_13886;
wire n_9123;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_4048;
wire n_4596;
wire n_12368;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_13193;
wire n_6100;
wire n_12796;
wire n_6516;
wire n_3919;
wire n_14489;
wire n_8462;
wire n_13774;
wire n_6977;
wire n_9380;
wire n_13847;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_12529;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_6522;
wire n_8979;
wire n_14053;
wire n_4952;
wire n_5023;
wire n_5906;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_14581;
wire n_5660;
wire n_3981;
wire n_7890;
wire n_12785;
wire n_3973;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_14155;
wire n_12461;
wire n_6808;
wire n_13603;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_6207;
wire n_6931;
wire n_7006;
wire n_5821;
wire n_14160;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_9082;
wire n_10925;
wire n_4770;
wire n_9879;
wire n_11158;
wire n_3474;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_4690;
wire n_11669;
wire n_14390;
wire n_3864;
wire n_8264;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_12078;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_8135;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_3592;
wire n_11739;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_10497;
wire n_14561;
wire n_9445;
wire n_7627;
wire n_13301;
wire n_9803;
wire n_13293;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_6346;
wire n_14381;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_8408;
wire n_12639;
wire n_14212;
wire n_5386;
wire n_10661;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_3817;
wire n_10028;
wire n_13878;
wire n_7811;
wire n_13158;
wire n_14649;
wire n_11676;
wire n_11044;
wire n_11771;
wire n_12266;
wire n_3659;
wire n_12175;
wire n_5003;
wire n_13536;
wire n_10512;
wire n_13833;
wire n_11384;
wire n_4827;
wire n_12287;
wire n_11679;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_12353;
wire n_14441;
wire n_14129;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_12398;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_13485;
wire n_9087;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_9043;
wire n_6075;
wire n_12991;
wire n_3657;
wire n_7397;
wire n_10789;
wire n_11134;
wire n_12705;
wire n_13735;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_11828;
wire n_14470;
wire n_12326;
wire n_14264;
wire n_7847;
wire n_8506;
wire n_14115;
wire n_6494;
wire n_13830;
wire n_13178;
wire n_6133;
wire n_3723;
wire n_11548;
wire n_13041;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_14184;
wire n_7822;
wire n_6453;
wire n_4380;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_6127;
wire n_14183;
wire n_10762;
wire n_11452;
wire n_4398;
wire n_11342;
wire n_11362;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_14200;
wire n_5031;
wire n_6006;
wire n_10797;
wire n_11266;
wire n_7289;
wire n_4193;
wire n_3570;
wire n_14110;
wire n_12309;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_5338;
wire n_3828;
wire n_12479;
wire n_7354;
wire n_8352;
wire n_12502;
wire n_13824;
wire n_4131;
wire n_10360;
wire n_7960;
wire n_9450;
wire n_3594;
wire n_5689;
wire n_13953;
wire n_7482;
wire n_12912;
wire n_10312;
wire n_4090;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_9223;
wire n_13191;
wire n_6048;
wire n_6416;
wire n_4144;
wire n_10131;
wire n_12537;
wire n_6838;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_11988;
wire n_12600;
wire n_12921;
wire n_14536;
wire n_13226;
wire n_3485;
wire n_5931;
wire n_6139;
wire n_4077;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_13686;
wire n_6256;
wire n_7965;
wire n_13645;
wire n_6613;
wire n_11438;
wire n_11244;
wire n_4008;
wire n_12919;
wire n_14432;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_6361;
wire n_9880;
wire n_13253;
wire n_4689;
wire n_14321;
wire n_8183;
wire n_11348;
wire n_4547;
wire n_11245;
wire n_9685;
wire n_6085;
wire n_7474;
wire n_11169;
wire n_11685;
wire n_5731;
wire n_12422;
wire n_6329;
wire n_11607;
wire n_8650;
wire n_6678;
wire n_11546;
wire n_14654;
wire n_8662;
wire n_10503;
wire n_14422;
wire n_9694;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_14664;
wire n_13215;
wire n_13400;
wire n_4601;
wire n_9905;
wire n_9948;
wire n_10465;
wire n_14630;
wire n_12429;
wire n_10590;
wire n_3647;
wire n_3681;
wire n_13782;
wire n_14494;
wire n_4300;
wire n_8526;
wire n_13331;
wire n_4623;
wire n_7325;
wire n_13751;
wire n_10887;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_14019;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_5883;
wire n_13743;
wire n_7166;
wire n_13812;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_13378;
wire n_3988;
wire n_6560;
wire n_14055;
wire n_11319;
wire n_3476;
wire n_7028;
wire n_7838;
wire n_4842;
wire n_9890;
wire n_5629;
wire n_11492;
wire n_4135;
wire n_7873;
wire n_6535;
wire n_12731;
wire n_12399;
wire n_7518;
wire n_12342;
wire n_12640;
wire n_7414;
wire n_9744;
wire n_9817;
wire n_6147;
wire n_10063;
wire n_9199;
wire n_13092;
wire n_11160;
wire n_9548;
wire n_8973;
wire n_6448;
wire n_13544;
wire n_7791;
wire n_14292;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_12533;
wire n_9862;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_12616;
wire n_11385;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_12535;
wire n_12178;
wire n_4111;
wire n_14375;
wire n_12653;
wire n_6643;
wire n_12327;
wire n_7146;
wire n_9471;
wire n_4608;
wire n_3712;
wire n_11346;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_9069;
wire n_13110;
wire n_3562;
wire n_5852;
wire n_14030;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_8249;
wire n_7052;
wire n_11343;
wire n_12348;
wire n_3665;
wire n_10496;
wire n_12257;
wire n_3528;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_14149;
wire n_13394;
wire n_4571;
wire n_10843;
wire n_13391;
wire n_3698;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_13384;
wire n_14680;
wire n_8234;
wire n_5321;
wire n_9960;
wire n_10997;
wire n_4215;
wire n_9010;
wire n_13707;
wire n_10998;
wire n_9003;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_12418;
wire n_14216;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_13498;
wire n_3752;
wire n_7312;
wire n_13263;
wire n_7919;
wire n_5145;
wire n_4219;
wire n_11269;
wire n_10800;
wire n_7085;
wire n_11491;
wire n_12065;
wire n_3958;
wire n_13950;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_11408;
wire n_14048;
wire n_3985;
wire n_11772;
wire n_4196;
wire n_14103;
wire n_4774;
wire n_5210;
wire n_13183;
wire n_6689;
wire n_13732;
wire n_10993;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_12519;
wire n_9172;
wire n_12769;
wire n_14653;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_5149;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_11311;
wire n_10112;
wire n_14443;
wire n_10765;
wire n_3899;
wire n_6698;
wire n_11792;
wire n_14285;
wire n_7304;
wire n_3713;
wire n_9734;
wire n_7288;
wire n_8558;
wire n_13242;
wire n_10489;
wire n_7707;
wire n_7223;
wire n_12421;
wire n_13282;
wire n_14436;
wire n_7833;
wire n_12113;
wire n_4987;
wire n_14599;
wire n_5512;
wire n_7274;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_4736;
wire n_14351;
wire n_3743;
wire n_6206;
wire n_9068;
wire n_13352;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_10612;
wire n_11086;
wire n_7466;
wire n_6529;
wire n_10260;
wire n_11293;
wire n_3759;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_12285;
wire n_13310;
wire n_11710;
wire n_8619;
wire n_11568;
wire n_3511;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_9150;
wire n_10134;
wire n_14508;
wire n_11603;
wire n_13798;
wire n_7277;
wire n_6455;
wire n_13804;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_13099;
wire n_12015;
wire n_8146;
wire n_4492;
wire n_13690;
wire n_8813;
wire n_5607;
wire n_11562;
wire n_3694;
wire n_7695;
wire n_10194;
wire n_14566;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_12157;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_13386;
wire n_13846;
wire n_8910;
wire n_12311;
wire n_6203;
wire n_4376;
wire n_6408;
wire n_14374;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_13064;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_4708;
wire n_13619;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_12031;
wire n_5341;
wire n_8643;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_11718;
wire n_8565;
wire n_10821;
wire n_13648;
wire n_11170;
wire n_11758;
wire n_12126;
wire n_14383;
wire n_8550;
wire n_14543;
wire n_4081;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_14450;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_14683;
wire n_10599;
wire n_9667;
wire n_14192;
wire n_14181;
wire n_6401;
wire n_7322;
wire n_9053;
wire n_11658;
wire n_11893;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_13492;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_14001;
wire n_14213;
wire n_5562;
wire n_7051;
wire n_4324;
wire n_10850;
wire n_9185;
wire n_8477;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_4382;
wire n_12195;
wire n_13376;
wire n_13115;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_13864;
wire n_5911;
wire n_3954;
wire n_11601;
wire n_13289;
wire n_11971;
wire n_13182;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_5622;
wire n_3503;
wire n_9919;
wire n_12135;
wire n_6574;
wire n_11116;
wire n_13324;
wire n_12604;
wire n_6571;
wire n_13305;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_8876;
wire n_5124;
wire n_9151;
wire n_3951;
wire n_8829;
wire n_9359;
wire n_7824;
wire n_13381;
wire n_13236;
wire n_3569;
wire n_14189;
wire n_14299;
wire n_7094;
wire n_3874;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8140;
wire n_8971;
wire n_8060;
wire n_10558;
wire n_4083;
wire n_7036;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_6392;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_13777;
wire n_9049;
wire n_7351;
wire n_13718;
wire n_4480;
wire n_9352;
wire n_7608;
wire n_5779;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_13202;
wire n_7909;
wire n_7413;
wire n_13638;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_14392;
wire n_11340;
wire n_10734;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_11903;
wire n_7027;
wire n_7992;
wire n_13279;
wire n_13644;
wire n_6912;
wire n_11560;
wire n_10330;
wire n_10395;
wire n_7175;
wire n_8276;
wire n_3617;
wire n_13291;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_3567;
wire n_11465;
wire n_7524;
wire n_4344;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_11564;
wire n_14015;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_11265;
wire n_9370;
wire n_11125;
wire n_9670;
wire n_13136;
wire n_13513;
wire n_4027;
wire n_12916;
wire n_9334;
wire n_7783;
wire n_13220;
wire n_6692;
wire n_3898;
wire n_10276;
wire n_14322;
wire n_12331;
wire n_3520;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_12531;
wire n_8245;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_12521;
wire n_11302;
wire n_12910;
wire n_13349;
wire n_9956;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_10991;
wire n_14173;
wire n_10098;
wire n_11745;
wire n_8891;
wire n_4947;
wire n_3551;
wire n_11690;
wire n_9487;
wire n_3897;
wire n_11707;
wire n_5591;
wire n_11373;
wire n_7697;
wire n_14608;
wire n_6403;
wire n_7306;
wire n_13835;
wire n_7947;
wire n_10118;
wire n_14350;
wire n_7470;
wire n_7547;
wire n_6013;
wire n_7733;
wire n_13815;
wire n_13800;
wire n_7693;
wire n_9557;
wire n_6491;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_14039;
wire n_14072;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_13039;
wire n_13773;
wire n_13130;
wire n_14109;
wire n_8582;
wire n_10441;
wire n_5518;
wire n_6982;
wire n_10002;
wire n_5068;
wire n_6293;
wire n_6661;
wire n_9124;
wire n_5847;
wire n_13719;
wire n_7345;
wire n_6049;
wire n_9762;
wire n_8847;
wire n_11242;
wire n_8957;
wire n_14136;
wire n_7385;
wire n_10923;
wire n_14548;
wire n_5159;
wire n_4068;
wire n_6558;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_3703;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_13694;
wire n_12313;
wire n_3962;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_9543;
wire n_13688;
wire n_14661;
wire n_4166;
wire n_11396;
wire n_8356;
wire n_6136;
wire n_9660;
wire n_11443;
wire n_9483;
wire n_6855;
wire n_3745;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_4188;
wire n_13467;
wire n_5357;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_13093;
wire n_13062;
wire n_9328;
wire n_14252;
wire n_7857;
wire n_7481;
wire n_14130;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_6312;
wire n_8747;
wire n_9539;
wire n_6668;
wire n_4817;
wire n_11532;
wire n_9415;
wire n_4115;
wire n_14343;
wire n_9385;
wire n_3697;
wire n_9147;
wire n_11209;
wire n_7653;
wire n_13462;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_14276;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_13752;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_13185;
wire n_9027;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_4383;
wire n_13596;
wire n_6995;
wire n_10902;
wire n_4491;
wire n_12889;
wire n_13855;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_4486;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_11304;
wire n_9642;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_7475;
wire n_10485;
wire n_14231;
wire n_12105;
wire n_4612;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_13219;
wire n_14329;
wire n_5673;
wire n_5443;
wire n_6351;
wire n_9079;
wire n_9382;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_10444;
wire n_4529;
wire n_11377;
wire n_3478;
wire n_8018;
wire n_8653;
wire n_13295;
wire n_3936;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_5823;
wire n_7305;
wire n_13388;
wire n_3496;
wire n_13160;
wire n_13731;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_14550;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_14503;
wire n_4390;
wire n_12248;
wire n_13818;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_13477;
wire n_8884;
wire n_8803;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_10978;
wire n_5537;
wire n_8222;
wire n_13808;
wire n_14644;
wire n_6822;
wire n_3902;
wire n_4062;
wire n_11715;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_9706;
wire n_10642;
wire n_4233;
wire n_12181;
wire n_10187;
wire n_10387;
wire n_11014;
wire n_13764;
wire n_14560;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_11864;
wire n_3876;
wire n_11007;
wire n_11224;
wire n_11006;
wire n_9564;
wire n_7391;
wire n_8790;
wire n_9230;
wire n_6617;
wire n_4293;
wire n_10219;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_4684;
wire n_14067;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_14108;
wire n_6389;
wire n_5027;
wire n_6137;
wire n_10364;
wire n_10479;
wire n_11422;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_13660;
wire n_8398;
wire n_4412;
wire n_14480;
wire n_8178;
wire n_13970;
wire n_6801;
wire n_12489;
wire n_8491;
wire n_14000;
wire n_14372;
wire n_3618;
wire n_4580;
wire n_5630;
wire n_4758;
wire n_10065;
wire n_4781;
wire n_12046;
wire n_10212;
wire n_9283;
wire n_8700;
wire n_4148;
wire n_12030;
wire n_12738;
wire n_13408;
wire n_4057;
wire n_13727;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_10268;
wire n_14098;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_12601;
wire n_14482;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_13641;
wire n_14223;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_10559;
wire n_13173;
wire n_8439;
wire n_9641;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_12059;
wire n_12488;
wire n_3795;
wire n_7321;
wire n_5289;
wire n_3852;
wire n_4138;
wire n_8200;
wire n_11110;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_8304;
wire n_3815;
wire n_3896;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_13328;
wire n_7537;
wire n_10516;
wire n_4093;
wire n_8675;
wire n_10892;
wire n_6254;
wire n_5989;
wire n_10493;
wire n_13542;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_4794;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_14604;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_9016;
wire n_14426;
wire n_13101;
wire n_11887;
wire n_14349;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_11545;
wire n_9729;
wire n_5073;
wire n_12691;
wire n_8846;
wire n_8315;
wire n_12471;
wire n_11033;
wire n_12451;
wire n_4834;
wire n_11040;
wire n_12665;
wire n_11754;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_14356;
wire n_5581;
wire n_4762;
wire n_13748;
wire n_9029;
wire n_9411;
wire n_11672;
wire n_6837;
wire n_10353;
wire n_3813;
wire n_3660;
wire n_10847;
wire n_12651;
wire n_3766;
wire n_10451;
wire n_11043;
wire n_5303;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_9414;
wire n_7023;
wire n_3574;
wire n_9615;
wire n_12003;
wire n_14205;
wire n_7496;
wire n_11277;
wire n_14564;
wire n_4154;
wire n_12165;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_10866;
wire n_14190;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_3844;
wire n_8777;
wire n_4975;
wire n_11061;
wire n_11763;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_8535;
wire n_10653;
wire n_11534;
wire n_6373;
wire n_5375;
wire n_11587;
wire n_12280;
wire n_9221;
wire n_12492;
wire n_13461;
wire n_13581;
wire n_14344;
wire n_12972;
wire n_5370;
wire n_13789;
wire n_4898;
wire n_5601;
wire n_4815;
wire n_5784;
wire n_9811;
wire n_7899;
wire n_8631;
wire n_13188;
wire n_4819;
wire n_14511;
wire n_7906;
wire n_13286;
wire n_5248;
wire n_9951;
wire n_7131;
wire n_6411;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_14488;
wire n_11032;
wire n_5112;
wire n_13582;
wire n_4134;
wire n_10507;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_11843;
wire n_4092;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_14614;
wire n_13531;
wire n_7797;
wire n_3668;
wire n_11335;
wire n_11629;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_13880;
wire n_7687;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_13988;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_4087;
wire n_5635;
wire n_7582;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_13609;
wire n_3487;
wire n_14587;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_4302;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_6534;
wire n_10614;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_13679;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_5778;
wire n_8425;
wire n_11257;
wire n_8087;
wire n_13276;
wire n_9910;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_14458;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_11801;
wire n_13217;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_10743;
wire n_5165;
wire n_13424;
wire n_14658;
wire n_4884;
wire n_14397;
wire n_10853;
wire n_7867;
wire n_9651;
wire n_13565;
wire n_14281;
wire n_13755;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_6135;
wire n_13802;
wire n_14594;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_10270;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_11115;
wire n_8669;
wire n_12978;
wire n_13784;
wire n_8001;
wire n_7525;
wire n_13468;
wire n_7257;
wire n_12363;
wire n_9372;
wire n_7553;
wire n_7529;
wire n_4692;
wire n_6791;
wire n_14233;
wire n_8496;
wire n_11915;
wire n_13704;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_11788;
wire n_12544;
wire n_3890;
wire n_13036;
wire n_3750;
wire n_14146;
wire n_3607;
wire n_7650;
wire n_12476;
wire n_13199;
wire n_8568;
wire n_6903;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_4311;
wire n_12023;
wire n_8637;
wire n_6168;
wire n_6881;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_13413;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_13002;
wire n_12620;
wire n_12632;
wire n_7520;
wire n_9831;
wire n_13203;
wire n_13868;
wire n_4187;
wire n_6309;
wire n_7903;
wire n_9697;
wire n_11303;
wire n_11877;
wire n_6733;
wire n_14462;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_13285;
wire n_5430;
wire n_8610;
wire n_5942;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_9902;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_3532;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_9039;
wire n_12598;
wire n_11854;
wire n_13374;
wire n_12416;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_8704;
wire n_8265;
wire n_4619;
wire n_7639;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_5211;
wire n_5336;
wire n_11609;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_13230;
wire n_9294;
wire n_5036;
wire n_12811;
wire n_4221;
wire n_12186;
wire n_11747;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_12494;
wire n_13032;
wire n_13826;
wire n_7054;
wire n_7605;
wire n_11556;
wire n_11529;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_5327;
wire n_10021;
wire n_13684;
wire n_14199;
wire n_9146;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_14027;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_3803;
wire n_8941;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_9073;
wire n_10075;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_4334;
wire n_6171;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_12272;
wire n_9302;
wire n_5519;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_14684;
wire n_11895;
wire n_13458;
wire n_6269;
wire n_4047;
wire n_5753;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_8279;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_12191;
wire n_9580;
wire n_8019;
wire n_14572;
wire n_13963;
wire n_9972;
wire n_3791;
wire n_13003;
wire n_6083;
wire n_13091;
wire n_12909;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_4320;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_3884;
wire n_9465;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_13811;
wire n_14316;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_13839;
wire n_5231;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_14011;
wire n_4141;
wire n_13954;
wire n_10436;
wire n_8464;
wire n_6547;
wire n_8799;
wire n_12794;
wire n_5193;
wire n_6423;
wire n_9442;
wire n_6342;
wire n_6641;
wire n_6984;
wire n_12467;
wire n_5789;
wire n_10763;
wire n_7441;
wire n_9957;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_12112;
wire n_13060;
wire n_14689;
wire n_3883;
wire n_10245;
wire n_5961;
wire n_10905;
wire n_14132;
wire n_11235;
wire n_9449;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_6399;
wire n_4499;
wire n_6687;
wire n_9313;
wire n_5822;
wire n_9173;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_5726;
wire n_3949;
wire n_9563;
wire n_11015;
wire n_14087;
wire n_9160;
wire n_5364;
wire n_9974;
wire n_12129;
wire n_11166;
wire n_7031;
wire n_9285;
wire n_13658;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_9631;
wire n_14671;
wire n_8033;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_14438;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_13572;
wire n_12032;
wire n_4720;
wire n_10784;
wire n_12202;
wire n_4893;
wire n_14674;
wire n_3857;
wire n_13836;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_12815;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_9945;
wire n_8661;
wire n_12431;
wire n_7424;
wire n_3714;
wire n_7523;
wire n_8654;
wire n_5039;
wire n_11855;
wire n_4772;
wire n_14229;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_11156;
wire n_8531;
wire n_14188;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_4468;
wire n_13799;
wire n_5718;
wire n_4161;
wire n_6505;
wire n_6459;
wire n_12333;
wire n_12636;
wire n_8379;
wire n_8609;
wire n_13854;
wire n_4172;
wire n_11227;
wire n_7626;
wire n_13576;
wire n_13100;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_12334;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_9209;
wire n_3686;
wire n_7669;
wire n_11218;
wire n_4502;
wire n_12119;
wire n_11787;
wire n_12618;
wire n_5958;
wire n_8793;
wire n_12355;
wire n_8103;
wire n_9767;
wire n_10195;
wire n_9838;
wire n_13722;
wire n_4277;
wire n_4526;
wire n_9300;
wire n_11500;
wire n_3490;
wire n_4849;
wire n_12943;
wire n_7327;
wire n_4319;
wire n_14306;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_8367;
wire n_11891;
wire n_7367;
wire n_5792;
wire n_11021;
wire n_3581;
wire n_12401;
wire n_8543;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_6905;
wire n_3715;
wire n_10243;
wire n_9700;
wire n_10564;
wire n_8682;
wire n_3725;
wire n_13829;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_3933;
wire n_8533;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_7244;
wire n_10745;
wire n_7368;
wire n_3691;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_7633;
wire n_13937;
wire n_4146;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_10263;
wire n_5790;
wire n_4340;
wire n_11509;
wire n_8640;
wire n_14359;
wire n_8063;
wire n_3961;
wire n_11960;
wire n_4855;
wire n_12599;
wire n_3917;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_12411;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_12465;
wire n_7427;
wire n_10605;
wire n_4004;
wire n_11029;
wire n_13532;
wire n_14013;
wire n_13250;
wire n_13118;
wire n_14419;
wire n_5404;
wire n_9933;
wire n_11449;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_4292;
wire n_9892;
wire n_8570;
wire n_6163;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_14448;
wire n_10519;
wire n_5549;
wire n_9408;
wire n_6785;
wire n_6553;
wire n_10163;
wire n_10454;
wire n_3983;
wire n_13339;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_12568;
wire n_13478;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_12970;
wire n_8902;
wire n_8916;
wire n_14295;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_3510;
wire n_8843;
wire n_10146;
wire n_9891;
wire n_7128;
wire n_9946;
wire n_12959;
wire n_14367;
wire n_9885;
wire n_6849;
wire n_12330;
wire n_7594;
wire n_13915;
wire n_8129;
wire n_8162;
wire n_13906;
wire n_7457;
wire n_10643;
wire n_8744;
wire n_10504;
wire n_5824;
wire n_3719;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_13783;
wire n_6760;
wire n_10701;
wire n_3827;
wire n_5154;
wire n_13664;
wire n_13987;
wire n_14265;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_3889;
wire n_13566;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_13416;
wire n_12798;
wire n_5329;
wire n_9015;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_9925;
wire n_10874;
wire n_6825;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_11831;
wire n_13726;
wire n_9628;
wire n_14399;
wire n_7767;
wire n_14412;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_12243;
wire n_6611;
wire n_8562;
wire n_13705;
wire n_4560;
wire n_12614;
wire n_11378;
wire n_4899;
wire n_10250;
wire n_14631;
wire n_5728;
wire n_5471;
wire n_10032;
wire n_10592;
wire n_11433;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_14063;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_13425;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_7744;
wire n_7021;
wire n_10595;
wire n_13591;
wire n_7748;
wire n_8537;
wire n_10126;
wire n_6827;
wire n_14421;
wire n_12041;
wire n_4663;
wire n_11713;
wire n_11073;
wire n_13653;
wire n_5484;
wire n_6355;
wire n_12566;
wire n_12931;
wire n_6227;
wire n_13680;
wire n_7215;
wire n_7485;
wire n_13074;
wire n_9066;
wire n_4802;
wire n_5523;
wire n_14332;
wire n_10302;
wire n_11974;
wire n_12881;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_10645;
wire n_13058;
wire n_5074;
wire n_10604;
wire n_11096;
wire n_12036;
wire n_12876;
wire n_4044;
wire n_6564;
wire n_11161;
wire n_9671;
wire n_8782;
wire n_8709;
wire n_12911;
wire n_6468;
wire n_12491;
wire n_3937;
wire n_10080;
wire n_11216;
wire n_14368;
wire n_12228;
wire n_10570;
wire n_9857;
wire n_4701;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_14323;
wire n_12929;
wire n_10882;
wire n_9338;
wire n_13071;
wire n_6857;
wire n_8144;
wire n_12261;
wire n_3576;
wire n_10435;
wire n_9542;
wire n_12536;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_12061;
wire n_12106;
wire n_3922;
wire n_14585;
wire n_11085;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_10609;
wire n_11157;
wire n_13649;
wire n_13739;
wire n_4991;
wire n_5594;
wire n_12291;
wire n_14510;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_12124;
wire n_11755;
wire n_9783;
wire n_13806;
wire n_14364;
wire n_9510;
wire n_9389;
wire n_12074;
wire n_4934;
wire n_13497;
wire n_9404;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5087;
wire n_14396;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_13234;
wire n_5292;
wire n_9314;
wire n_11918;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_14466;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5000;
wire n_5403;
wire n_14473;
wire n_12887;
wire n_5551;
wire n_7652;
wire n_10220;
wire n_10341;
wire n_8701;
wire n_11347;
wire n_4479;
wire n_6499;
wire n_10550;
wire n_7830;
wire n_14673;
wire n_4011;
wire n_5131;
wire n_12217;
wire n_12365;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_13738;
wire n_13851;
wire n_9679;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_14138;
wire n_13272;
wire n_4688;
wire n_4753;
wire n_8712;
wire n_10232;
wire n_4058;
wire n_14113;
wire n_10461;
wire n_14586;
wire n_8289;
wire n_11178;
wire n_3611;
wire n_7966;
wire n_4848;
wire n_8591;
wire n_5059;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_8824;
wire n_11673;
wire n_11432;
wire n_14641;
wire n_14179;
wire n_14031;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_10412;
wire n_4475;
wire n_5242;
wire n_10326;
wire n_12650;
wire n_5219;
wire n_8417;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_3537;
wire n_10499;
wire n_8340;
wire n_6008;
wire n_3887;
wire n_4443;
wire n_12487;
wire n_12658;
wire n_14324;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_5460;
wire n_4587;
wire n_4114;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_13613;
wire n_9210;
wire n_12185;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_6893;
wire n_5686;
wire n_5899;
wire n_7406;
wire n_8681;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_10617;
wire n_12271;
wire n_12704;
wire n_7807;
wire n_4749;
wire n_9592;
wire n_5155;
wire n_14198;
wire n_7680;
wire n_9180;
wire n_10922;
wire n_10544;
wire n_12958;
wire n_13030;
wire n_3654;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_12056;
wire n_14539;
wire n_8106;
wire n_9502;
wire n_4100;
wire n_13821;
wire n_6447;
wire n_13712;
wire n_4264;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_3788;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_6422;
wire n_13896;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_3837;
wire n_14420;
wire n_11087;
wire n_11477;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_4085;
wire n_13299;
wire n_13243;
wire n_4464;
wire n_14314;
wire n_8612;
wire n_13042;
wire n_14144;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_10095;
wire n_14227;
wire n_4659;
wire n_13725;
wire n_10309;
wire n_3600;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_14164;
wire n_6160;
wire n_9871;
wire n_10050;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_7066;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_7789;
wire n_13197;
wire n_10306;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_7193;
wire n_3987;
wire n_6039;
wire n_4487;
wire n_11919;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_10450;
wire n_5721;
wire n_11472;
wire n_11414;
wire n_3638;
wire n_9114;
wire n_11978;
wire n_4816;
wire n_12520;
wire n_8515;
wire n_10529;
wire n_13632;
wire n_5719;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_8812;
wire n_14505;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_9392;
wire n_13148;
wire n_10429;
wire n_4937;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_14531;
wire n_3615;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_11538;
wire n_10037;
wire n_12808;
wire n_13871;
wire n_4222;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_13435;
wire n_4401;
wire n_12744;
wire n_6064;
wire n_11136;
wire n_9903;
wire n_4015;
wire n_13801;
wire n_5793;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_4709;
wire n_9228;
wire n_10179;
wire n_11539;
wire n_4976;
wire n_7710;
wire n_12143;
wire n_9499;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_13879;
wire n_6647;
wire n_6275;
wire n_4120;
wire n_14038;
wire n_9522;
wire n_5578;
wire n_11215;
wire n_4658;
wire n_5296;
wire n_11076;
wire n_9366;
wire n_11890;
wire n_14339;
wire n_14253;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_9148;
wire n_11806;
wire n_11054;
wire n_8406;
wire n_6277;
wire n_10754;
wire n_5742;
wire n_5207;
wire n_11050;
wire n_3705;
wire n_12443;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_11683;
wire n_8554;
wire n_10920;
wire n_9275;
wire n_10223;
wire n_6051;
wire n_8896;
wire n_14398;
wire n_4665;
wire n_3582;
wire n_11484;
wire n_7206;
wire n_4223;
wire n_11126;
wire n_7538;
wire n_5674;
wire n_12934;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_5282;
wire n_10295;
wire n_9409;
wire n_5464;
wire n_6799;
wire n_10336;
wire n_10228;
wire n_12555;
wire n_4362;
wire n_3913;
wire n_7716;
wire n_6487;
wire n_11646;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_8818;
wire n_4430;
wire n_8617;
wire n_4348;
wire n_12980;
wire n_13966;
wire n_9881;
wire n_12530;
wire n_5013;
wire n_8954;
wire n_6807;
wire n_9463;
wire n_7251;
wire n_4839;
wire n_7254;
wire n_4489;
wire n_12212;
wire n_10466;
wire n_12973;
wire n_7540;
wire n_11953;
wire n_4404;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_13231;
wire n_12624;
wire n_7882;
wire n_8552;
wire n_10425;
wire n_7554;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_8373;
wire n_10848;
wire n_13165;
wire n_6481;
wire n_5628;
wire n_4825;
wire n_7765;
wire n_11482;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_12151;
wire n_4006;
wire n_11089;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_13422;
wire n_6384;
wire n_3869;
wire n_7421;
wire n_13828;
wire n_10166;
wire n_7489;
wire n_7541;
wire n_6906;
wire n_4747;
wire n_13179;
wire n_14562;
wire n_5251;
wire n_3753;
wire n_12033;
wire n_11839;
wire n_3742;
wire n_9844;
wire n_3683;
wire n_8318;
wire n_4801;
wire n_12826;
wire n_14376;
wire n_13834;
wire n_10366;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_11365;
wire n_9595;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_11217;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_13923;
wire n_9287;
wire n_7991;
wire n_13051;
wire n_6233;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_14686;
wire n_12214;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_13330;
wire n_8926;
wire n_6257;
wire n_4386;
wire n_4132;
wire n_10361;
wire n_11228;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_13924;
wire n_4955;
wire n_8965;
wire n_11290;
wire n_5936;
wire n_4149;
wire n_12518;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_9052;
wire n_13476;
wire n_14047;
wire n_8817;
wire n_8190;
wire n_11488;
wire n_13671;
wire n_12162;
wire n_6587;
wire n_14627;
wire n_6987;
wire n_7781;
wire n_7360;
wire n_11037;
wire n_14568;
wire n_11702;
wire n_6069;
wire n_13699;
wire n_14319;
wire n_7497;
wire n_4655;
wire n_11372;
wire n_5706;
wire n_7665;
wire n_9354;
wire n_10817;
wire n_10501;
wire n_11829;
wire n_14026;
wire n_11517;
wire n_7793;
wire n_8355;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_12741;
wire n_7101;
wire n_7671;
wire n_9436;
wire n_7530;
wire n_8489;
wire n_13150;
wire n_13776;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_13343;
wire n_7654;
wire n_13152;
wire n_8303;
wire n_6153;
wire n_5132;
wire n_4374;
wire n_6637;
wire n_8369;
wire n_9022;
wire n_9238;
wire n_13809;
wire n_8059;
wire n_6633;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_6579;
wire n_11665;
wire n_13590;
wire n_13907;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_11138;
wire n_11731;
wire n_5187;
wire n_5875;
wire n_9839;
wire n_12821;
wire n_4024;
wire n_8831;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_6569;
wire n_7120;
wire n_6335;
wire n_8728;
wire n_10807;
wire n_12478;
wire n_12837;
wire n_12233;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_8853;
wire n_14070;
wire n_4582;
wire n_14330;
wire n_13491;
wire n_6252;
wire n_13545;
wire n_13471;
wire n_13760;
wire n_13883;
wire n_4860;
wire n_6211;
wire n_10511;
wire n_5844;
wire n_8862;
wire n_10580;
wire n_14235;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_9675;
wire n_7786;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_10058;
wire n_10873;
wire n_14484;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_11454;
wire n_13442;
wire n_8900;
wire n_12523;
wire n_14444;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_10484;
wire n_4304;
wire n_4558;
wire n_6737;
wire n_11744;
wire n_4488;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_14307;
wire n_8478;
wire n_6606;
wire n_13450;
wire n_6695;
wire n_3550;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_4211;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_14178;
wire n_11626;
wire n_12148;
wire n_4016;
wire n_11072;
wire n_5867;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_12907;
wire n_3839;
wire n_8497;
wire n_10770;
wire n_8820;
wire n_6410;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_5597;
wire n_9028;
wire n_13944;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_9374;
wire n_7419;
wire n_6506;
wire n_5515;
wire n_5662;
wire n_13634;
wire n_12132;
wire n_3730;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_10593;
wire n_13019;
wire n_14452;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_13464;
wire n_4397;
wire n_12182;
wire n_12670;
wire n_5050;
wire n_10636;
wire n_12043;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_10203;
wire n_3498;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_8992;
wire n_12708;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_6234;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_9983;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_13573;
wire n_6608;
wire n_10467;
wire n_3533;
wire n_9109;
wire n_9849;
wire n_13622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_11207;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_5498;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_9237;
wire n_13931;
wire n_11668;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_14404;
wire n_8466;
wire n_6753;
wire n_12137;
wire n_6527;
wire n_7341;
wire n_11328;
wire n_9349;
wire n_12306;
wire n_4908;
wire n_11200;
wire n_12088;
wire n_14442;
wire n_11091;
wire n_8094;
wire n_4109;
wire n_4192;
wire n_10940;
wire n_14377;
wire n_6639;
wire n_4824;
wire n_4567;
wire n_12096;
wire n_6430;
wire n_12508;
wire n_5150;
wire n_13418;
wire n_8832;
wire n_10987;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_4595;
wire n_4174;
wire n_12891;
wire n_11098;
wire n_11615;
wire n_10533;
wire n_11059;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_14616;
wire n_11965;
wire n_4904;
wire n_10938;
wire n_10176;
wire n_7517;
wire n_6627;
wire n_8080;
wire n_3544;
wire n_5988;
wire n_4150;
wire n_5585;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_7745;
wire n_12941;
wire n_13551;
wire n_14006;
wire n_6666;
wire n_3692;
wire n_10927;
wire n_14258;
wire n_12200;
wire n_4616;
wire n_8321;
wire n_14024;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_4982;
wire n_11722;
wire n_8592;
wire n_8786;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_4643;
wire n_13682;
wire n_6249;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_9805;
wire n_5480;
wire n_10155;
wire n_4323;
wire n_13593;
wire n_8157;
wire n_4831;
wire n_7095;
wire n_3821;
wire n_11461;
wire n_13902;
wire n_10714;
wire n_11701;
wire n_6969;
wire n_6615;
wire n_7459;
wire n_6161;
wire n_7294;
wire n_8206;
wire n_3676;
wire n_4896;
wire n_3666;
wire n_3675;
wire n_4260;
wire n_4017;
wire n_4916;
wire n_9110;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_8622;
wire n_5904;
wire n_13917;
wire n_4739;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_9335;
wire n_13546;
wire n_14595;
wire n_14468;
wire n_6062;
wire n_7908;
wire n_12550;
wire n_9452;
wire n_4122;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_13350;
wire n_13861;
wire n_10051;
wire n_4209;
wire n_8104;
wire n_10414;
wire n_11255;
wire n_8344;
wire n_13592;
wire n_3858;
wire n_5284;
wire n_11720;
wire n_4298;
wire n_12673;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_9075;
wire n_12961;
wire n_13874;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_4128;
wire n_10746;
wire n_12225;
wire n_9188;
wire n_6294;
wire n_5147;
wire n_9611;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_8779;
wire n_9810;
wire n_14469;
wire n_8621;
wire n_5503;
wire n_9250;
wire n_5845;
wire n_5945;
wire n_11212;
wire n_9550;
wire n_12884;
wire n_13145;
wire n_10697;
wire n_11714;
wire n_11263;
wire n_10641;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_12207;
wire n_9975;
wire n_7250;
wire n_5600;
wire n_5755;
wire n_8762;
wire n_12011;
wire n_13195;
wire n_8043;
wire n_8694;
wire n_14492;
wire n_13965;
wire n_5048;
wire n_6053;
wire n_11994;
wire n_7252;
wire n_13419;
wire n_9207;
wire n_13358;
wire n_14134;
wire n_4944;
wire n_11860;
wire n_11990;
wire n_10103;
wire n_5245;
wire n_6843;
wire n_4343;
wire n_10926;
wire n_14519;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_10626;
wire n_6901;
wire n_14345;
wire n_4935;
wire n_13273;
wire n_4694;
wire n_11503;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_8376;
wire n_8171;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_7698;
wire n_5749;
wire n_6774;
wire n_12854;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_8710;
wire n_12806;
wire n_4045;
wire n_3517;
wire n_3893;
wire n_4598;
wire n_3932;
wire n_14302;
wire n_3469;
wire n_8599;
wire n_8549;
wire n_13460;
wire n_10172;
wire n_5993;
wire n_8054;
wire n_11273;
wire n_13904;
wire n_10400;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_6020;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_14035;
wire n_14496;
wire n_14467;
wire n_13218;
wire n_9096;
wire n_9081;
wire n_13952;
wire n_11697;
wire n_13076;
wire n_4084;
wire n_9236;
wire n_6844;
wire n_11762;
wire n_11969;
wire n_12950;
wire n_7914;
wire n_8628;
wire n_7891;
wire n_6521;
wire n_13028;
wire n_14413;
wire n_8857;
wire n_8517;
wire n_4850;
wire n_14243;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_6162;
wire n_10433;
wire n_6779;
wire n_8010;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_9116;
wire n_14096;
wire n_10774;
wire n_3972;
wire n_12332;
wire n_4153;
wire n_11034;
wire n_10901;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_3506;
wire n_7216;
wire n_3855;
wire n_12762;
wire n_11499;
wire n_13574;
wire n_10825;
wire n_14583;
wire n_4317;
wire n_8275;
wire n_6198;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_4088;
wire n_5685;
wire n_10761;
wire n_3776;
wire n_4235;
wire n_3711;
wire n_5459;
wire n_14057;
wire n_9035;
wire n_11579;
wire n_10398;
wire n_8291;
wire n_4143;
wire n_4170;
wire n_11535;
wire n_3642;
wire n_12558;
wire n_4650;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_7477;
wire n_5173;
wire n_4719;
wire n_5016;
wire n_12975;
wire n_11402;
wire n_6458;
wire n_4967;
wire n_7642;
wire n_9678;
wire n_11401;
wire n_8247;
wire n_6577;
wire n_12506;
wire n_13850;
wire n_6740;
wire n_12718;
wire n_12956;
wire n_11510;
wire n_6315;
wire n_10581;
wire n_12638;
wire n_14116;
wire n_4912;
wire n_4799;
wire n_9284;
wire n_12736;
wire n_4423;
wire n_5283;
wire n_5086;
wire n_9111;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_3602;
wire n_12086;
wire n_5170;
wire n_6910;
wire n_7604;
wire n_6262;
wire n_7703;
wire n_3515;
wire n_9606;
wire n_6319;
wire n_13459;
wire n_10470;
wire n_14268;
wire n_11589;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_5028;
wire n_5839;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_14127;
wire n_6536;
wire n_12747;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_8827;
wire n_10625;
wire n_8280;
wire n_12561;
wire n_12390;
wire n_14460;
wire n_5514;
wire n_13216;
wire n_8388;
wire n_12849;
wire n_10235;
wire n_11312;
wire n_3866;
wire n_6978;
wire n_13786;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_4543;
wire n_10445;
wire n_7378;
wire n_10738;
wire n_12866;
wire n_4157;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_9190;
wire n_6947;
wire n_11612;
wire n_4229;
wire n_9482;
wire n_5293;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_12900;
wire n_13414;
wire n_3865;
wire n_4073;
wire n_8569;
wire n_3629;
wire n_5400;
wire n_14598;
wire n_3920;
wire n_4892;
wire n_6140;
wire n_8877;
wire n_9412;
wire n_7498;
wire n_10679;
wire n_11323;
wire n_10799;
wire n_3846;
wire n_6321;
wire n_12914;
wire n_11916;
wire n_3512;
wire n_6819;
wire n_7501;
wire n_5201;
wire n_9506;
wire n_10136;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_10585;
wire n_12764;
wire n_13696;
wire n_4783;
wire n_11356;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_13322;
wire n_14238;
wire n_9092;
wire n_10034;
wire n_9451;
wire n_4910;
wire n_11148;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_13934;
wire n_6899;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_6592;
wire n_11280;
wire n_12337;
wire n_13254;
wire n_13466;
wire n_8686;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_14042;
wire n_7613;
wire n_3541;
wire n_11493;
wire n_6101;
wire n_9220;
wire n_14440;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_10860;
wire n_12763;
wire n_4930;
wire n_8588;
wire n_11339;
wire n_5623;
wire n_12273;
wire n_13875;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_4112;
wire n_12712;
wire n_14076;
wire n_11220;
wire n_9012;
wire n_4557;
wire n_13012;
wire n_4917;
wire n_8698;
wire n_8924;
wire n_12584;
wire n_14435;
wire n_3739;
wire n_4432;
wire n_14638;
wire n_10376;
wire n_12752;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_4593;
wire n_7238;
wire n_9994;
wire n_4465;
wire n_14226;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_11596;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_14278;
wire n_11885;
wire n_5117;
wire n_5663;
wire n_7572;
wire n_8214;
wire n_10224;
wire n_11955;
wire n_12777;
wire n_5990;
wire n_7043;
wire n_10777;
wire n_3721;
wire n_11462;
wire n_11732;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_13306;
wire n_12819;
wire n_14159;
wire n_14515;
wire n_8722;
wire n_11654;
wire n_12268;
wire n_10214;
wire n_8241;
wire n_8589;
wire n_12077;
wire n_3969;
wire n_12982;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_6281;
wire n_4231;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_4256;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_6311;
wire n_10469;
wire n_9229;
wire n_11194;
wire n_11480;
wire n_7590;
wire n_9342;
wire n_12237;
wire n_13271;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_5426;
wire n_10175;
wire n_11481;
wire n_5803;
wire n_13372;
wire n_9868;
wire n_11375;
wire n_5285;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_4335;
wire n_9311;
wire n_12275;
wire n_6593;
wire n_13742;
wire n_8630;
wire n_12376;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_4521;
wire n_8405;
wire n_8145;
wire n_10447;
wire n_9260;
wire n_7176;
wire n_14534;
wire n_8928;
wire n_13630;
wire n_7682;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_11925;
wire n_13700;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_10406;
wire n_5715;
wire n_12509;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_11985;
wire n_13527;
wire n_8447;
wire n_7901;
wire n_5395;
wire n_10522;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_13793;
wire n_11782;
wire n_6446;
wire n_10278;
wire n_14290;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_3802;
wire n_6996;
wire n_7218;
wire n_8828;
wire n_9430;
wire n_11407;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_12710;
wire n_6749;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_7005;
wire n_10408;
wire n_8572;
wire n_10798;
wire n_10965;
wire n_7732;
wire n_13325;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_9776;
wire n_11911;
wire n_6777;
wire n_4265;
wire n_11987;
wire n_11442;
wire n_8227;
wire n_12936;
wire n_12721;
wire n_5634;
wire n_5672;
wire n_8475;
wire n_11730;
wire n_10482;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_4105;
wire n_14064;
wire n_14524;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_12039;
wire n_4926;
wire n_11388;
wire n_11651;
wire n_14151;
wire n_8314;
wire n_9386;
wire n_10154;
wire n_5617;
wire n_7922;
wire n_13089;
wire n_10377;
wire n_5266;
wire n_5580;
wire n_4828;
wire n_10033;
wire n_9926;
wire n_11121;
wire n_13167;
wire n_11270;
wire n_12329;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_8311;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_3769;
wire n_12253;
wire n_11147;
wire n_12928;
wire n_5310;
wire n_9661;
wire n_9843;
wire n_9877;
wire n_8764;
wire n_14284;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_13001;
wire n_5390;
wire n_13232;
wire n_9901;
wire n_13320;
wire n_5593;
wire n_12990;
wire n_14246;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_8567;
wire n_11817;
wire n_13278;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_5237;
wire n_13597;
wire n_5133;
wire n_13488;
wire n_11042;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_13447;
wire n_3989;
wire n_7089;
wire n_7144;
wire n_7286;
wire n_11479;
wire n_11737;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_14681;
wire n_12028;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_13016;
wire n_11272;
wire n_13668;
wire n_13095;
wire n_14230;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_6332;
wire n_4303;
wire n_5853;
wire n_12048;
wire n_8283;
wire n_5982;
wire n_10930;
wire n_11600;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_14546;
wire n_7129;
wire n_4909;
wire n_13938;
wire n_12057;
wire n_6696;
wire n_3925;
wire n_13251;
wire n_9882;
wire n_9527;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_3472;
wire n_8516;
wire n_8302;
wire n_10637;
wire n_8317;
wire n_5376;
wire n_12229;
wire n_14003;
wire n_5106;
wire n_6116;
wire n_9205;
wire n_9511;
wire n_8167;
wire n_7859;
wire n_14315;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_13670;
wire n_7972;
wire n_11254;
wire n_13319;
wire n_4768;
wire n_11617;
wire n_13858;
wire n_13512;
wire n_9071;
wire n_7916;
wire n_3717;
wire n_9368;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_10415;
wire n_13069;
wire n_11711;
wire n_5410;
wire n_12362;
wire n_8944;
wire n_6167;
wire n_13233;
wire n_11931;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_8109;
wire n_13297;
wire n_9459;
wire n_14185;
wire n_5156;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_6307;
wire n_10410;
wire n_6094;
wire n_9098;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_9133;
wire n_12664;
wire n_7434;
wire n_4826;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_9504;
wire n_8975;
wire n_6267;
wire n_9063;
wire n_7787;
wire n_3903;
wire n_12360;
wire n_5998;
wire n_9268;
wire n_5304;
wire n_3854;
wire n_6568;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_10456;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_14083;
wire n_13186;
wire n_5916;
wire n_11907;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_10627;
wire n_10025;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_6299;
wire n_6813;
wire n_8825;
wire n_12969;
wire n_11753;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_8266;
wire n_5691;
wire n_12457;
wire n_4951;
wire n_8981;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_13519;
wire n_14170;
wire n_4039;
wire n_3800;
wire n_13496;
wire n_4566;
wire n_12939;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_13884;
wire n_10404;
wire n_8639;
wire n_8058;
wire n_8138;
wire n_9308;
wire n_3504;
wire n_6638;
wire n_12779;
wire n_11838;
wire n_10508;
wire n_7719;
wire n_4272;
wire n_10811;
wire n_14049;
wire n_8333;
wire n_5615;
wire n_6220;
wire n_7562;
wire n_13547;
wire n_12816;
wire n_7619;
wire n_6985;
wire n_12783;
wire n_7170;
wire n_13853;
wire n_9211;
wire n_12019;
wire n_8176;
wire n_8124;
wire n_14529;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_10891;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_10803;
wire n_8147;
wire n_13190;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_14195;
wire n_5262;
wire n_10700;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_11695;
wire n_4620;
wire n_7935;
wire n_4738;
wire n_5421;
wire n_3579;
wire n_8458;
wire n_14247;
wire n_6772;
wire n_8113;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_14300;
wire n_11453;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_6318;
wire n_11970;
wire n_4099;
wire n_14678;
wire n_7918;
wire n_13599;
wire n_4517;
wire n_13354;
wire n_4168;
wire n_14690;
wire n_5188;
wire n_13647;
wire n_6916;
wire n_4490;
wire n_13683;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_10783;
wire n_11862;
wire n_10147;
wire n_12163;
wire n_10725;
wire n_3952;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_12944;
wire n_3911;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_11660;
wire n_4285;
wire n_10812;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_14249;
wire n_6230;
wire n_14241;
wire n_6604;
wire n_14497;
wire n_5161;
wire n_5373;
wire n_10001;
wire n_3708;
wire n_11107;
wire n_14280;
wire n_4078;
wire n_13724;
wire n_13280;
wire n_9301;
wire n_12145;
wire n_11088;
wire n_5573;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_8160;
wire n_10284;
wire n_12757;
wire n_12054;
wire n_14379;
wire n_5659;
wire n_8099;
wire n_14446;
wire n_11595;
wire n_8840;
wire n_3619;
wire n_11405;
wire n_13768;
wire n_13189;
wire n_5881;
wire n_8522;
wire n_12971;
wire n_7222;
wire n_7942;
wire n_8578;
wire n_6473;
wire n_13103;
wire n_13838;
wire n_4198;
wire n_3754;
wire n_10046;
wire n_12328;
wire n_14558;
wire n_11318;
wire n_9083;
wire n_7725;
wire n_10977;
wire n_4213;
wire n_11299;
wire n_10397;
wire n_6483;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_4065;
wire n_14004;
wire n_5863;
wire n_7647;
wire n_8626;
wire n_10936;
wire n_12442;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_9835;
wire n_7300;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_4446;
wire n_14666;
wire n_13605;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_13995;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_4733;
wire n_13441;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_14237;
wire n_3879;
wire n_11240;
wire n_4743;
wire n_10207;
wire n_13857;
wire n_13841;
wire n_13556;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_13367;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_13816;
wire n_11487;
wire n_11441;
wire n_8441;
wire n_14203;
wire n_6076;
wire n_8933;
wire n_7778;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_11287;
wire n_4060;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_4879;
wire n_6390;
wire n_10139;
wire n_13246;
wire n_13409;
wire n_14061;
wire n_5796;
wire n_10104;
wire n_8726;
wire n_12986;
wire n_11381;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_9117;
wire n_9720;
wire n_7746;
wire n_3662;
wire n_9381;
wire n_10169;
wire n_6958;
wire n_12049;
wire n_12690;
wire n_14498;
wire n_7563;
wire n_12475;
wire n_3624;
wire n_4556;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_14667;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_12526;
wire n_4687;
wire n_14414;
wire n_7531;
wire n_12377;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_13214;
wire n_8615;
wire n_11062;
wire n_13650;
wire n_7721;
wire n_7192;
wire n_14202;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_14554;
wire n_9887;
wire n_9149;
wire n_4600;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_13211;
wire n_8316;
wire n_4250;
wire n_9990;
wire n_5829;
wire n_3906;
wire n_10005;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_4954;
wire n_5191;
wire n_8505;
wire n_9273;
wire n_3963;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_13061;
wire n_9682;
wire n_4881;
wire n_12513;
wire n_4253;
wire n_10640;
wire n_6582;
wire n_5734;
wire n_13395;
wire n_4255;
wire n_4071;
wire n_10729;
wire n_12545;
wire n_14656;
wire n_7388;
wire n_3568;
wire n_3850;
wire n_11657;
wire n_9924;
wire n_8717;
wire n_13336;
wire n_5770;
wire n_5705;
wire n_4605;
wire n_9064;
wire n_7635;
wire n_5525;
wire n_13102;
wire n_11268;
wire n_12753;
wire n_7090;
wire n_4691;
wire n_9254;
wire n_12894;
wire n_14135;
wire n_3943;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_4305;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_13390;
wire n_13375;
wire n_13691;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_4297;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_14194;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_12010;
wire n_9738;
wire n_5675;
wire n_9570;
wire n_12026;
wire n_4227;
wire n_12356;
wire n_11857;
wire n_13825;
wire n_11077;
wire n_6240;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_9593;
wire n_7689;
wire n_9846;
wire n_13262;
wire n_13482;
wire n_6511;
wire n_5297;
wire n_7121;
wire n_9469;
wire n_10764;
wire n_13398;
wire n_9677;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_14676;
wire n_8449;
wire n_6358;
wire n_13204;
wire n_4094;
wire n_14331;
wire n_6603;
wire n_4765;
wire n_13873;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_8201;
wire n_8967;
wire n_6986;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_8801;
wire n_9322;
wire n_10438;
wire n_5959;
wire n_11201;
wire n_3720;
wire n_10531;
wire n_8031;
wire n_8918;
wire n_12878;
wire n_9348;
wire n_14262;
wire n_12188;
wire n_8219;
wire n_8696;
wire n_4745;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_12630;
wire n_4581;
wire n_6890;
wire n_11028;
wire n_12171;
wire n_4377;
wire n_12299;
wire n_12022;
wire n_9249;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_8180;
wire n_10741;
wire n_6109;
wire n_10760;
wire n_4792;
wire n_12425;
wire n_9444;
wire n_7731;
wire n_3842;
wire n_10772;
wire n_11527;
wire n_7114;
wire n_4878;
wire n_13507;
wire n_3514;
wire n_11327;
wire n_10915;
wire n_4979;
wire n_9535;
wire n_6770;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_5302;
wire n_12000;
wire n_4511;
wire n_9707;
wire n_12490;
wire n_13594;
wire n_5639;
wire n_5781;
wire n_14182;
wire n_3895;
wire n_8943;
wire n_8486;
wire n_10279;
wire n_4520;
wire n_5299;
wire n_12829;
wire n_4118;
wire n_4503;
wire n_14352;
wire n_13889;
wire n_10680;
wire n_10127;
wire n_3599;
wire n_5543;
wire n_13654;
wire n_5361;
wire n_11610;
wire n_7081;
wire n_7132;
wire n_11814;
wire n_12255;
wire n_12739;
wire n_13015;
wire n_4199;
wire n_5885;
wire n_6663;
wire n_14228;
wire n_9723;
wire n_5356;
wire n_12609;
wire n_7319;
wire n_4441;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_11176;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_11360;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5038;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_10039;
wire n_11726;
wire n_10854;
wire n_11358;
wire n_5463;
wire n_13366;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_12904;
wire n_8833;
wire n_9191;
wire n_5489;
wire n_5892;
wire n_7828;
wire n_10142;
wire n_4773;
wire n_14623;
wire n_7940;
wire n_9918;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_6009;
wire n_9034;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_9390;
wire n_5113;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_8074;
wire n_8485;
wire n_13639;
wire n_8860;
wire n_5510;
wire n_11958;
wire n_3940;
wire n_6621;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_13070;
wire n_8271;
wire n_5692;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_4800;
wire n_9266;
wire n_14491;
wire n_12728;
wire n_5555;
wire n_10027;
wire n_12784;
wire n_3768;
wire n_4958;
wire n_4043;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_13678;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_14582;
wire n_8699;
wire n_3785;
wire n_14261;
wire n_14677;
wire n_6897;
wire n_13523;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_5366;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_13778;
wire n_14250;
wire n_4886;
wire n_9931;
wire n_13198;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_13741;
wire n_13819;
wire n_4055;
wire n_12610;
wire n_14634;
wire n_11671;
wire n_10328;
wire n_14416;
wire n_5968;
wire n_11251;
wire n_14424;
wire n_14523;
wire n_12293;
wire n_11063;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_13174;
wire n_4200;
wire n_7108;
wire n_14455;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_8368;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_11879;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_8546;
wire n_10963;
wire n_8300;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_14161;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_8148;
wire n_11400;
wire n_13290;
wire n_8150;
wire n_13500;
wire n_3578;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_10483;
wire n_12160;
wire n_4737;
wire n_11563;
wire n_4925;
wire n_9620;
wire n_4116;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_5419;
wire n_11243;
wire n_3805;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_14513;
wire n_7260;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_6409;
wire n_11939;
wire n_7954;
wire n_9824;
wire n_11119;
wire n_14347;
wire n_7951;
wire n_7552;
wire n_8096;
wire n_11468;
wire n_14602;
wire n_13901;
wire n_12166;
wire n_8233;
wire n_6130;
wire n_4603;
wire n_7273;
wire n_9683;
wire n_10646;
wire n_7231;
wire n_5080;
wire n_5976;
wire n_11704;
wire n_14074;
wire n_5732;
wire n_5372;
wire n_14050;
wire n_11878;
wire n_4471;
wire n_7449;
wire n_7772;
wire n_8763;
wire n_12800;
wire n_5208;
wire n_14197;
wire n_8679;
wire n_7239;
wire n_14289;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_6623;
wire n_9561;
wire n_13951;
wire n_10378;
wire n_13968;
wire n_13979;
wire n_12070;
wire n_9714;
wire n_9740;
wire n_9773;
wire n_13316;
wire n_10313;
wire n_3838;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_13689;
wire n_3941;
wire n_3793;
wire n_10216;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_12354;
wire n_12666;
wire n_14297;
wire n_14395;
wire n_13528;
wire n_6047;
wire n_12581;
wire n_8292;
wire n_12631;
wire n_10133;
wire n_3729;
wire n_8601;
wire n_10773;
wire n_4994;
wire n_6652;
wire n_9377;
wire n_11932;
wire n_10971;
wire n_8830;
wire n_5347;
wire n_4483;
wire n_6921;
wire n_6970;
wire n_5168;
wire n_4661;
wire n_13027;
wire n_12867;
wire n_4988;
wire n_7674;
wire n_14675;
wire n_9826;
wire n_12607;
wire n_14516;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_12075;
wire n_4540;
wire n_11942;
wire n_6344;
wire n_12305;
wire n_13489;
wire n_12123;
wire n_9772;
wire n_12170;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_6624;
wire n_9630;
wire n_6956;
wire n_4284;
wire n_13313;
wire n_13927;
wire n_12966;
wire n_13877;
wire n_6305;
wire n_9255;
wire n_6209;
wire n_8310;
wire n_10231;
wire n_12547;
wire n_9758;
wire n_11922;
wire n_4971;
wire n_14020;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_5125;
wire n_5857;
wire n_12358;
wire n_7329;
wire n_14502;
wire n_8646;
wire n_7408;
wire n_13415;
wire n_9691;
wire n_12997;
wire n_14533;
wire n_10259;
wire n_14005;
wire n_7107;
wire n_14293;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_14334;
wire n_7690;
wire n_8969;
wire n_14187;
wire n_7123;
wire n_10752;
wire n_11577;
wire n_5499;
wire n_8117;
wire n_10067;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_13562;
wire n_14537;
wire n_12498;
wire n_13888;
wire n_11475;
wire n_6950;
wire n_8208;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_11010;
wire n_10274;
wire n_9590;
wire n_11588;
wire n_6694;
wire n_3497;
wire n_13956;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_9168;
wire n_3580;
wire n_14220;
wire n_11221;
wire n_13837;
wire n_12387;
wire n_9497;
wire n_8536;
wire n_13255;
wire n_9435;
wire n_7229;
wire n_14245;
wire n_8350;
wire n_3704;
wire n_11448;
wire n_9219;
wire n_5507;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_8914;
wire n_12576;
wire n_7258;
wire n_5190;
wire n_13892;
wire n_8391;
wire n_14221;
wire n_10579;
wire n_10832;
wire n_13345;
wire n_13964;
wire n_13749;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_6466;
wire n_14559;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_14360;
wire n_10584;
wire n_4218;
wire n_5392;
wire n_12862;
wire n_11445;
wire n_13151;
wire n_3880;
wire n_13601;
wire n_13621;
wire n_14052;
wire n_14311;
wire n_3685;
wire n_8216;
wire n_11552;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_11874;
wire n_13926;
wire n_3609;
wire n_9982;
wire n_10171;
wire n_14157;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_14317;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_12656;
wire n_9852;
wire n_6820;
wire n_11623;
wire n_8313;
wire n_3471;
wire n_5511;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_4175;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_10540;
wire n_11936;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_4771;
wire n_10200;
wire n_13392;
wire n_7332;
wire n_12734;
wire n_10382;
wire n_13164;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_13662;
wire n_3867;
wire n_10269;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_12262;
wire n_13223;
wire n_13340;
wire n_9169;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_5834;
wire n_10229;
wire n_5584;
wire n_13728;
wire n_7512;
wire n_14385;
wire n_4140;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_7766;
wire n_11018;
wire n_8738;
wire n_10981;
wire n_14499;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_12797;
wire n_6223;
wire n_11376;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_9481;
wire n_13379;
wire n_9600;
wire n_13781;
wire n_9122;
wire n_8085;
wire n_11274;
wire n_5098;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_5707;
wire n_12012;
wire n_5140;
wire n_4992;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_9927;
wire n_14613;
wire n_5497;
wire n_10076;
wire n_11515;
wire n_8721;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_3505;
wire n_13558;
wire n_3540;
wire n_3577;
wire n_11554;
wire n_7637;
wire n_10148;
wire n_10318;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_7127;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_4533;
wire n_9635;
wire n_13890;
wire n_5481;
wire n_12890;
wire n_3590;
wire n_8666;
wire n_5344;
wire n_9264;
wire n_13994;
wire n_14483;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_14308;
wire n_5408;
wire n_7801;
wire n_13484;
wire n_9155;
wire n_4053;
wire n_10234;
wire n_8460;
wire n_3848;
wire n_10416;
wire n_14370;
wire n_14593;
wire n_8836;
wire n_7959;
wire n_13430;
wire n_7019;
wire n_8181;
wire n_11325;
wire n_8254;
wire n_13452;
wire n_13521;
wire n_4167;
wire n_8071;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_10731;
wire n_10583;
wire n_10735;
wire n_9878;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_13807;
wire n_14591;
wire n_14363;
wire n_9825;
wire n_5494;
wire n_7444;
wire n_11628;
wire n_14576;
wire n_5234;
wire n_7546;
wire n_4431;
wire n_6272;
wire n_4387;
wire n_14274;
wire n_6588;
wire n_11549;
wire n_5128;
wire n_3755;
wire n_4042;
wire n_14033;
wire n_12286;
wire n_9001;
wire n_10393;
wire n_11498;
wire n_13081;
wire n_10513;
wire n_12252;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_14545;
wire n_12627;
wire n_4890;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_12281;
wire n_14272;
wire n_11237;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_9373;
wire n_14337;
wire n_6268;
wire n_5827;
wire n_4176;
wire n_12347;
wire n_5199;
wire n_14551;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_11181;
wire n_13651;
wire n_9967;
wire n_13553;
wire n_7521;
wire n_14088;
wire n_5992;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_13817;
wire n_3856;
wire n_4236;
wire n_7187;
wire n_9971;
wire n_10894;
wire n_3894;
wire n_14118;
wire n_13974;
wire n_9524;
wire n_12277;
wire n_12698;
wire n_5312;
wire n_3623;
wire n_6467;
wire n_9243;
wire n_9182;
wire n_9282;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_9224;
wire n_3646;
wire n_10347;
wire n_5513;
wire n_5614;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_12410;
wire n_4830;
wire n_4706;
wire n_13225;
wire n_5225;
wire n_4570;
wire n_10208;
wire n_7722;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_8141;
wire n_14612;
wire n_12294;
wire n_14180;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_14058;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_13355;
wire n_12957;
wire n_4693;
wire n_13141;
wire n_4206;
wire n_11616;
wire n_14065;
wire n_8791;
wire n_11920;
wire n_10793;
wire n_8288;
wire n_14672;
wire n_3862;
wire n_14366;
wire n_4267;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_12786;
wire n_5049;
wire n_13382;
wire n_12711;
wire n_11675;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_5846;
wire n_8323;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_10440;
wire n_10391;
wire n_7636;
wire n_9695;
wire n_9799;
wire n_11083;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_7866;
wire n_4609;
wire n_11306;
wire n_13176;
wire n_9784;
wire n_11198;
wire n_7205;
wire n_8757;
wire n_7990;
wire n_7020;
wire n_13035;
wire n_10036;
wire n_13021;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_8596;
wire n_3525;
wire n_5157;
wire n_11840;
wire n_4754;
wire n_11698;
wire n_4647;
wire n_9556;
wire n_3688;
wire n_11292;
wire n_8590;
wire n_8720;
wire n_10261;
wire n_13157;
wire n_5708;
wire n_4003;
wire n_3751;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_4894;
wire n_5474;
wire n_14084;
wire n_12289;
wire n_4113;
wire n_10813;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_11326;
wire n_13046;
wire n_6421;
wire n_13935;
wire n_11870;
wire n_7407;
wire n_9827;
wire n_14009;
wire n_3466;
wire n_13334;
wire n_10907;
wire n_5704;
wire n_11431;
wire n_4983;
wire n_7148;
wire n_14002;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_13646;
wire n_6236;
wire n_9417;
wire n_11834;
wire n_13361;
wire n_12020;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_3907;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_6835;
wire n_8834;
wire n_3636;
wire n_11624;
wire n_13399;
wire n_14010;
wire n_8826;
wire n_11352;
wire n_5516;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_10822;
wire n_11234;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_13967;
wire n_12099;
wire n_12858;
wire n_3539;
wire n_7467;
wire n_4399;
wire n_14609;
wire n_7799;
wire n_8364;
wire n_5698;
wire n_11092;
wire n_9534;
wire n_14310;
wire n_13380;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_3572;
wire n_11836;
wire n_6602;
wire n_10924;
wire n_3886;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_9647;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_10885;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_13201;
wire n_3637;
wire n_6242;
wire n_12527;
wire n_4574;
wire n_13274;
wire n_12379;
wire n_9312;
wire n_9019;
wire n_13891;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_4234;
wire n_12477;
wire n_7469;
wire n_5538;
wire n_14325;
wire n_14078;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_14309;
wire n_10895;
wire n_3974;
wire n_10875;
wire n_3634;
wire n_11736;
wire n_11977;
wire n_7560;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_14222;
wire n_11696;
wire n_12400;
wire n_5096;
wire n_11734;
wire n_12114;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_11507;
wire n_14430;
wire n_9145;
wire n_13996;
wire n_7082;
wire n_12092;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_4270;
wire n_11837;
wire n_5428;
wire n_4151;
wire n_13709;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_13898;
wire n_9000;
wire n_5677;
wire n_9454;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_8307;
wire n_5153;
wire n_11967;
wire n_9383;
wire n_9253;
wire n_13559;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_5927;
wire n_7392;
wire n_7495;
wire n_9566;
wire n_11338;
wire n_11996;
wire n_5435;
wire n_13426;
wire n_12174;
wire n_9765;
wire n_9807;
wire n_4333;
wire n_9057;
wire n_5200;
wire n_3820;
wire n_8706;
wire n_6400;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_6941;
wire n_5115;
wire n_12053;
wire n_5566;
wire n_11250;
wire n_7829;
wire n_12619;
wire n_7543;
wire n_13504;
wire n_8680;
wire n_11289;
wire n_13169;
wire n_7877;
wire n_7963;
wire n_13555;
wire n_9672;
wire n_12582;
wire n_4152;
wire n_5487;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_5486;
wire n_9503;
wire n_12423;
wire n_11391;
wire n_5244;
wire n_5092;
wire n_14137;
wire n_13265;
wire n_8270;
wire n_4832;
wire n_12714;
wire n_12153;
wire n_5889;
wire n_11738;
wire n_7284;
wire n_7264;
wire n_5391;
wire n_11522;
wire n_9763;
wire n_14163;
wire n_7737;
wire n_13666;
wire n_6537;
wire n_8614;
wire n_11070;
wire n_7328;
wire n_10702;
wire n_13337;
wire n_10958;
wire n_9479;
wire n_9162;
wire n_9568;
wire n_13730;
wire n_3536;
wire n_12405;
wire n_8816;
wire n_3957;
wire n_14041;
wire n_3710;
wire n_9119;
wire n_4195;
wire n_10319;
wire n_5849;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_13529;
wire n_6224;
wire n_6578;
wire n_8802;
wire n_9859;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_6092;
wire n_10879;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_10639;
wire n_3475;
wire n_3501;
wire n_8121;
wire n_3905;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_12554;
wire n_13351;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_10491;
wire n_12037;
wire n_13453;
wire n_5152;
wire n_5265;
wire n_12792;
wire n_11717;
wire n_9943;
wire n_4927;
wire n_5574;
wire n_12391;
wire n_14242;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_7152;
wire n_11723;
wire n_9575;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_11830;
wire n_12438;
wire n_5469;
wire n_14393;
wire n_8766;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_12838;
wire n_6567;
wire n_9165;
wire n_13505;
wire n_14016;
wire n_12323;
wire n_5910;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_14369;
wire n_7240;
wire n_7570;
wire n_4553;
wire n_7033;
wire n_10476;
wire n_4875;
wire n_9966;
wire n_13156;
wire n_7817;
wire n_5682;
wire n_10710;
wire n_5387;
wire n_5557;
wire n_11394;
wire n_8850;
wire n_11906;
wire n_9928;
wire n_11820;
wire n_14647;
wire n_14298;
wire n_8002;
wire n_9741;
wire n_13897;
wire n_11486;
wire n_12677;
wire n_4321;
wire n_10180;
wire n_4183;
wire n_14248;
wire n_14112;
wire n_8370;
wire n_7237;
wire n_13300;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_9090;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_4901;
wire n_4145;
wire n_4821;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_12901;
wire n_4040;
wire n_10518;
wire n_8301;
wire n_12895;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_9771;
wire n_13401;
wire n_5316;
wire n_7718;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_13844;
wire n_14122;
wire n_7396;
wire n_10942;
wire n_12668;
wire n_12726;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_13010;
wire n_6320;
wire n_8126;
wire n_11239;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4943;
wire n_10953;
wire n_12432;
wire n_4757;
wire n_7561;
wire n_6810;
wire n_7842;
wire n_12352;
wire n_9969;
wire n_6202;
wire n_10099;
wire n_11437;
wire n_4682;
wire n_9961;
wire n_12898;
wire n_14068;
wire n_12879;
wire n_5564;
wire n_11869;
wire n_13746;
wire n_12559;
wire n_13508;
wire n_5620;
wire n_14660;
wire n_7163;
wire n_4530;
wire n_10343;
wire n_10836;
wire n_4942;
wire n_9899;
wire n_9258;
wire n_13004;
wire n_10181;
wire n_10286;
wire n_5406;
wire n_8072;
wire n_10371;
wire n_13479;
wire n_8277;
wire n_7236;
wire n_4604;
wire n_13117;
wire n_10257;
wire n_5724;
wire n_7130;
wire n_7201;
wire n_11219;
wire n_4841;
wire n_14437;
wire n_10047;
wire n_14541;
wire n_13759;
wire n_5806;
wire n_10949;
wire n_4338;
wire n_13766;
wire n_10486;
wire n_11282;
wire n_11226;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_11413;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_5355;
wire n_5320;
wire n_3984;
wire n_7491;
wire n_13969;
wire n_5353;
wire n_9995;
wire n_13710;
wire n_5186;
wire n_5710;
wire n_9076;
wire n_11232;
wire n_12351;
wire n_12693;
wire n_9105;
wire n_6792;
wire n_12080;
wire n_5093;
wire n_4052;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_13359;
wire n_9668;
wire n_3558;
wire n_10372;
wire n_7559;
wire n_5438;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_13259;
wire n_4326;
wire n_13335;
wire n_14022;
wire n_12702;
wire n_13175;
wire n_5517;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_10744;
wire n_12648;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_5907;
wire n_11334;
wire n_6045;
wire n_13075;
wire n_13129;
wire n_13736;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_14186;
wire n_7526;
wire n_5040;
wire n_14023;
wire n_6063;
wire n_10736;
wire n_10917;
wire n_6504;
wire n_3761;
wire n_11575;
wire n_4315;
wire n_7004;
wire n_7821;
wire n_14418;
wire n_12407;
wire n_13586;
wire n_8308;
wire n_6154;
wire n_11284;
wire n_6943;
wire n_4301;
wire n_10597;
wire n_14668;
wire n_11827;
wire n_13049;
wire n_3744;
wire n_8165;
wire n_13961;
wire n_14283;
wire n_12038;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_8210;
wire n_11656;
wire n_12644;
wire n_5977;
wire n_10446;
wire n_13134;
wire n_11826;
wire n_7879;
wire n_10271;
wire n_3814;
wire n_3781;
wire n_10888;
wire n_10116;
wire n_7696;
wire n_11570;
wire n_6003;
wire n_12952;
wire n_6684;
wire n_3843;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_5451;
wire n_9323;
wire n_14140;
wire n_3687;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_9331;
wire n_3621;
wire n_6031;
wire n_9922;
wire n_10170;
wire n_13252;
wire n_11909;
wire n_8331;
wire n_12024;
wire n_13084;
wire n_14479;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_12004;
wire n_12830;
wire n_12637;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_4365;
wire n_6060;
wire n_7929;
wire n_10255;
wire n_10572;
wire n_14172;
wire n_3726;
wire n_12009;
wire n_13612;
wire n_7270;
wire n_13985;
wire n_11490;
wire n_3758;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_14124;
wire n_10113;
wire n_7550;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_6853;
wire n_6742;
wire n_10188;
wire n_13525;
wire n_4923;
wire n_5864;
wire n_10686;
wire n_9841;
wire n_13552;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_12681;
wire n_14207;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_12634;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_13863;
wire n_8627;
wire n_14305;
wire n_9513;
wire n_9863;
wire n_12680;
wire n_11613;
wire n_4885;
wire n_13659;
wire n_10233;
wire n_12034;
wire n_10500;
wire n_10555;
wire n_5432;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_11929;
wire n_10810;
wire n_11075;
wire n_7851;
wire n_6894;
wire n_13303;
wire n_13346;
wire n_12176;
wire n_9791;
wire n_13702;
wire n_10311;
wire n_9179;
wire n_5453;
wire n_13656;
wire n_3658;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_11177;
wire n_13667;
wire n_4408;
wire n_4577;
wire n_6817;
wire n_4748;
wire n_5842;
wire n_10937;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_12449;
wire n_5814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_11310;
wire n_13275;
wire n_12094;
wire n_6215;
wire n_11165;
wire n_4212;
wire n_9736;
wire n_5699;
wire n_5531;
wire n_14411;
wire n_5765;
wire n_12823;
wire n_12517;
wire n_6517;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_10167;
wire n_7862;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_6883;
wire n_4225;
wire n_8808;
wire n_10061;
wire n_12963;
wire n_10428;
wire n_13087;
wire n_13972;
wire n_11865;
wire n_12366;
wire n_8528;
wire n_8204;
wire n_13024;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_5495;
wire n_10694;
wire n_12339;
wire n_10602;
wire n_7100;
wire n_12729;
wire n_3583;
wire n_13292;
wire n_12198;
wire n_3860;
wire n_11041;
wire n_14632;
wire n_9420;
wire n_3851;
wire n_14490;
wire n_5655;
wire n_6393;
wire n_9708;
wire n_14336;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_8154;
wire n_6966;
wire n_8889;
wire n_13986;
wire n_9790;
wire n_13849;
wire n_13796;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_4009;
wire n_5002;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_13258;
wire n_6035;
wire n_3473;
wire n_7874;
wire n_8490;
wire n_7622;
wire n_13329;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_13166;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_13946;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_6364;
wire n_14464;
wire n_8635;
wire n_7102;
wire n_7420;
wire n_4342;
wire n_12605;
wire n_13618;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_7831;
wire n_6253;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_8532;
wire n_14327;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_14097;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_11140;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_8796;
wire n_12218;
wire n_4106;
wire n_5737;
wire n_3604;
wire n_12343;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_12597;
wire n_12316;
wire n_14454;
wire n_4711;
wire n_13744;
wire n_11478;
wire n_12834;
wire n_10066;
wire n_13017;
wire n_12236;
wire n_14335;
wire n_12902;
wire n_6419;
wire n_8372;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_3553;
wire n_10088;
wire n_13038;
wire n_7225;
wire n_8077;
wire n_12892;
wire n_3811;
wire n_11294;
wire n_3494;
wire n_6244;
wire n_9812;
wire n_6900;
wire n_9337;
wire n_3486;
wire n_4086;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_9432;
wire n_9949;
wire n_10289;
wire n_6942;
wire n_7705;
wire n_11819;
wire n_7228;
wire n_13762;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_7932;
wire n_4812;
wire n_11573;
wire n_4409;
wire n_9576;
wire n_7509;
wire n_10145;
wire n_13420;
wire n_5872;
wire n_6862;
wire n_14225;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_6840;
wire n_13005;
wire n_6338;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_6037;
wire n_7981;
wire n_9577;
wire n_9874;
wire n_3699;
wire n_12588;
wire n_4913;
wire n_12589;
wire n_5874;
wire n_6266;
wire n_14143;
wire n_6488;
wire n_8337;
wire n_7164;
wire n_9231;
wire n_11844;
wire n_14044;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_11364;
wire n_3868;
wire n_9569;
wire n_13184;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_13535;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_8358;
wire n_10009;
wire n_9552;
wire n_12927;
wire n_11100;
wire n_9279;
wire n_13822;
wire n_11902;
wire n_6317;
wire n_8199;
wire n_5588;
wire n_11993;
wire n_4012;
wire n_10443;
wire n_8656;
wire n_7167;
wire n_10756;
wire n_12813;
wire n_6480;
wire n_3645;
wire n_14387;
wire n_10918;
wire n_13122;
wire n_13534;
wire n_5075;
wire n_11797;
wire n_3682;
wire n_4968;
wire n_3771;
wire n_12765;
wire n_14106;
wire n_7865;
wire n_13616;
wire n_12663;
wire n_10384;
wire n_9289;
wire n_5085;
wire n_11315;
wire n_5736;
wire n_4259;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_7134;
wire n_9633;
wire n_11153;
wire n_12312;
wire n_10074;
wire n_4572;
wire n_4845;
wire n_9547;
wire n_4104;
wire n_13097;
wire n_6875;
wire n_13627;
wire n_10934;
wire n_10197;
wire n_8346;
wire n_5120;
wire n_4208;
wire n_8761;
wire n_13112;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_13734;
wire n_8226;
wire n_11949;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_9084;
wire n_5928;
wire n_12256;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_11746;
wire n_11812;
wire n_9371;
wire n_14051;
wire n_13163;
wire n_3702;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_4779;
wire n_14650;
wire n_7267;
wire n_10367;
wire n_14610;
wire n_4599;
wire n_12315;
wire n_11505;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_14100;
wire n_12375;
wire n_12556;
wire n_12998;
wire n_7812;
wire n_7103;
wire n_13723;
wire n_13143;
wire n_9080;
wire n_4061;
wire n_14601;
wire n_14549;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_9519;
wire n_6367;
wire n_3881;
wire n_11363;
wire n_12156;
wire n_13564;
wire n_14459;
wire n_13128;
wire n_4508;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_11530;
wire n_12671;
wire n_10621;
wire n_13411;
wire n_7056;
wire n_14645;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_13260;
wire n_4642;
wire n_4051;
wire n_7813;
wire n_10085;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_6080;
wire n_4865;
wire n_8182;
wire n_8387;
wire n_12525;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_12076;
wire n_14090;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_13758;
wire n_7200;
wire n_11359;
wire n_7688;
wire n_4562;
wire n_8707;
wire n_12357;
wire n_4903;
wire n_3709;
wire n_10561;
wire n_11434;
wire n_3738;
wire n_9208;
wire n_11791;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_13212;
wire n_14463;
wire n_8494;
wire n_5812;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_11848;
wire n_13503;
wire n_3610;
wire n_11152;
wire n_4998;
wire n_10749;
wire n_11632;
wire n_7795;
wire n_14166;
wire n_12180;
wire n_8788;
wire n_14405;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_14081;
wire n_7723;
wire n_4341;
wire n_11621;
wire n_10160;
wire n_9327;
wire n_10560;
wire n_7404;
wire n_12857;
wire n_13171;
wire n_5368;
wire n_4263;
wire n_8177;
wire n_3555;
wire n_9854;
wire n_14271;
wire n_7059;
wire n_7450;
wire n_11667;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_12208;
wire n_6145;
wire n_11964;
wire n_6539;
wire n_6926;
wire n_13421;
wire n_7271;
wire n_7826;
wire n_9713;
wire n_14565;
wire n_11298;
wire n_5933;
wire n_13495;
wire n_8993;
wire n_6204;
wire n_7076;
wire n_13474;
wire n_4780;
wire n_10300;
wire n_13949;
wire n_13314;
wire n_9588;
wire n_11403;
wire n_14218;
wire n_11741;
wire n_12383;
wire n_11912;
wire n_3908;
wire n_4973;
wire n_6842;
wire n_3467;
wire n_12773;
wire n_6866;
wire n_13876;
wire n_9044;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_3950;
wire n_9423;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_14487;
wire n_4750;
wire n_12962;
wire n_6451;
wire n_9813;
wire n_9127;
wire n_14596;
wire n_6514;
wire n_3740;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_9244;
wire n_9869;
wire n_11142;
wire n_7049;
wire n_5903;
wire n_14449;
wire n_5986;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_12885;
wire n_11644;
wire n_6345;
wire n_9715;
wire n_8618;
wire n_12108;
wire n_9094;
wire n_13108;
wire n_5782;
wire n_7535;
wire n_5041;
wire n_13170;
wire n_4275;
wire n_10862;
wire n_11531;
wire n_4283;
wire n_4959;
wire n_8248;
wire n_9056;
wire n_8911;
wire n_11357;
wire n_14471;
wire n_4426;
wire n_9407;
wire n_11476;
wire n_14476;
wire n_4425;
wire n_13633;
wire n_9985;
wire n_4449;
wire n_12089;
wire n_12496;
wire n_14538;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_11959;
wire n_11367;
wire n_6957;
wire n_9361;
wire n_11921;
wire n_4809;
wire n_8495;
wire n_14532;
wire n_12676;
wire n_13976;
wire n_8783;
wire n_12987;
wire n_13579;
wire n_14557;
wire n_11566;
wire n_13913;
wire n_8529;
wire n_8733;
wire n_14639;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_10254;
wire n_14340;
wire n_14032;
wire n_7944;
wire n_13080;
wire n_11208;
wire n_7262;
wire n_3773;
wire n_8647;
wire n_11374;
wire n_12967;
wire n_12452;
wire n_13403;
wire n_8574;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_13557;
wire n_12232;
wire n_4241;
wire n_11859;
wire n_12818;
wire n_10386;
wire n_12128;
wire n_6379;
wire n_14060;
wire n_14018;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_5563;
wire n_13583;
wire n_11026;
wire n_14111;
wire n_8044;
wire n_13309;
wire n_5840;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9439;
wire n_9553;
wire n_11633;
wire n_11467;
wire n_7506;
wire n_12672;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_14361;
wire n_8330;
wire n_12760;
wire n_4050;
wire n_13455;
wire n_6232;
wire n_9132;
wire n_13172;
wire n_5717;
wire n_6017;
wire n_9696;
wire n_10861;
wire n_9120;
wire n_8879;
wire n_11203;
wire n_11159;
wire n_8052;
wire n_12168;
wire n_4578;
wire n_6362;
wire n_4777;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_14148;
wire n_8903;
wire n_11030;
wire n_4702;
wire n_12590;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_12924;
wire n_7142;
wire n_12577;
wire n_10182;
wire n_12732;
wire n_13928;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_9464;
wire n_9252;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_10073;
wire n_4531;
wire n_11655;
wire n_14619;
wire n_5072;
wire n_3626;
wire n_11017;
wire n_12843;
wire n_7241;
wire n_7247;
wire n_14279;
wire n_12069;
wire n_10419;
wire n_7172;
wire n_14622;
wire n_10333;
wire n_12430;
wire n_10317;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_4029;
wire n_7235;
wire n_8540;
wire n_11248;
wire n_12613;
wire n_6239;
wire n_12270;
wire n_14365;
wire n_9915;
wire n_4617;
wire n_9325;
wire n_9196;
wire n_13407;
wire n_4010;
wire n_5896;
wire n_5882;
wire n_4555;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_13676;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_13788;
wire n_14555;
wire n_11141;
wire n_5105;
wire n_12695;
wire n_10893;
wire n_4308;
wire n_11093;
wire n_5021;
wire n_14219;
wire n_9251;
wire n_11576;
wire n_8939;
wire n_13584;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_8468;
wire n_4325;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_13181;
wire n_5134;
wire n_7096;
wire n_12210;
wire n_13327;
wire n_8778;
wire n_11197;
wire n_3998;
wire n_7442;
wire n_3632;
wire n_10093;
wire n_5567;
wire n_8343;
wire n_6174;
wire n_12006;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_14168;
wire n_6087;
wire n_7593;
wire n_12246;
wire n_5249;
wire n_14085;
wire n_8068;
wire n_9955;
wire n_3829;
wire n_10539;
wire n_14080;
wire n_4164;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_4919;
wire n_3737;
wire n_10107;
wire n_13975;
wire n_5969;
wire n_3655;
wire n_10196;
wire n_10121;
wire n_8198;
wire n_14573;
wire n_3825;
wire n_13085;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_13224;
wire n_11469;
wire n_6454;
wire n_5022;
wire n_12625;
wire n_9270;
wire n_14046;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_14142;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_14512;
wire n_8557;
wire n_6041;
wire n_6918;
wire n_9099;
wire n_12389;
wire n_13761;
wire n_9309;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_10814;
wire n_5276;
wire n_9627;
wire n_13971;
wire n_11252;
wire n_8012;
wire n_14456;
wire n_13364;
wire n_7672;
wire n_11494;
wire n_6664;
wire n_5047;
wire n_7318;
wire n_6472;
wire n_10218;
wire n_8114;
wire n_13131;
wire n_3792;
wire n_4202;
wire n_12995;
wire n_14406;
wire n_3938;
wire n_13209;
wire n_4791;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_5879;
wire n_14563;
wire n_8062;
wire n_4403;
wire n_11883;
wire n_5238;
wire n_11256;
wire n_11832;
wire n_6166;
wire n_5855;
wire n_12370;
wire n_3531;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_10975;
wire n_11901;
wire n_6352;
wire n_12974;
wire n_9460;
wire n_8542;
wire n_12136;
wire n_10859;
wire n_13078;
wire n_7063;
wire n_7047;
wire n_11652;
wire n_4139;
wire n_14320;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_13885;
wire n_6238;
wire n_10542;
wire n_8038;
wire n_13631;
wire n_13932;
wire n_3931;
wire n_4349;
wire n_10681;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_11572;
wire n_13370;
wire n_5141;
wire n_11894;
wire n_3603;
wire n_14493;
wire n_10222;
wire n_6724;
wire n_13113;
wire n_13387;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_8716;
wire n_11336;
wire n_6705;
wire n_3822;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_4163;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_7074;
wire n_3910;
wire n_3812;
wire n_8734;
wire n_9204;
wire n_9689;
wire n_9476;
wire n_11849;
wire n_12142;
wire n_10659;
wire n_6591;
wire n_7585;
wire n_4948;
wire n_12564;
wire n_5268;
wire n_13643;
wire n_9780;
wire n_6946;
wire n_3482;
wire n_6002;
wire n_4080;
wire n_13433;
wire n_10403;
wire n_13607;
wire n_12983;
wire n_6289;
wire n_7037;
wire n_3748;
wire n_13697;
wire n_11784;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_14244;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_12886;
wire n_14114;
wire n_13980;
wire n_6532;
wire n_4372;
wire n_7293;
wire n_13000;
wire n_12035;
wire n_14362;
wire n_13006;
wire n_5640;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3978;
wire n_6721;
wire n_5560;
wire n_13205;
wire n_6644;
wire n_6512;
wire n_5544;
wire n_4074;
wire n_4795;
wire n_3716;
wire n_12810;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_4918;
wire n_3824;
wire n_9597;
wire n_5067;
wire n_13820;
wire n_13947;
wire n_11322;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_11892;
wire n_12122;
wire n_5384;
wire n_4544;
wire n_13428;
wire n_5841;
wire n_12241;
wire n_12396;
wire n_7614;
wire n_9343;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_4032;
wire n_6086;
wire n_9837;
wire n_11421;
wire n_11057;
wire n_4147;
wire n_10969;
wire n_10896;
wire n_4477;
wire n_11966;
wire n_14474;
wire n_12748;
wire n_7383;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_10562;
wire n_5941;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_14417;
wire n_3601;
wire n_5611;
wire n_6340;
wire n_10054;
wire n_10355;
wire n_6219;
wire n_7479;
wire n_6706;
wire n_11551;
wire n_3966;
wire n_12571;
wire n_11853;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_10598;
wire n_13034;
wire n_8947;
wire n_4742;
wire n_3734;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_7078;
wire n_8188;
wire n_13831;
wire n_6761;
wire n_8972;
wire n_10007;
wire n_3649;
wire n_11751;
wire n_11423;
wire n_11725;
wire n_5701;
wire n_3746;
wire n_13635;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_12674;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_9567;
wire n_14637;
wire n_6811;
wire n_9061;
wire n_11495;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_4478;
wire n_7372;
wire n_5367;
wire n_3794;
wire n_12220;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_10704;
wire n_11520;
wire n_11622;
wire n_4838;
wire n_5970;
wire n_12169;
wire n_12283;
wire n_12336;
wire n_7174;
wire n_13268;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_13383;
wire n_10457;
wire n_12543;
wire n_4965;
wire n_8021;
wire n_9705;
wire n_7803;
wire n_11012;
wire n_6111;
wire n_14158;
wire n_12595;
wire n_9624;
wire n_3861;
wire n_9701;
wire n_11502;
wire n_14236;
wire n_11429;
wire n_10389;
wire n_11631;
wire n_13588;
wire n_13510;
wire n_13570;
wire n_14640;
wire n_3891;
wire n_6659;
wire n_4523;
wire n_9709;
wire n_13677;
wire n_13983;
wire n_6011;
wire n_9295;
wire n_9416;
wire n_13757;
wire n_14036;
wire n_4371;
wire n_6225;
wire n_11842;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_5502;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_9929;
wire n_12920;
wire n_10264;
wire n_5850;
wire n_13317;
wire n_4673;
wire n_13910;
wire n_9953;
wire n_13737;
wire n_7086;
wire n_6648;
wire n_4607;
wire n_14286;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_12717;
wire n_4041;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_12141;
wire n_8584;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_13196;
wire n_13520;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_10301;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_13018;
wire n_7025;
wire n_9364;
wire n_8228;
wire n_8076;
wire n_6826;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_9836;
wire n_10929;
wire n_14357;
wire n_9107;
wire n_3809;
wire n_11279;
wire n_11724;
wire n_13044;
wire n_11789;
wire n_14152;
wire n_13228;
wire n_11525;
wire n_13518;
wire n_13862;
wire n_8100;
wire n_4070;
wire n_11999;
wire n_13446;
wire n_13086;
wire n_10837;
wire n_3545;
wire n_3885;
wire n_14008;
wire n_10554;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_12746;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_10149;
wire n_10970;
wire n_7768;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_14651;
wire n_5491;
wire n_5496;
wire n_3780;
wire n_5802;
wire n_13887;
wire n_7982;
wire n_12190;
wire n_12787;
wire n_8804;
wire n_13881;
wire n_11383;
wire n_12799;
wire n_4002;
wire n_11847;
wire n_11976;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_5547;
wire n_13747;
wire n_8158;
wire n_12511;
wire n_11167;
wire n_6879;
wire n_12532;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_3477;
wire n_8433;
wire n_10102;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_8213;
wire n_5983;
wire n_14472;
wire n_3953;
wire n_4588;
wire n_10534;
wire n_11825;
wire n_4653;
wire n_4435;
wire n_11049;
wire n_10619;
wire n_7684;
wire n_10932;
wire n_14354;
wire n_5604;
wire n_8451;
wire n_5411;
wire n_8334;
wire n_12743;
wire n_4019;
wire n_8731;
wire n_10589;
wire n_11681;
wire n_11611;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_11202;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_7370;
wire n_5815;
wire n_3616;
wire n_9748;
wire n_13365;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_13539;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_8539;
wire n_10205;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_14618;
wire n_9226;
wire n_3727;
wire n_5235;
wire n_10110;
wire n_13899;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_11688;
wire n_6888;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_12715;
wire n_11709;
wire n_12434;
wire n_14328;
wire n_12628;
wire n_8122;
wire n_6095;
wire n_13444;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_14209;
wire n_11331;
wire n_14429;
wire n_5311;
wire n_12979;
wire n_9528;
wire n_6590;
wire n_14348;
wire n_10638;
wire n_7583;
wire n_12201;
wire n_14086;
wire n_3522;
wire n_6559;
wire n_12499;
wire n_3924;
wire n_9112;
wire n_12448;
wire n_4621;
wire n_4216;
wire n_11876;
wire n_5797;
wire n_9235;
wire n_10610;
wire n_11187;
wire n_4240;
wire n_12761;
wire n_5572;
wire n_3491;
wire n_13852;
wire n_9333;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_14270;
wire n_8950;
wire n_14089;
wire n_10758;
wire n_13431;
wire n_10190;
wire n_5520;
wire n_11804;
wire n_14234;
wire n_3975;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_6287;
wire n_12809;
wire n_13614;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_14552;
wire n_7353;
wire n_9330;
wire n_12538;
wire n_14208;
wire n_14025;
wire n_7758;
wire n_4021;
wire n_13779;
wire n_12446;
wire n_9490;
wire n_12029;
wire n_4103;
wire n_9355;
wire n_11052;
wire n_5060;
wire n_9523;
wire n_14584;
wire n_4986;
wire n_4022;
wire n_14620;
wire n_5888;
wire n_5669;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_9582;
wire n_4775;
wire n_5884;
wire n_10060;
wire n_6671;
wire n_13470;
wire n_11009;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_9686;
wire n_9288;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_13068;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_11446;
wire n_10910;
wire n_10162;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_13248;
wire n_7792;
wire n_13842;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_14501;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_8703;
wire n_10014;
wire n_7109;
wire n_12642;
wire n_3731;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_8822;
wire n_6029;
wire n_10677;
wire n_12187;
wire n_5751;
wire n_5264;
wire n_4525;
wire n_12321;
wire n_5924;
wire n_9992;
wire n_11247;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_12669;
wire n_13106;
wire n_8476;
wire n_14296;
wire n_14294;
wire n_6702;
wire n_11927;
wire n_3620;
wire n_13720;
wire n_11179;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_13706;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_13903;
wire n_3693;
wire n_9051;
wire n_8545;
wire n_8736;
wire n_4497;
wire n_7749;
wire n_10078;
wire n_10105;
wire n_10385;
wire n_11514;
wire n_12470;
wire n_12994;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_8705;
wire n_14574;
wire n_10215;
wire n_14451;
wire n_11779;
wire n_14059;
wire n_7508;
wire n_3674;
wire n_5694;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_14211;
wire n_10834;
wire n_7574;
wire n_14092;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_14509;
wire n_4306;
wire n_14394;
wire n_11882;
wire n_13516;
wire n_11647;
wire n_4224;
wire n_12064;
wire n_14273;
wire n_10706;
wire n_12462;
wire n_6005;
wire n_8872;
wire n_12696;
wire n_4453;
wire n_9555;
wire n_11133;
wire n_5449;
wire n_3559;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_3546;
wire n_3661;
wire n_12735;
wire n_7713;
wire n_4564;
wire n_13560;
wire n_11222;
wire n_9200;
wire n_5146;
wire n_10709;
wire n_12646;
wire n_10871;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_10304;
wire n_5398;
wire n_4573;
wire n_5860;
wire n_6936;
wire n_4535;
wire n_14624;
wire n_10244;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_14120;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_7641;
wire n_13794;
wire n_6106;
wire n_3627;
wire n_3480;
wire n_7203;
wire n_12999;
wire n_13537;
wire n_14260;
wire n_14407;
wire n_9397;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_12682;
wire n_3612;
wire n_9673;
wire n_14434;
wire n_14175;
wire n_4695;
wire n_6848;
wire n_8642;
wire n_3509;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11941;
wire n_11875;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_12111;
wire n_8912;
wire n_14346;
wire n_7439;
wire n_13463;
wire n_9496;
wire n_8110;
wire n_14275;
wire n_5319;
wire n_10796;
wire n_14506;
wire n_10016;
wire n_12903;
wire n_9008;
wire n_12079;
wire n_6343;
wire n_12593;
wire n_14615;
wire n_5270;
wire n_10030;
wire n_8805;
wire n_6850;
wire n_12864;
wire n_5005;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_13294;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_13895;
wire n_11307;
wire n_5181;
wire n_13936;
wire n_13933;
wire n_6979;
wire n_7815;
wire n_13222;
wire n_7934;
wire n_9545;
wire n_13813;
wire n_8111;
wire n_9603;
wire n_9629;
wire n_11578;
wire n_6865;
wire n_10432;
wire n_12719;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_5043;
wire n_8739;
wire n_6747;
wire n_9674;
wire n_13714;
wire n_5583;
wire n_4654;
wire n_13438;
wire n_6433;
wire n_10462;
wire n_12725;
wire n_3640;
wire n_3481;
wire n_6640;
wire n_11769;
wire n_8856;
wire n_6142;
wire n_9930;
wire n_11908;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_6034;
wire n_10291;
wire n_9781;
wire n_13159;
wire n_4597;
wire n_9659;
wire n_4020;
wire n_14333;
wire n_7233;
wire n_8732;
wire n_13636;
wire n_13506;
wire n_13287;
wire n_11913;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_14590;
wire n_11341;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_13256;
wire n_10669;
wire n_13389;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_14603;
wire n_8231;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_13905;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_4063;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_4237;
wire n_13717;
wire n_5029;
wire n_5127;
wire n_12317;
wire n_13302;
wire n_6071;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_8908;
wire n_10185;
wire n_11182;
wire n_10092;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_12782;
wire n_4721;
wire n_11231;
wire n_14145;
wire n_8090;
wire n_13740;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_12875;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_13918;
wire n_8137;
wire n_7045;
wire n_13775;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_11727;
wire n_13615;
wire n_6788;
wire n_7014;
wire n_12192;
wire n_12633;
wire n_10430;
wire n_8305;
wire n_4614;
wire n_10277;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_6709;
wire n_14465;
wire n_13412;
wire n_4422;
wire n_10948;
wire n_11749;
wire n_6550;
wire n_6712;
wire n_10525;
wire n_9507;
wire n_14287;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_8841;
wire n_14553;
wire n_3870;
wire n_13457;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_6743;
wire n_12497;
wire n_4632;
wire n_10354;
wire n_12412;
wire n_11880;
wire n_5785;
wire n_7465;
wire n_14528;
wire n_13177;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_12724;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_9457;
wire n_4966;
wire n_9485;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_13940;
wire n_7936;
wire n_8966;
wire n_6084;
wire n_11249;
wire n_4847;
wire n_10287;
wire n_4054;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_14342;
wire n_12101;
wire n_10119;
wire n_13693;
wire n_11145;
wire n_3586;
wire n_12606;
wire n_11986;
wire n_3653;
wire n_8395;
wire n_10900;
wire n_5966;
wire n_10349;
wire n_6634;
wire n_14107;
wire n_4668;
wire n_5213;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_13333;
wire n_4635;
wire n_13229;
wire n_5735;
wire n_12118;
wire n_13311;
wire n_14409;
wire n_7490;
wire n_11380;
wire n_14291;
wire n_7545;
wire n_10792;
wire n_11513;
wire n_8625;
wire n_13296;
wire n_7160;
wire n_7464;
wire n_8937;
wire n_4214;
wire n_9809;
wire n_6919;
wire n_14611;
wire n_10750;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_7115;
wire n_7295;
wire n_12087;
wire n_13675;
wire n_9192;
wire n_3595;
wire n_14338;
wire n_7348;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_10537;
wire n_11861;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_10426;
wire n_4405;
wire n_4413;
wire n_9558;
wire n_11594;
wire n_7453;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_4036;
wire n_10684;
wire n_4759;
wire n_7162;
wire n_3670;
wire n_11436;
wire n_12346;
wire n_4667;
wire n_5081;
wire n_11729;
wire n_4182;
wire n_8371;
wire n_8702;
wire n_13916;
wire n_8116;
wire n_7946;
wire n_8195;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_14069;
wire n_12244;
wire n_5877;
wire n_9991;
wire n_14255;
wire n_11670;
wire n_11366;
wire n_11872;
wire n_7681;
wire n_8845;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_13620;
wire n_5189;
wire n_13930;
wire n_7702;
wire n_6676;
wire n_13981;
wire n_8149;
wire n_10823;
wire n_4637;
wire n_9976;
wire n_8042;
wire n_11516;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_8392;
wire n_9560;
wire n_14592;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_14659;
wire n_10830;
wire n_11132;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_6854;
wire n_4155;
wire n_4238;
wire n_4977;
wire n_13624;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_14277;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_13493;
wire n_6032;
wire n_9047;
wire n_13805;
wire n_12953;
wire n_12842;
wire n_3650;
wire n_8968;
wire n_12481;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_5446;
wire n_11316;
wire n_7855;
wire n_14029;
wire n_11047;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_4590;
wire n_8399;
wire n_5090;
wire n_14648;
wire n_11767;
wire n_9599;
wire n_14056;
wire n_3560;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_13866;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_13695;
wire n_12435;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_11586;
wire n_6981;
wire n_13288;
wire n_7065;
wire n_12149;
wire n_13669;
wire n_9216;
wire n_3529;
wire n_12002;
wire n_12836;
wire n_4835;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_13840;
wire n_11229;
wire n_13548;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_14251;
wire n_6122;
wire n_4038;
wire n_11397;
wire n_11225;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_4565;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_4159;
wire n_12840;
wire n_3784;
wire n_7330;
wire n_14605;
wire n_5437;
wire n_8883;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_13543;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_10577;
wire n_13772;
wire n_14679;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_7357;
wire n_8756;
wire n_11324;
wire n_8737;
wire n_13925;
wire n_10334;
wire n_4434;
wire n_12945;
wire n_13406;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_10151;
wire n_6439;
wire n_11614;
wire n_4290;
wire n_14040;
wire n_8602;
wire n_14054;
wire n_13368;
wire n_8240;
wire n_12850;
wire n_13469;
wire n_14507;
wire n_7714;
wire n_5407;
wire n_10411;
wire n_13249;
wire n_9484;
wire n_12984;
wire n_10989;
wire n_8422;
wire n_10939;
wire n_13587;
wire n_12224;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_8878;
wire n_11144;
wire n_10090;
wire n_6406;
wire n_7440;
wire n_11361;
wire n_6945;
wire n_8112;
wire n_14034;
wire n_11567;
wire n_3790;
wire n_10962;
wire n_7029;
wire n_11128;
wire n_9622;
wire n_9292;
wire n_10721;
wire n_8593;
wire n_12197;
wire n_14177;
wire n_14093;
wire n_10186;
wire n_14607;
wire n_4833;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_6618;
wire n_13326;
wire n_6474;
wire n_13082;
wire n_14453;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_13094;
wire n_7317;
wire n_10856;
wire n_12403;
wire n_6000;
wire n_12679;
wire n_13481;
wire n_9584;
wire n_3977;
wire n_8194;
wire n_9461;
wire n_8055;
wire n_11168;
wire n_13692;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_8360;
wire n_3588;
wire n_5008;
wire n_4279;
wire n_12018;
wire n_6425;
wire n_14457;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_9845;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_14382;
wire n_14389;
wire n_11937;
wire n_12872;
wire n_13396;
wire n_7522;
wire n_6492;
wire n_10071;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_6046;
wire n_11460;
wire n_14517;
wire n_8251;
wire n_13713;
wire n_5323;
wire n_11565;
wire n_4790;
wire n_4181;
wire n_14621;
wire n_12372;
wire n_9618;
wire n_6118;
wire n_13608;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_7046;
wire n_11192;
wire n_11808;
wire n_4007;
wire n_13257;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_4239;
wire n_8677;
wire n_13052;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_5991;
wire n_4184;
wire n_13914;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_14663;
wire n_5702;
wire n_10035;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_13922;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_3489;
wire n_13423;
wire n_8108;
wire n_14578;
wire n_5243;
wire n_5914;
wire n_12955;
wire n_12068;
wire n_10252;
wire n_5250;
wire n_11555;
wire n_13494;
wire n_6869;
wire n_10041;
wire n_9321;
wire n_14625;
wire n_5590;
wire n_10345;
wire n_14514;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_5809;
wire n_14256;
wire n_10543;
wire n_7924;
wire n_4782;
wire n_12394;
wire n_13578;
wire n_7659;
wire n_9005;
wire n_3530;
wire n_9161;
wire n_14204;
wire n_8875;
wire n_5349;
wire n_4378;
wire n_8274;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_12954;
wire n_7836;
wire n_10737;
wire n_12662;
wire n_4876;
wire n_14082;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_7280;
wire n_10644;
wire n_12801;
wire n_13448;
wire n_14688;
wire n_5813;
wire n_9293;
wire n_12503;
wire n_13708;
wire n_10365;
wire n_13767;
wire n_5833;
wire n_11781;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_12965;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_14571;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_5816;
wire n_10809;
wire n_8927;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_6228;
wire n_6711;
wire n_11997;
wire n_3483;
wire n_11884;
wire n_5416;
wire n_8946;
wire n_13090;
wire n_14527;
wire n_12822;
wire n_13541;
wire n_13307;
wire n_13371;
wire n_11863;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_12264;
wire n_13312;
wire n_11761;
wire n_8474;
wire n_9984;
wire n_3524;
wire n_7275;
wire n_8232;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_9649;
wire n_8904;
wire n_11199;
wire n_13533;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_10629;
wire n_9562;
wire n_7007;
wire n_7070;
wire n_4539;
wire n_8382;
wire n_4421;
wire n_13023;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_4793;
wire n_13856;
wire n_4498;
wire n_10006;
wire n_7259;
wire n_11757;
wire n_12274;
wire n_12320;
wire n_14588;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_12622;
wire n_6992;
wire n_11185;
wire n_8128;
wire n_12659;
wire n_13440;
wire n_6818;
wire n_3831;
wire n_13436;
wire n_10206;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5932;
wire n_5830;
wire n_3589;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12629;
wire n_7539;
wire n_12586;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_10275;
wire n_11081;
wire n_7775;
wire n_13011;
wire n_4505;
wire n_11392;
wire n_9981;
wire n_7930;
wire n_5558;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_13911;
wire n_5383;
wire n_14495;
wire n_5126;
wire n_8205;
wire n_14165;
wire n_5051;
wire n_9907;
wire n_13088;
wire n_5587;
wire n_6976;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_12269;
wire n_13538;
wire n_7640;
wire n_14617;
wire n_13701;
wire n_9816;
wire n_13787;
wire n_10498;
wire n_11424;
wire n_13486;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_13674;
wire n_14263;
wire n_11463;
wire n_13912;
wire n_14303;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_8605;
wire n_11278;
wire n_14445;
wire n_10358;
wire n_3787;
wire n_7548;
wire n_3585;
wire n_10635;
wire n_13626;
wire n_3565;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_12832;
wire n_12913;
wire n_5025;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_12301;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_14427;
wire n_7197;
wire n_5645;
wire n_9676;
wire n_3990;
wire n_11881;
wire n_7393;
wire n_11332;
wire n_6917;
wire n_13629;
wire n_6937;
wire n_7591;
wire n_13207;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_7727;
wire n_7358;
wire n_7324;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_11935;
wire n_13589;
wire n_4534;
wire n_6301;
wire n_9788;
wire n_6929;
wire n_11309;
wire n_8719;
wire n_8045;
wire n_10785;
wire n_7729;
wire n_13872;
wire n_12341;
wire n_12615;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_14475;
wire n_8209;
wire n_13357;
wire n_10802;
wire n_14477;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_6699;
wire n_12926;
wire n_9213;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_14522;
wire n_8784;
wire n_7382;
wire n_4811;
wire n_13869;
wire n_13955;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_13561;
wire n_12167;
wire n_9473;
wire n_14400;
wire n_4857;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_6677;
wire n_12161;
wire n_13499;
wire n_12085;
wire n_11735;
wire n_7618;
wire n_4282;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_6764;
wire n_8575;
wire n_13554;
wire n_12298;
wire n_10081;
wire n_5733;
wire n_3774;
wire n_10324;
wire n_11189;
wire n_6780;
wire n_8815;
wire n_11582;
wire n_12569;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_9303;
wire n_11105;
wire n_11705;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_7673;
wire n_13698;
wire n_6830;
wire n_13894;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_7282;
wire n_6586;
wire n_9968;
wire n_10808;
wire n_11474;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_13595;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_13943;
wire n_7953;
wire n_13540;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_14642;
wire n_9722;
wire n_13283;
wire n_12042;
wire n_12155;
wire n_5657;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_13465;
wire n_8695;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_4911;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_4436;
wire n_14579;
wire n_8363;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_8665;
wire n_13098;
wire n_13733;
wire n_6510;
wire n_8282;
wire n_9388;
wire n_5938;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_12654;
wire n_14141;
wire n_5602;
wire n_9379;
wire n_11992;
wire n_5097;
wire n_4985;
wire n_7751;
wire n_10869;
wire n_3823;
wire n_4384;
wire n_13142;
wire n_7581;
wire n_13180;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_14589;
wire n_5246;
wire n_3584;
wire n_10453;
wire n_12386;
wire n_14257;
wire n_4858;
wire n_4678;
wire n_13308;
wire n_9952;
wire n_3556;
wire n_9911;
wire n_12183;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_13785;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_12964;
wire n_10473;
wire n_14007;
wire n_5107;
wire n_5095;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_10957;
wire n_13373;
wire n_4243;
wire n_7579;
wire n_13517;
wire n_12863;
wire n_10352;
wire n_4025;
wire n_11188;
wire n_7428;
wire n_5666;
wire n_12221;
wire n_4059;
wire n_9195;
wire n_10442;
wire n_11687;
wire n_4121;
wire n_8870;
wire n_13973;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_11774;
wire n_7283;
wire n_3671;
wire n_6475;
wire n_7015;
wire n_4142;
wire n_4313;
wire n_3982;
wire n_7699;
wire n_8507;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_13206;
wire n_9623;
wire n_6103;
wire n_7249;
wire n_5546;
wire n_10713;
wire n_3796;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_14102;
wire n_6680;
wire n_7985;
wire n_10954;
wire n_13637;
wire n_4246;
wire n_12267;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_13941;
wire n_13978;
wire n_4532;
wire n_13439;
wire n_13780;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_14133;
wire n_14433;
wire n_11329;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_9516;
wire n_4244;
wire n_13241;
wire n_13187;
wire n_13162;
wire n_4049;
wire n_6752;
wire n_12768;
wire n_8976;
wire n_6426;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_8156;
wire n_11661;
wire n_7494;
wire n_4353;
wire n_11120;
wire n_9222;
wire n_13031;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_7736;
wire n_4787;
wire n_10622;
wire n_5633;
wire n_13661;
wire n_13155;
wire n_9546;
wire n_5664;
wire n_7589;
wire n_14259;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_13410;
wire n_4537;
wire n_14012;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_13066;
wire n_8660;
wire n_13360;
wire n_11296;
wire n_13665;
wire n_8479;
wire n_14214;
wire n_13770;
wire n_12993;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_3521;
wire n_11314;
wire n_8723;
wire n_13511;
wire n_11019;
wire n_8606;
wire n_9663;
wire n_7843;
wire n_6235;
wire n_8235;
wire n_13083;
wire n_3764;
wire n_12647;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_9820;
wire n_14569;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_14071;
wire n_9743;
wire n_6496;
wire n_7756;
wire n_12749;
wire n_8342;
wire n_8940;
wire n_13048;
wire n_11584;
wire n_5280;
wire n_8448;
wire n_13563;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_14169;
wire n_4332;
wire n_7555;
wire n_10000;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_10582;
wire n_12066;
wire n_12812;
wire n_3695;
wire n_10427;
wire n_11816;
wire n_12060;
wire n_3976;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_14174;
wire n_3563;
wire n_6513;
wire n_7500;
wire n_10246;
wire n_11910;
wire n_11693;
wire n_3495;
wire n_13347;
wire n_14269;
wire n_5925;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_9822;
wire n_10835;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_13991;
wire n_13823;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_13323;
wire n_12164;
wire n_5272;
wire n_11368;
wire n_10125;
wire n_12824;
wire n_13111;
wire n_13434;
wire n_6330;
wire n_10117;
wire n_9065;
wire n_12716;
wire n_10844;
wire n_14153;
wire n_8457;
wire n_6802;
wire n_13456;
wire n_10654;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_9339;
wire n_10198;
wire n_6909;
wire n_7157;
wire n_11064;
wire n_13237;
wire n_6908;
wire n_14312;
wire n_8237;
wire n_13445;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_11409;
wire n_4201;
wire n_4336;
wire n_7266;
wire n_8046;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_13284;
wire n_12437;
wire n_5624;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_10840;
wire n_12052;
wire n_6477;
wire n_9746;
wire n_14606;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_5440;
wire n_6490;
wire n_11605;
wire n_11533;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_7198;
wire n_8335;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_9440;
wire n_10144;
wire n_3955;
wire n_9684;
wire n_6184;
wire n_3945;
wire n_5817;
wire n_5214;
wire n_10973;
wire n_4936;
wire n_4205;
wire n_13472;
wire n_9493;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_11330;
wire n_12720;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_6038;
wire n_10551;
wire n_13318;
wire n_5861;
wire n_3833;
wire n_10553;
wire n_13127;
wire n_8309;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_12687;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_14075;
wire n_9032;
wire n_9814;
wire n_6313;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_13208;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_13867;
wire n_5859;
wire n_12325;
wire n_14423;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_13443;
wire n_5776;
wire n_8166;
wire n_5606;
wire n_4433;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_14626;
wire n_5826;
wire n_10108;
wire n_8960;
wire n_13865;
wire n_12789;
wire n_5920;
wire n_10307;
wire n_5030;
wire n_14530;
wire n_4194;
wire n_7994;
wire n_14206;
wire n_4703;
wire n_8443;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_6180;
wire n_8683;
wire n_14481;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_12127;
wire n_12382;
wire n_12504;
wire n_5756;
wire n_12602;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_13673;
wire n_12062;
wire n_14119;
wire n_4030;
wire n_12573;

CKINVDCx5p33_ASAP7_75t_R g3466 ( 
.A(n_2751),
.Y(n_3466)
);

CKINVDCx5p33_ASAP7_75t_R g3467 ( 
.A(n_3346),
.Y(n_3467)
);

CKINVDCx5p33_ASAP7_75t_R g3468 ( 
.A(n_2987),
.Y(n_3468)
);

CKINVDCx5p33_ASAP7_75t_R g3469 ( 
.A(n_3265),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2739),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3124),
.Y(n_3471)
);

CKINVDCx5p33_ASAP7_75t_R g3472 ( 
.A(n_3268),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_2996),
.Y(n_3473)
);

CKINVDCx5p33_ASAP7_75t_R g3474 ( 
.A(n_3038),
.Y(n_3474)
);

INVxp67_ASAP7_75t_SL g3475 ( 
.A(n_848),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_592),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_1835),
.Y(n_3477)
);

CKINVDCx5p33_ASAP7_75t_R g3478 ( 
.A(n_2367),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_1569),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3195),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3225),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3329),
.Y(n_3482)
);

CKINVDCx5p33_ASAP7_75t_R g3483 ( 
.A(n_703),
.Y(n_3483)
);

CKINVDCx5p33_ASAP7_75t_R g3484 ( 
.A(n_873),
.Y(n_3484)
);

CKINVDCx5p33_ASAP7_75t_R g3485 ( 
.A(n_1804),
.Y(n_3485)
);

CKINVDCx5p33_ASAP7_75t_R g3486 ( 
.A(n_670),
.Y(n_3486)
);

CKINVDCx5p33_ASAP7_75t_R g3487 ( 
.A(n_409),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_1179),
.Y(n_3488)
);

CKINVDCx5p33_ASAP7_75t_R g3489 ( 
.A(n_2516),
.Y(n_3489)
);

CKINVDCx20_ASAP7_75t_R g3490 ( 
.A(n_2468),
.Y(n_3490)
);

CKINVDCx5p33_ASAP7_75t_R g3491 ( 
.A(n_2682),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_1015),
.Y(n_3492)
);

CKINVDCx5p33_ASAP7_75t_R g3493 ( 
.A(n_171),
.Y(n_3493)
);

CKINVDCx5p33_ASAP7_75t_R g3494 ( 
.A(n_3317),
.Y(n_3494)
);

CKINVDCx5p33_ASAP7_75t_R g3495 ( 
.A(n_2670),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_725),
.Y(n_3496)
);

CKINVDCx5p33_ASAP7_75t_R g3497 ( 
.A(n_399),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2421),
.Y(n_3498)
);

CKINVDCx5p33_ASAP7_75t_R g3499 ( 
.A(n_3229),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3013),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_3364),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_199),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_2693),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_477),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_891),
.Y(n_3505)
);

CKINVDCx5p33_ASAP7_75t_R g3506 ( 
.A(n_3312),
.Y(n_3506)
);

CKINVDCx5p33_ASAP7_75t_R g3507 ( 
.A(n_684),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2697),
.Y(n_3508)
);

CKINVDCx5p33_ASAP7_75t_R g3509 ( 
.A(n_3277),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_1764),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_2525),
.Y(n_3511)
);

CKINVDCx5p33_ASAP7_75t_R g3512 ( 
.A(n_83),
.Y(n_3512)
);

CKINVDCx5p33_ASAP7_75t_R g3513 ( 
.A(n_1961),
.Y(n_3513)
);

CKINVDCx5p33_ASAP7_75t_R g3514 ( 
.A(n_1952),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_245),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_2925),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_2132),
.Y(n_3517)
);

CKINVDCx5p33_ASAP7_75t_R g3518 ( 
.A(n_1064),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_2417),
.Y(n_3519)
);

CKINVDCx5p33_ASAP7_75t_R g3520 ( 
.A(n_1530),
.Y(n_3520)
);

CKINVDCx5p33_ASAP7_75t_R g3521 ( 
.A(n_2050),
.Y(n_3521)
);

CKINVDCx5p33_ASAP7_75t_R g3522 ( 
.A(n_3286),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_1927),
.Y(n_3523)
);

BUFx10_ASAP7_75t_L g3524 ( 
.A(n_808),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_347),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_3336),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_3250),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_2148),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_1889),
.Y(n_3529)
);

CKINVDCx5p33_ASAP7_75t_R g3530 ( 
.A(n_141),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2115),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3086),
.Y(n_3532)
);

CKINVDCx5p33_ASAP7_75t_R g3533 ( 
.A(n_2891),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3087),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3331),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_2354),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_2543),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_650),
.Y(n_3538)
);

CKINVDCx5p33_ASAP7_75t_R g3539 ( 
.A(n_836),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_437),
.Y(n_3540)
);

BUFx10_ASAP7_75t_L g3541 ( 
.A(n_2605),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_958),
.Y(n_3542)
);

CKINVDCx5p33_ASAP7_75t_R g3543 ( 
.A(n_1469),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_2569),
.Y(n_3544)
);

CKINVDCx5p33_ASAP7_75t_R g3545 ( 
.A(n_2979),
.Y(n_3545)
);

CKINVDCx5p33_ASAP7_75t_R g3546 ( 
.A(n_2434),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_3171),
.Y(n_3547)
);

CKINVDCx5p33_ASAP7_75t_R g3548 ( 
.A(n_3128),
.Y(n_3548)
);

CKINVDCx5p33_ASAP7_75t_R g3549 ( 
.A(n_47),
.Y(n_3549)
);

CKINVDCx5p33_ASAP7_75t_R g3550 ( 
.A(n_2493),
.Y(n_3550)
);

CKINVDCx5p33_ASAP7_75t_R g3551 ( 
.A(n_1997),
.Y(n_3551)
);

CKINVDCx5p33_ASAP7_75t_R g3552 ( 
.A(n_2776),
.Y(n_3552)
);

CKINVDCx20_ASAP7_75t_R g3553 ( 
.A(n_2767),
.Y(n_3553)
);

CKINVDCx5p33_ASAP7_75t_R g3554 ( 
.A(n_1770),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_821),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_3409),
.Y(n_3556)
);

CKINVDCx5p33_ASAP7_75t_R g3557 ( 
.A(n_2049),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3023),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_3096),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3388),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_77),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_1002),
.Y(n_3562)
);

CKINVDCx5p33_ASAP7_75t_R g3563 ( 
.A(n_114),
.Y(n_3563)
);

INVx1_ASAP7_75t_SL g3564 ( 
.A(n_1962),
.Y(n_3564)
);

CKINVDCx5p33_ASAP7_75t_R g3565 ( 
.A(n_3138),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2006),
.Y(n_3566)
);

BUFx10_ASAP7_75t_L g3567 ( 
.A(n_157),
.Y(n_3567)
);

CKINVDCx5p33_ASAP7_75t_R g3568 ( 
.A(n_2710),
.Y(n_3568)
);

CKINVDCx5p33_ASAP7_75t_R g3569 ( 
.A(n_2707),
.Y(n_3569)
);

CKINVDCx5p33_ASAP7_75t_R g3570 ( 
.A(n_3411),
.Y(n_3570)
);

BUFx5_ASAP7_75t_L g3571 ( 
.A(n_711),
.Y(n_3571)
);

CKINVDCx5p33_ASAP7_75t_R g3572 ( 
.A(n_1412),
.Y(n_3572)
);

CKINVDCx5p33_ASAP7_75t_R g3573 ( 
.A(n_640),
.Y(n_3573)
);

CKINVDCx16_ASAP7_75t_R g3574 ( 
.A(n_2510),
.Y(n_3574)
);

CKINVDCx5p33_ASAP7_75t_R g3575 ( 
.A(n_3334),
.Y(n_3575)
);

INVx1_ASAP7_75t_SL g3576 ( 
.A(n_578),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_935),
.Y(n_3577)
);

BUFx6f_ASAP7_75t_L g3578 ( 
.A(n_1275),
.Y(n_3578)
);

CKINVDCx5p33_ASAP7_75t_R g3579 ( 
.A(n_1031),
.Y(n_3579)
);

CKINVDCx5p33_ASAP7_75t_R g3580 ( 
.A(n_351),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_2904),
.Y(n_3581)
);

CKINVDCx5p33_ASAP7_75t_R g3582 ( 
.A(n_990),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_131),
.Y(n_3583)
);

CKINVDCx5p33_ASAP7_75t_R g3584 ( 
.A(n_2671),
.Y(n_3584)
);

INVx2_ASAP7_75t_SL g3585 ( 
.A(n_2320),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_2165),
.Y(n_3586)
);

CKINVDCx5p33_ASAP7_75t_R g3587 ( 
.A(n_1814),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3281),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3095),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_3413),
.Y(n_3590)
);

CKINVDCx20_ASAP7_75t_R g3591 ( 
.A(n_2146),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3325),
.Y(n_3592)
);

CKINVDCx20_ASAP7_75t_R g3593 ( 
.A(n_631),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_670),
.Y(n_3594)
);

BUFx10_ASAP7_75t_L g3595 ( 
.A(n_3293),
.Y(n_3595)
);

CKINVDCx5p33_ASAP7_75t_R g3596 ( 
.A(n_1772),
.Y(n_3596)
);

BUFx3_ASAP7_75t_L g3597 ( 
.A(n_944),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3421),
.Y(n_3598)
);

CKINVDCx5p33_ASAP7_75t_R g3599 ( 
.A(n_1369),
.Y(n_3599)
);

CKINVDCx5p33_ASAP7_75t_R g3600 ( 
.A(n_378),
.Y(n_3600)
);

INVx1_ASAP7_75t_SL g3601 ( 
.A(n_879),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_1289),
.Y(n_3602)
);

CKINVDCx5p33_ASAP7_75t_R g3603 ( 
.A(n_3264),
.Y(n_3603)
);

CKINVDCx20_ASAP7_75t_R g3604 ( 
.A(n_2080),
.Y(n_3604)
);

CKINVDCx20_ASAP7_75t_R g3605 ( 
.A(n_756),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_2163),
.Y(n_3606)
);

CKINVDCx5p33_ASAP7_75t_R g3607 ( 
.A(n_88),
.Y(n_3607)
);

CKINVDCx5p33_ASAP7_75t_R g3608 ( 
.A(n_83),
.Y(n_3608)
);

BUFx6f_ASAP7_75t_L g3609 ( 
.A(n_3234),
.Y(n_3609)
);

BUFx10_ASAP7_75t_L g3610 ( 
.A(n_1740),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_2952),
.Y(n_3611)
);

BUFx3_ASAP7_75t_L g3612 ( 
.A(n_2020),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_805),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_3258),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_3430),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_3210),
.Y(n_3616)
);

CKINVDCx20_ASAP7_75t_R g3617 ( 
.A(n_1347),
.Y(n_3617)
);

CKINVDCx5p33_ASAP7_75t_R g3618 ( 
.A(n_2619),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_2190),
.Y(n_3619)
);

INVx2_ASAP7_75t_SL g3620 ( 
.A(n_1605),
.Y(n_3620)
);

CKINVDCx5p33_ASAP7_75t_R g3621 ( 
.A(n_375),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_2436),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2618),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3239),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_1757),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_2079),
.Y(n_3626)
);

CKINVDCx5p33_ASAP7_75t_R g3627 ( 
.A(n_3031),
.Y(n_3627)
);

CKINVDCx5p33_ASAP7_75t_R g3628 ( 
.A(n_3069),
.Y(n_3628)
);

INVx1_ASAP7_75t_SL g3629 ( 
.A(n_2380),
.Y(n_3629)
);

CKINVDCx5p33_ASAP7_75t_R g3630 ( 
.A(n_467),
.Y(n_3630)
);

CKINVDCx20_ASAP7_75t_R g3631 ( 
.A(n_1932),
.Y(n_3631)
);

CKINVDCx5p33_ASAP7_75t_R g3632 ( 
.A(n_717),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_1557),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_1345),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3181),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_2664),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_1157),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_821),
.Y(n_3638)
);

CKINVDCx20_ASAP7_75t_R g3639 ( 
.A(n_907),
.Y(n_3639)
);

CKINVDCx5p33_ASAP7_75t_R g3640 ( 
.A(n_1873),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_112),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_3379),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_1385),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_2537),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_1453),
.Y(n_3645)
);

CKINVDCx5p33_ASAP7_75t_R g3646 ( 
.A(n_649),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_3017),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_745),
.Y(n_3648)
);

CKINVDCx5p33_ASAP7_75t_R g3649 ( 
.A(n_3013),
.Y(n_3649)
);

CKINVDCx5p33_ASAP7_75t_R g3650 ( 
.A(n_1701),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_701),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_1444),
.Y(n_3652)
);

CKINVDCx5p33_ASAP7_75t_R g3653 ( 
.A(n_2752),
.Y(n_3653)
);

CKINVDCx5p33_ASAP7_75t_R g3654 ( 
.A(n_597),
.Y(n_3654)
);

CKINVDCx20_ASAP7_75t_R g3655 ( 
.A(n_1254),
.Y(n_3655)
);

CKINVDCx20_ASAP7_75t_R g3656 ( 
.A(n_2529),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_1583),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_2678),
.Y(n_3658)
);

CKINVDCx5p33_ASAP7_75t_R g3659 ( 
.A(n_569),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_3221),
.Y(n_3660)
);

CKINVDCx5p33_ASAP7_75t_R g3661 ( 
.A(n_1027),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_3355),
.Y(n_3662)
);

CKINVDCx5p33_ASAP7_75t_R g3663 ( 
.A(n_2064),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_1683),
.Y(n_3664)
);

CKINVDCx5p33_ASAP7_75t_R g3665 ( 
.A(n_3294),
.Y(n_3665)
);

BUFx2_ASAP7_75t_L g3666 ( 
.A(n_3144),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_2485),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3053),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_3087),
.Y(n_3669)
);

CKINVDCx5p33_ASAP7_75t_R g3670 ( 
.A(n_1594),
.Y(n_3670)
);

HB1xp67_ASAP7_75t_L g3671 ( 
.A(n_2540),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_3298),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_2240),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_1945),
.Y(n_3674)
);

CKINVDCx5p33_ASAP7_75t_R g3675 ( 
.A(n_379),
.Y(n_3675)
);

INVx2_ASAP7_75t_SL g3676 ( 
.A(n_3393),
.Y(n_3676)
);

CKINVDCx5p33_ASAP7_75t_R g3677 ( 
.A(n_2302),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_2073),
.Y(n_3678)
);

CKINVDCx5p33_ASAP7_75t_R g3679 ( 
.A(n_408),
.Y(n_3679)
);

CKINVDCx5p33_ASAP7_75t_R g3680 ( 
.A(n_2165),
.Y(n_3680)
);

BUFx10_ASAP7_75t_L g3681 ( 
.A(n_1704),
.Y(n_3681)
);

CKINVDCx5p33_ASAP7_75t_R g3682 ( 
.A(n_3370),
.Y(n_3682)
);

CKINVDCx5p33_ASAP7_75t_R g3683 ( 
.A(n_1670),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_2820),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_556),
.Y(n_3685)
);

CKINVDCx5p33_ASAP7_75t_R g3686 ( 
.A(n_447),
.Y(n_3686)
);

CKINVDCx5p33_ASAP7_75t_R g3687 ( 
.A(n_305),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_877),
.Y(n_3688)
);

CKINVDCx5p33_ASAP7_75t_R g3689 ( 
.A(n_3103),
.Y(n_3689)
);

CKINVDCx5p33_ASAP7_75t_R g3690 ( 
.A(n_1710),
.Y(n_3690)
);

INVx1_ASAP7_75t_SL g3691 ( 
.A(n_3270),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3296),
.Y(n_3692)
);

BUFx10_ASAP7_75t_L g3693 ( 
.A(n_3392),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_3243),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_1092),
.Y(n_3695)
);

CKINVDCx16_ASAP7_75t_R g3696 ( 
.A(n_928),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_1768),
.Y(n_3697)
);

CKINVDCx5p33_ASAP7_75t_R g3698 ( 
.A(n_581),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_2513),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_1728),
.Y(n_3700)
);

BUFx2_ASAP7_75t_L g3701 ( 
.A(n_671),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_79),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_1096),
.Y(n_3703)
);

CKINVDCx5p33_ASAP7_75t_R g3704 ( 
.A(n_2172),
.Y(n_3704)
);

CKINVDCx5p33_ASAP7_75t_R g3705 ( 
.A(n_849),
.Y(n_3705)
);

INVx2_ASAP7_75t_SL g3706 ( 
.A(n_1665),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3332),
.Y(n_3707)
);

CKINVDCx5p33_ASAP7_75t_R g3708 ( 
.A(n_212),
.Y(n_3708)
);

INVx1_ASAP7_75t_SL g3709 ( 
.A(n_1086),
.Y(n_3709)
);

CKINVDCx20_ASAP7_75t_R g3710 ( 
.A(n_1230),
.Y(n_3710)
);

CKINVDCx5p33_ASAP7_75t_R g3711 ( 
.A(n_2172),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_2146),
.Y(n_3712)
);

CKINVDCx14_ASAP7_75t_R g3713 ( 
.A(n_261),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_2479),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_734),
.Y(n_3715)
);

CKINVDCx5p33_ASAP7_75t_R g3716 ( 
.A(n_3386),
.Y(n_3716)
);

INVx2_ASAP7_75t_SL g3717 ( 
.A(n_417),
.Y(n_3717)
);

CKINVDCx5p33_ASAP7_75t_R g3718 ( 
.A(n_3406),
.Y(n_3718)
);

HB1xp67_ASAP7_75t_L g3719 ( 
.A(n_2419),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_58),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3078),
.Y(n_3721)
);

CKINVDCx5p33_ASAP7_75t_R g3722 ( 
.A(n_3356),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_1697),
.Y(n_3723)
);

CKINVDCx5p33_ASAP7_75t_R g3724 ( 
.A(n_3374),
.Y(n_3724)
);

CKINVDCx5p33_ASAP7_75t_R g3725 ( 
.A(n_1906),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_2686),
.Y(n_3726)
);

BUFx3_ASAP7_75t_L g3727 ( 
.A(n_2120),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_880),
.Y(n_3728)
);

BUFx10_ASAP7_75t_L g3729 ( 
.A(n_799),
.Y(n_3729)
);

CKINVDCx5p33_ASAP7_75t_R g3730 ( 
.A(n_1346),
.Y(n_3730)
);

CKINVDCx5p33_ASAP7_75t_R g3731 ( 
.A(n_267),
.Y(n_3731)
);

CKINVDCx5p33_ASAP7_75t_R g3732 ( 
.A(n_1037),
.Y(n_3732)
);

CKINVDCx5p33_ASAP7_75t_R g3733 ( 
.A(n_1388),
.Y(n_3733)
);

CKINVDCx5p33_ASAP7_75t_R g3734 ( 
.A(n_3282),
.Y(n_3734)
);

CKINVDCx5p33_ASAP7_75t_R g3735 ( 
.A(n_2445),
.Y(n_3735)
);

CKINVDCx16_ASAP7_75t_R g3736 ( 
.A(n_3422),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_1312),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_2063),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_662),
.Y(n_3739)
);

CKINVDCx5p33_ASAP7_75t_R g3740 ( 
.A(n_3258),
.Y(n_3740)
);

CKINVDCx5p33_ASAP7_75t_R g3741 ( 
.A(n_2791),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_2253),
.Y(n_3742)
);

CKINVDCx5p33_ASAP7_75t_R g3743 ( 
.A(n_3316),
.Y(n_3743)
);

BUFx10_ASAP7_75t_L g3744 ( 
.A(n_3373),
.Y(n_3744)
);

CKINVDCx20_ASAP7_75t_R g3745 ( 
.A(n_2746),
.Y(n_3745)
);

CKINVDCx5p33_ASAP7_75t_R g3746 ( 
.A(n_2014),
.Y(n_3746)
);

CKINVDCx20_ASAP7_75t_R g3747 ( 
.A(n_2183),
.Y(n_3747)
);

CKINVDCx20_ASAP7_75t_R g3748 ( 
.A(n_528),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_3231),
.Y(n_3749)
);

CKINVDCx5p33_ASAP7_75t_R g3750 ( 
.A(n_2070),
.Y(n_3750)
);

CKINVDCx5p33_ASAP7_75t_R g3751 ( 
.A(n_3410),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_880),
.Y(n_3752)
);

CKINVDCx5p33_ASAP7_75t_R g3753 ( 
.A(n_873),
.Y(n_3753)
);

CKINVDCx5p33_ASAP7_75t_R g3754 ( 
.A(n_3368),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_2300),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3233),
.Y(n_3756)
);

BUFx10_ASAP7_75t_L g3757 ( 
.A(n_1198),
.Y(n_3757)
);

CKINVDCx5p33_ASAP7_75t_R g3758 ( 
.A(n_109),
.Y(n_3758)
);

CKINVDCx5p33_ASAP7_75t_R g3759 ( 
.A(n_1252),
.Y(n_3759)
);

CKINVDCx5p33_ASAP7_75t_R g3760 ( 
.A(n_1141),
.Y(n_3760)
);

CKINVDCx5p33_ASAP7_75t_R g3761 ( 
.A(n_2770),
.Y(n_3761)
);

BUFx5_ASAP7_75t_L g3762 ( 
.A(n_2748),
.Y(n_3762)
);

CKINVDCx5p33_ASAP7_75t_R g3763 ( 
.A(n_982),
.Y(n_3763)
);

CKINVDCx20_ASAP7_75t_R g3764 ( 
.A(n_228),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_1119),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_2320),
.Y(n_3766)
);

CKINVDCx5p33_ASAP7_75t_R g3767 ( 
.A(n_478),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_2477),
.Y(n_3768)
);

CKINVDCx5p33_ASAP7_75t_R g3769 ( 
.A(n_2075),
.Y(n_3769)
);

CKINVDCx5p33_ASAP7_75t_R g3770 ( 
.A(n_1062),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_1561),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_1007),
.Y(n_3772)
);

CKINVDCx5p33_ASAP7_75t_R g3773 ( 
.A(n_759),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_1396),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_2837),
.Y(n_3775)
);

CKINVDCx14_ASAP7_75t_R g3776 ( 
.A(n_3082),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_1489),
.Y(n_3777)
);

INVx1_ASAP7_75t_SL g3778 ( 
.A(n_928),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_1732),
.Y(n_3779)
);

CKINVDCx5p33_ASAP7_75t_R g3780 ( 
.A(n_1681),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3119),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_913),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_1099),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_1271),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3460),
.Y(n_3785)
);

CKINVDCx5p33_ASAP7_75t_R g3786 ( 
.A(n_3235),
.Y(n_3786)
);

INVx2_ASAP7_75t_SL g3787 ( 
.A(n_1198),
.Y(n_3787)
);

CKINVDCx5p33_ASAP7_75t_R g3788 ( 
.A(n_1539),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_1581),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_277),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3256),
.Y(n_3791)
);

CKINVDCx5p33_ASAP7_75t_R g3792 ( 
.A(n_2516),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_343),
.Y(n_3793)
);

BUFx8_ASAP7_75t_SL g3794 ( 
.A(n_2491),
.Y(n_3794)
);

CKINVDCx5p33_ASAP7_75t_R g3795 ( 
.A(n_825),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3287),
.Y(n_3796)
);

CKINVDCx5p33_ASAP7_75t_R g3797 ( 
.A(n_1788),
.Y(n_3797)
);

BUFx10_ASAP7_75t_L g3798 ( 
.A(n_809),
.Y(n_3798)
);

CKINVDCx5p33_ASAP7_75t_R g3799 ( 
.A(n_3404),
.Y(n_3799)
);

CKINVDCx5p33_ASAP7_75t_R g3800 ( 
.A(n_1400),
.Y(n_3800)
);

CKINVDCx5p33_ASAP7_75t_R g3801 ( 
.A(n_442),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_2367),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_233),
.Y(n_3803)
);

BUFx3_ASAP7_75t_L g3804 ( 
.A(n_437),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3237),
.Y(n_3805)
);

CKINVDCx5p33_ASAP7_75t_R g3806 ( 
.A(n_701),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3310),
.Y(n_3807)
);

CKINVDCx5p33_ASAP7_75t_R g3808 ( 
.A(n_1371),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3241),
.Y(n_3809)
);

BUFx10_ASAP7_75t_L g3810 ( 
.A(n_1969),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_946),
.Y(n_3811)
);

CKINVDCx5p33_ASAP7_75t_R g3812 ( 
.A(n_2591),
.Y(n_3812)
);

CKINVDCx5p33_ASAP7_75t_R g3813 ( 
.A(n_3257),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_1649),
.Y(n_3814)
);

BUFx6f_ASAP7_75t_L g3815 ( 
.A(n_1241),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_337),
.Y(n_3816)
);

CKINVDCx5p33_ASAP7_75t_R g3817 ( 
.A(n_1971),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_1210),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_2519),
.Y(n_3819)
);

CKINVDCx5p33_ASAP7_75t_R g3820 ( 
.A(n_3251),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_1754),
.Y(n_3821)
);

CKINVDCx5p33_ASAP7_75t_R g3822 ( 
.A(n_2569),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_2537),
.Y(n_3823)
);

CKINVDCx5p33_ASAP7_75t_R g3824 ( 
.A(n_3399),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3365),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_1926),
.Y(n_3826)
);

CKINVDCx20_ASAP7_75t_R g3827 ( 
.A(n_1538),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_3262),
.Y(n_3828)
);

HB1xp67_ASAP7_75t_L g3829 ( 
.A(n_2030),
.Y(n_3829)
);

CKINVDCx20_ASAP7_75t_R g3830 ( 
.A(n_3349),
.Y(n_3830)
);

CKINVDCx5p33_ASAP7_75t_R g3831 ( 
.A(n_2753),
.Y(n_3831)
);

CKINVDCx5p33_ASAP7_75t_R g3832 ( 
.A(n_2939),
.Y(n_3832)
);

CKINVDCx5p33_ASAP7_75t_R g3833 ( 
.A(n_240),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_525),
.Y(n_3834)
);

CKINVDCx5p33_ASAP7_75t_R g3835 ( 
.A(n_2423),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_1917),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_1999),
.Y(n_3837)
);

CKINVDCx5p33_ASAP7_75t_R g3838 ( 
.A(n_3305),
.Y(n_3838)
);

CKINVDCx5p33_ASAP7_75t_R g3839 ( 
.A(n_667),
.Y(n_3839)
);

CKINVDCx5p33_ASAP7_75t_R g3840 ( 
.A(n_113),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_1297),
.Y(n_3841)
);

CKINVDCx5p33_ASAP7_75t_R g3842 ( 
.A(n_1668),
.Y(n_3842)
);

BUFx2_ASAP7_75t_SL g3843 ( 
.A(n_3267),
.Y(n_3843)
);

INVx1_ASAP7_75t_SL g3844 ( 
.A(n_1981),
.Y(n_3844)
);

INVx1_ASAP7_75t_SL g3845 ( 
.A(n_3248),
.Y(n_3845)
);

INVx2_ASAP7_75t_SL g3846 ( 
.A(n_1746),
.Y(n_3846)
);

BUFx6f_ASAP7_75t_L g3847 ( 
.A(n_576),
.Y(n_3847)
);

CKINVDCx5p33_ASAP7_75t_R g3848 ( 
.A(n_680),
.Y(n_3848)
);

INVx1_ASAP7_75t_SL g3849 ( 
.A(n_3441),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_740),
.Y(n_3850)
);

CKINVDCx5p33_ASAP7_75t_R g3851 ( 
.A(n_3019),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_2358),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2708),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3363),
.Y(n_3854)
);

HB1xp67_ASAP7_75t_L g3855 ( 
.A(n_2022),
.Y(n_3855)
);

CKINVDCx5p33_ASAP7_75t_R g3856 ( 
.A(n_3207),
.Y(n_3856)
);

HB1xp67_ASAP7_75t_L g3857 ( 
.A(n_2788),
.Y(n_3857)
);

CKINVDCx5p33_ASAP7_75t_R g3858 ( 
.A(n_2100),
.Y(n_3858)
);

CKINVDCx5p33_ASAP7_75t_R g3859 ( 
.A(n_2327),
.Y(n_3859)
);

CKINVDCx5p33_ASAP7_75t_R g3860 ( 
.A(n_3326),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_2148),
.Y(n_3861)
);

CKINVDCx5p33_ASAP7_75t_R g3862 ( 
.A(n_1244),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_404),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_1775),
.Y(n_3864)
);

BUFx10_ASAP7_75t_L g3865 ( 
.A(n_838),
.Y(n_3865)
);

CKINVDCx5p33_ASAP7_75t_R g3866 ( 
.A(n_3279),
.Y(n_3866)
);

CKINVDCx5p33_ASAP7_75t_R g3867 ( 
.A(n_1534),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_2642),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_517),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_2951),
.Y(n_3870)
);

CKINVDCx5p33_ASAP7_75t_R g3871 ( 
.A(n_301),
.Y(n_3871)
);

CKINVDCx5p33_ASAP7_75t_R g3872 ( 
.A(n_2317),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_707),
.Y(n_3873)
);

BUFx3_ASAP7_75t_L g3874 ( 
.A(n_908),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3191),
.Y(n_3875)
);

CKINVDCx5p33_ASAP7_75t_R g3876 ( 
.A(n_3390),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_1915),
.Y(n_3877)
);

CKINVDCx5p33_ASAP7_75t_R g3878 ( 
.A(n_149),
.Y(n_3878)
);

CKINVDCx5p33_ASAP7_75t_R g3879 ( 
.A(n_368),
.Y(n_3879)
);

CKINVDCx5p33_ASAP7_75t_R g3880 ( 
.A(n_248),
.Y(n_3880)
);

CKINVDCx5p33_ASAP7_75t_R g3881 ( 
.A(n_2944),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_111),
.Y(n_3882)
);

BUFx3_ASAP7_75t_L g3883 ( 
.A(n_2422),
.Y(n_3883)
);

CKINVDCx5p33_ASAP7_75t_R g3884 ( 
.A(n_3274),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_177),
.Y(n_3885)
);

CKINVDCx5p33_ASAP7_75t_R g3886 ( 
.A(n_3133),
.Y(n_3886)
);

CKINVDCx5p33_ASAP7_75t_R g3887 ( 
.A(n_385),
.Y(n_3887)
);

CKINVDCx20_ASAP7_75t_R g3888 ( 
.A(n_2939),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_3397),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_2883),
.Y(n_3890)
);

INVx2_ASAP7_75t_SL g3891 ( 
.A(n_2770),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3254),
.Y(n_3892)
);

CKINVDCx5p33_ASAP7_75t_R g3893 ( 
.A(n_347),
.Y(n_3893)
);

CKINVDCx5p33_ASAP7_75t_R g3894 ( 
.A(n_2871),
.Y(n_3894)
);

CKINVDCx5p33_ASAP7_75t_R g3895 ( 
.A(n_1666),
.Y(n_3895)
);

CKINVDCx5p33_ASAP7_75t_R g3896 ( 
.A(n_3432),
.Y(n_3896)
);

CKINVDCx5p33_ASAP7_75t_R g3897 ( 
.A(n_2055),
.Y(n_3897)
);

CKINVDCx5p33_ASAP7_75t_R g3898 ( 
.A(n_2773),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3249),
.Y(n_3899)
);

CKINVDCx5p33_ASAP7_75t_R g3900 ( 
.A(n_1812),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_2364),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3259),
.Y(n_3902)
);

CKINVDCx20_ASAP7_75t_R g3903 ( 
.A(n_92),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_274),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_1779),
.Y(n_3905)
);

CKINVDCx5p33_ASAP7_75t_R g3906 ( 
.A(n_2861),
.Y(n_3906)
);

CKINVDCx20_ASAP7_75t_R g3907 ( 
.A(n_2451),
.Y(n_3907)
);

CKINVDCx5p33_ASAP7_75t_R g3908 ( 
.A(n_499),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_1943),
.Y(n_3909)
);

CKINVDCx5p33_ASAP7_75t_R g3910 ( 
.A(n_466),
.Y(n_3910)
);

CKINVDCx5p33_ASAP7_75t_R g3911 ( 
.A(n_2064),
.Y(n_3911)
);

CKINVDCx5p33_ASAP7_75t_R g3912 ( 
.A(n_2126),
.Y(n_3912)
);

CKINVDCx20_ASAP7_75t_R g3913 ( 
.A(n_3436),
.Y(n_3913)
);

CKINVDCx16_ASAP7_75t_R g3914 ( 
.A(n_2355),
.Y(n_3914)
);

INVxp67_ASAP7_75t_L g3915 ( 
.A(n_203),
.Y(n_3915)
);

CKINVDCx5p33_ASAP7_75t_R g3916 ( 
.A(n_3432),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3345),
.Y(n_3917)
);

BUFx10_ASAP7_75t_L g3918 ( 
.A(n_2660),
.Y(n_3918)
);

CKINVDCx5p33_ASAP7_75t_R g3919 ( 
.A(n_1251),
.Y(n_3919)
);

CKINVDCx5p33_ASAP7_75t_R g3920 ( 
.A(n_2763),
.Y(n_3920)
);

CKINVDCx5p33_ASAP7_75t_R g3921 ( 
.A(n_622),
.Y(n_3921)
);

CKINVDCx5p33_ASAP7_75t_R g3922 ( 
.A(n_1275),
.Y(n_3922)
);

BUFx10_ASAP7_75t_L g3923 ( 
.A(n_2089),
.Y(n_3923)
);

CKINVDCx5p33_ASAP7_75t_R g3924 ( 
.A(n_1332),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_3402),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_1146),
.Y(n_3926)
);

CKINVDCx5p33_ASAP7_75t_R g3927 ( 
.A(n_56),
.Y(n_3927)
);

BUFx6f_ASAP7_75t_L g3928 ( 
.A(n_2616),
.Y(n_3928)
);

CKINVDCx5p33_ASAP7_75t_R g3929 ( 
.A(n_3012),
.Y(n_3929)
);

BUFx3_ASAP7_75t_L g3930 ( 
.A(n_2752),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_1614),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_1103),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3339),
.Y(n_3933)
);

CKINVDCx5p33_ASAP7_75t_R g3934 ( 
.A(n_1450),
.Y(n_3934)
);

CKINVDCx5p33_ASAP7_75t_R g3935 ( 
.A(n_2125),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_1038),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_2282),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_363),
.Y(n_3938)
);

CKINVDCx5p33_ASAP7_75t_R g3939 ( 
.A(n_122),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_1095),
.Y(n_3940)
);

BUFx6f_ASAP7_75t_L g3941 ( 
.A(n_1624),
.Y(n_3941)
);

CKINVDCx5p33_ASAP7_75t_R g3942 ( 
.A(n_422),
.Y(n_3942)
);

CKINVDCx5p33_ASAP7_75t_R g3943 ( 
.A(n_314),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_1879),
.Y(n_3944)
);

CKINVDCx5p33_ASAP7_75t_R g3945 ( 
.A(n_3383),
.Y(n_3945)
);

CKINVDCx5p33_ASAP7_75t_R g3946 ( 
.A(n_3007),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_213),
.Y(n_3947)
);

CKINVDCx5p33_ASAP7_75t_R g3948 ( 
.A(n_465),
.Y(n_3948)
);

CKINVDCx5p33_ASAP7_75t_R g3949 ( 
.A(n_2319),
.Y(n_3949)
);

CKINVDCx5p33_ASAP7_75t_R g3950 ( 
.A(n_3415),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_479),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_2549),
.Y(n_3952)
);

CKINVDCx14_ASAP7_75t_R g3953 ( 
.A(n_2905),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_2748),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_1796),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_1195),
.Y(n_3956)
);

BUFx6f_ASAP7_75t_L g3957 ( 
.A(n_2614),
.Y(n_3957)
);

CKINVDCx5p33_ASAP7_75t_R g3958 ( 
.A(n_1410),
.Y(n_3958)
);

CKINVDCx20_ASAP7_75t_R g3959 ( 
.A(n_3315),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3425),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_1242),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_2373),
.Y(n_3962)
);

INVx2_ASAP7_75t_SL g3963 ( 
.A(n_2636),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_176),
.Y(n_3964)
);

CKINVDCx20_ASAP7_75t_R g3965 ( 
.A(n_2144),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_822),
.Y(n_3966)
);

CKINVDCx5p33_ASAP7_75t_R g3967 ( 
.A(n_1433),
.Y(n_3967)
);

CKINVDCx5p33_ASAP7_75t_R g3968 ( 
.A(n_98),
.Y(n_3968)
);

CKINVDCx5p33_ASAP7_75t_R g3969 ( 
.A(n_3046),
.Y(n_3969)
);

CKINVDCx5p33_ASAP7_75t_R g3970 ( 
.A(n_3082),
.Y(n_3970)
);

CKINVDCx5p33_ASAP7_75t_R g3971 ( 
.A(n_2964),
.Y(n_3971)
);

CKINVDCx5p33_ASAP7_75t_R g3972 ( 
.A(n_1740),
.Y(n_3972)
);

CKINVDCx5p33_ASAP7_75t_R g3973 ( 
.A(n_2954),
.Y(n_3973)
);

CKINVDCx5p33_ASAP7_75t_R g3974 ( 
.A(n_3268),
.Y(n_3974)
);

BUFx10_ASAP7_75t_L g3975 ( 
.A(n_2045),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_1641),
.Y(n_3976)
);

CKINVDCx5p33_ASAP7_75t_R g3977 ( 
.A(n_1994),
.Y(n_3977)
);

BUFx6f_ASAP7_75t_L g3978 ( 
.A(n_3196),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_916),
.Y(n_3979)
);

CKINVDCx20_ASAP7_75t_R g3980 ( 
.A(n_2217),
.Y(n_3980)
);

CKINVDCx5p33_ASAP7_75t_R g3981 ( 
.A(n_3355),
.Y(n_3981)
);

CKINVDCx5p33_ASAP7_75t_R g3982 ( 
.A(n_2566),
.Y(n_3982)
);

CKINVDCx5p33_ASAP7_75t_R g3983 ( 
.A(n_3260),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_1691),
.Y(n_3984)
);

CKINVDCx5p33_ASAP7_75t_R g3985 ( 
.A(n_812),
.Y(n_3985)
);

CKINVDCx5p33_ASAP7_75t_R g3986 ( 
.A(n_165),
.Y(n_3986)
);

CKINVDCx5p33_ASAP7_75t_R g3987 ( 
.A(n_1886),
.Y(n_3987)
);

CKINVDCx5p33_ASAP7_75t_R g3988 ( 
.A(n_3220),
.Y(n_3988)
);

CKINVDCx5p33_ASAP7_75t_R g3989 ( 
.A(n_1725),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_392),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_1551),
.Y(n_3991)
);

BUFx10_ASAP7_75t_L g3992 ( 
.A(n_3397),
.Y(n_3992)
);

BUFx10_ASAP7_75t_L g3993 ( 
.A(n_2302),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_3340),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_850),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3344),
.Y(n_3996)
);

CKINVDCx5p33_ASAP7_75t_R g3997 ( 
.A(n_246),
.Y(n_3997)
);

CKINVDCx5p33_ASAP7_75t_R g3998 ( 
.A(n_1717),
.Y(n_3998)
);

BUFx3_ASAP7_75t_L g3999 ( 
.A(n_178),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_1006),
.Y(n_4000)
);

CKINVDCx5p33_ASAP7_75t_R g4001 ( 
.A(n_1552),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_758),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_1128),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_2246),
.Y(n_4004)
);

CKINVDCx5p33_ASAP7_75t_R g4005 ( 
.A(n_1097),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_3047),
.Y(n_4006)
);

CKINVDCx5p33_ASAP7_75t_R g4007 ( 
.A(n_59),
.Y(n_4007)
);

CKINVDCx5p33_ASAP7_75t_R g4008 ( 
.A(n_3193),
.Y(n_4008)
);

BUFx10_ASAP7_75t_L g4009 ( 
.A(n_2550),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_718),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_2233),
.Y(n_4011)
);

CKINVDCx14_ASAP7_75t_R g4012 ( 
.A(n_2977),
.Y(n_4012)
);

BUFx6f_ASAP7_75t_L g4013 ( 
.A(n_210),
.Y(n_4013)
);

INVx1_ASAP7_75t_SL g4014 ( 
.A(n_2234),
.Y(n_4014)
);

CKINVDCx5p33_ASAP7_75t_R g4015 ( 
.A(n_1698),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3285),
.Y(n_4016)
);

CKINVDCx20_ASAP7_75t_R g4017 ( 
.A(n_1949),
.Y(n_4017)
);

CKINVDCx5p33_ASAP7_75t_R g4018 ( 
.A(n_1632),
.Y(n_4018)
);

CKINVDCx5p33_ASAP7_75t_R g4019 ( 
.A(n_3378),
.Y(n_4019)
);

CKINVDCx5p33_ASAP7_75t_R g4020 ( 
.A(n_2975),
.Y(n_4020)
);

CKINVDCx5p33_ASAP7_75t_R g4021 ( 
.A(n_1187),
.Y(n_4021)
);

CKINVDCx5p33_ASAP7_75t_R g4022 ( 
.A(n_1968),
.Y(n_4022)
);

CKINVDCx5p33_ASAP7_75t_R g4023 ( 
.A(n_1371),
.Y(n_4023)
);

CKINVDCx20_ASAP7_75t_R g4024 ( 
.A(n_3171),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3341),
.Y(n_4025)
);

CKINVDCx5p33_ASAP7_75t_R g4026 ( 
.A(n_2638),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3403),
.Y(n_4027)
);

BUFx8_ASAP7_75t_SL g4028 ( 
.A(n_1621),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_1313),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_2838),
.Y(n_4030)
);

CKINVDCx5p33_ASAP7_75t_R g4031 ( 
.A(n_3321),
.Y(n_4031)
);

CKINVDCx20_ASAP7_75t_R g4032 ( 
.A(n_1907),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_2394),
.Y(n_4033)
);

CKINVDCx5p33_ASAP7_75t_R g4034 ( 
.A(n_599),
.Y(n_4034)
);

BUFx6f_ASAP7_75t_L g4035 ( 
.A(n_1151),
.Y(n_4035)
);

CKINVDCx5p33_ASAP7_75t_R g4036 ( 
.A(n_1495),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_1628),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_929),
.Y(n_4038)
);

CKINVDCx5p33_ASAP7_75t_R g4039 ( 
.A(n_1850),
.Y(n_4039)
);

CKINVDCx5p33_ASAP7_75t_R g4040 ( 
.A(n_919),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_1624),
.Y(n_4041)
);

CKINVDCx5p33_ASAP7_75t_R g4042 ( 
.A(n_1287),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_1886),
.Y(n_4043)
);

INVx2_ASAP7_75t_SL g4044 ( 
.A(n_960),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_422),
.Y(n_4045)
);

CKINVDCx5p33_ASAP7_75t_R g4046 ( 
.A(n_34),
.Y(n_4046)
);

CKINVDCx5p33_ASAP7_75t_R g4047 ( 
.A(n_1767),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_2450),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_2618),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_2887),
.Y(n_4050)
);

CKINVDCx5p33_ASAP7_75t_R g4051 ( 
.A(n_2343),
.Y(n_4051)
);

CKINVDCx20_ASAP7_75t_R g4052 ( 
.A(n_610),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_2324),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_1889),
.Y(n_4054)
);

CKINVDCx5p33_ASAP7_75t_R g4055 ( 
.A(n_1028),
.Y(n_4055)
);

CKINVDCx20_ASAP7_75t_R g4056 ( 
.A(n_2556),
.Y(n_4056)
);

CKINVDCx5p33_ASAP7_75t_R g4057 ( 
.A(n_2371),
.Y(n_4057)
);

INVxp67_ASAP7_75t_SL g4058 ( 
.A(n_1506),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3340),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_172),
.Y(n_4060)
);

CKINVDCx5p33_ASAP7_75t_R g4061 ( 
.A(n_3453),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_944),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_2123),
.Y(n_4063)
);

BUFx6f_ASAP7_75t_L g4064 ( 
.A(n_1953),
.Y(n_4064)
);

BUFx10_ASAP7_75t_L g4065 ( 
.A(n_1030),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_2384),
.Y(n_4066)
);

CKINVDCx5p33_ASAP7_75t_R g4067 ( 
.A(n_472),
.Y(n_4067)
);

CKINVDCx5p33_ASAP7_75t_R g4068 ( 
.A(n_1931),
.Y(n_4068)
);

CKINVDCx5p33_ASAP7_75t_R g4069 ( 
.A(n_1238),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_1762),
.Y(n_4070)
);

CKINVDCx5p33_ASAP7_75t_R g4071 ( 
.A(n_1883),
.Y(n_4071)
);

BUFx10_ASAP7_75t_L g4072 ( 
.A(n_1494),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_1368),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_2439),
.Y(n_4074)
);

CKINVDCx5p33_ASAP7_75t_R g4075 ( 
.A(n_510),
.Y(n_4075)
);

CKINVDCx5p33_ASAP7_75t_R g4076 ( 
.A(n_2104),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3190),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_407),
.Y(n_4078)
);

CKINVDCx5p33_ASAP7_75t_R g4079 ( 
.A(n_3433),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_2529),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3183),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_2004),
.Y(n_4082)
);

CKINVDCx5p33_ASAP7_75t_R g4083 ( 
.A(n_1300),
.Y(n_4083)
);

CKINVDCx20_ASAP7_75t_R g4084 ( 
.A(n_3207),
.Y(n_4084)
);

CKINVDCx5p33_ASAP7_75t_R g4085 ( 
.A(n_1023),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_1026),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_283),
.Y(n_4087)
);

CKINVDCx5p33_ASAP7_75t_R g4088 ( 
.A(n_1087),
.Y(n_4088)
);

CKINVDCx5p33_ASAP7_75t_R g4089 ( 
.A(n_1585),
.Y(n_4089)
);

CKINVDCx5p33_ASAP7_75t_R g4090 ( 
.A(n_3128),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_1062),
.Y(n_4091)
);

CKINVDCx5p33_ASAP7_75t_R g4092 ( 
.A(n_1212),
.Y(n_4092)
);

BUFx10_ASAP7_75t_L g4093 ( 
.A(n_1686),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_2634),
.Y(n_4094)
);

CKINVDCx5p33_ASAP7_75t_R g4095 ( 
.A(n_3227),
.Y(n_4095)
);

CKINVDCx5p33_ASAP7_75t_R g4096 ( 
.A(n_176),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_1576),
.Y(n_4097)
);

HB1xp67_ASAP7_75t_L g4098 ( 
.A(n_1678),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_853),
.Y(n_4099)
);

CKINVDCx5p33_ASAP7_75t_R g4100 ( 
.A(n_3378),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_144),
.Y(n_4101)
);

BUFx5_ASAP7_75t_L g4102 ( 
.A(n_2207),
.Y(n_4102)
);

CKINVDCx5p33_ASAP7_75t_R g4103 ( 
.A(n_3211),
.Y(n_4103)
);

CKINVDCx5p33_ASAP7_75t_R g4104 ( 
.A(n_410),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_154),
.Y(n_4105)
);

CKINVDCx20_ASAP7_75t_R g4106 ( 
.A(n_438),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_985),
.Y(n_4107)
);

CKINVDCx16_ASAP7_75t_R g4108 ( 
.A(n_3113),
.Y(n_4108)
);

BUFx6f_ASAP7_75t_L g4109 ( 
.A(n_1388),
.Y(n_4109)
);

CKINVDCx16_ASAP7_75t_R g4110 ( 
.A(n_3371),
.Y(n_4110)
);

INVx2_ASAP7_75t_SL g4111 ( 
.A(n_1476),
.Y(n_4111)
);

CKINVDCx5p33_ASAP7_75t_R g4112 ( 
.A(n_2433),
.Y(n_4112)
);

CKINVDCx20_ASAP7_75t_R g4113 ( 
.A(n_1231),
.Y(n_4113)
);

CKINVDCx5p33_ASAP7_75t_R g4114 ( 
.A(n_3382),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_306),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_1748),
.Y(n_4116)
);

CKINVDCx5p33_ASAP7_75t_R g4117 ( 
.A(n_2791),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_2921),
.Y(n_4118)
);

CKINVDCx5p33_ASAP7_75t_R g4119 ( 
.A(n_876),
.Y(n_4119)
);

CKINVDCx5p33_ASAP7_75t_R g4120 ( 
.A(n_2573),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_2705),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_1695),
.Y(n_4122)
);

CKINVDCx20_ASAP7_75t_R g4123 ( 
.A(n_3051),
.Y(n_4123)
);

CKINVDCx16_ASAP7_75t_R g4124 ( 
.A(n_630),
.Y(n_4124)
);

BUFx10_ASAP7_75t_L g4125 ( 
.A(n_3031),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_2775),
.Y(n_4126)
);

CKINVDCx16_ASAP7_75t_R g4127 ( 
.A(n_3283),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_1954),
.Y(n_4128)
);

CKINVDCx5p33_ASAP7_75t_R g4129 ( 
.A(n_2948),
.Y(n_4129)
);

INVx1_ASAP7_75t_SL g4130 ( 
.A(n_1898),
.Y(n_4130)
);

CKINVDCx5p33_ASAP7_75t_R g4131 ( 
.A(n_302),
.Y(n_4131)
);

CKINVDCx5p33_ASAP7_75t_R g4132 ( 
.A(n_334),
.Y(n_4132)
);

CKINVDCx20_ASAP7_75t_R g4133 ( 
.A(n_2642),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_2183),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_3389),
.Y(n_4135)
);

CKINVDCx5p33_ASAP7_75t_R g4136 ( 
.A(n_571),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_371),
.Y(n_4137)
);

BUFx6f_ASAP7_75t_L g4138 ( 
.A(n_352),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_1495),
.Y(n_4139)
);

CKINVDCx5p33_ASAP7_75t_R g4140 ( 
.A(n_387),
.Y(n_4140)
);

INVx2_ASAP7_75t_SL g4141 ( 
.A(n_917),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_1257),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_3351),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_1949),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_1722),
.Y(n_4145)
);

BUFx6f_ASAP7_75t_L g4146 ( 
.A(n_2671),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_304),
.Y(n_4147)
);

CKINVDCx5p33_ASAP7_75t_R g4148 ( 
.A(n_3244),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_1277),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_913),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_2850),
.Y(n_4151)
);

CKINVDCx5p33_ASAP7_75t_R g4152 ( 
.A(n_1678),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_422),
.Y(n_4153)
);

CKINVDCx5p33_ASAP7_75t_R g4154 ( 
.A(n_1625),
.Y(n_4154)
);

CKINVDCx5p33_ASAP7_75t_R g4155 ( 
.A(n_3292),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_1928),
.Y(n_4156)
);

INVx2_ASAP7_75t_SL g4157 ( 
.A(n_3181),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_3314),
.Y(n_4158)
);

CKINVDCx5p33_ASAP7_75t_R g4159 ( 
.A(n_894),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3284),
.Y(n_4160)
);

BUFx6f_ASAP7_75t_L g4161 ( 
.A(n_2985),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_2531),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_1343),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_1793),
.Y(n_4164)
);

CKINVDCx5p33_ASAP7_75t_R g4165 ( 
.A(n_516),
.Y(n_4165)
);

CKINVDCx5p33_ASAP7_75t_R g4166 ( 
.A(n_2037),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_159),
.Y(n_4167)
);

CKINVDCx20_ASAP7_75t_R g4168 ( 
.A(n_1506),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_1429),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_2118),
.Y(n_4170)
);

CKINVDCx20_ASAP7_75t_R g4171 ( 
.A(n_122),
.Y(n_4171)
);

CKINVDCx5p33_ASAP7_75t_R g4172 ( 
.A(n_674),
.Y(n_4172)
);

CKINVDCx5p33_ASAP7_75t_R g4173 ( 
.A(n_764),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_308),
.Y(n_4174)
);

CKINVDCx5p33_ASAP7_75t_R g4175 ( 
.A(n_2513),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3225),
.Y(n_4176)
);

HB1xp67_ASAP7_75t_L g4177 ( 
.A(n_1542),
.Y(n_4177)
);

INVx1_ASAP7_75t_SL g4178 ( 
.A(n_366),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_1747),
.Y(n_4179)
);

CKINVDCx5p33_ASAP7_75t_R g4180 ( 
.A(n_2106),
.Y(n_4180)
);

CKINVDCx5p33_ASAP7_75t_R g4181 ( 
.A(n_72),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_1269),
.Y(n_4182)
);

CKINVDCx5p33_ASAP7_75t_R g4183 ( 
.A(n_2928),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3276),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_1384),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3141),
.Y(n_4186)
);

BUFx10_ASAP7_75t_L g4187 ( 
.A(n_1342),
.Y(n_4187)
);

CKINVDCx5p33_ASAP7_75t_R g4188 ( 
.A(n_3308),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3263),
.Y(n_4189)
);

BUFx6f_ASAP7_75t_L g4190 ( 
.A(n_1133),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_1087),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3306),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_2300),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_3271),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_908),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_2443),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_1510),
.Y(n_4197)
);

CKINVDCx5p33_ASAP7_75t_R g4198 ( 
.A(n_545),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_831),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3330),
.Y(n_4200)
);

INVx1_ASAP7_75t_SL g4201 ( 
.A(n_1672),
.Y(n_4201)
);

BUFx2_ASAP7_75t_L g4202 ( 
.A(n_3327),
.Y(n_4202)
);

CKINVDCx5p33_ASAP7_75t_R g4203 ( 
.A(n_3395),
.Y(n_4203)
);

CKINVDCx5p33_ASAP7_75t_R g4204 ( 
.A(n_1618),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3302),
.Y(n_4205)
);

CKINVDCx5p33_ASAP7_75t_R g4206 ( 
.A(n_1033),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3278),
.Y(n_4207)
);

INVx1_ASAP7_75t_SL g4208 ( 
.A(n_1130),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_2024),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_226),
.Y(n_4210)
);

CKINVDCx20_ASAP7_75t_R g4211 ( 
.A(n_2467),
.Y(n_4211)
);

CKINVDCx5p33_ASAP7_75t_R g4212 ( 
.A(n_3227),
.Y(n_4212)
);

CKINVDCx5p33_ASAP7_75t_R g4213 ( 
.A(n_2461),
.Y(n_4213)
);

BUFx3_ASAP7_75t_L g4214 ( 
.A(n_2111),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_3318),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_2922),
.Y(n_4216)
);

CKINVDCx5p33_ASAP7_75t_R g4217 ( 
.A(n_3328),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_1708),
.Y(n_4218)
);

CKINVDCx5p33_ASAP7_75t_R g4219 ( 
.A(n_1006),
.Y(n_4219)
);

BUFx8_ASAP7_75t_SL g4220 ( 
.A(n_2895),
.Y(n_4220)
);

CKINVDCx5p33_ASAP7_75t_R g4221 ( 
.A(n_2414),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_3226),
.Y(n_4222)
);

CKINVDCx5p33_ASAP7_75t_R g4223 ( 
.A(n_3347),
.Y(n_4223)
);

CKINVDCx5p33_ASAP7_75t_R g4224 ( 
.A(n_1291),
.Y(n_4224)
);

CKINVDCx5p33_ASAP7_75t_R g4225 ( 
.A(n_3320),
.Y(n_4225)
);

CKINVDCx5p33_ASAP7_75t_R g4226 ( 
.A(n_680),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_2672),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_2547),
.Y(n_4228)
);

CKINVDCx5p33_ASAP7_75t_R g4229 ( 
.A(n_1244),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_34),
.Y(n_4230)
);

CKINVDCx5p33_ASAP7_75t_R g4231 ( 
.A(n_2942),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_2293),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_2917),
.Y(n_4233)
);

CKINVDCx20_ASAP7_75t_R g4234 ( 
.A(n_2430),
.Y(n_4234)
);

CKINVDCx20_ASAP7_75t_R g4235 ( 
.A(n_365),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_2167),
.Y(n_4236)
);

CKINVDCx5p33_ASAP7_75t_R g4237 ( 
.A(n_231),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_1894),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_1858),
.Y(n_4239)
);

CKINVDCx5p33_ASAP7_75t_R g4240 ( 
.A(n_2797),
.Y(n_4240)
);

BUFx3_ASAP7_75t_L g4241 ( 
.A(n_1395),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_882),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3288),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_2971),
.Y(n_4244)
);

CKINVDCx5p33_ASAP7_75t_R g4245 ( 
.A(n_3230),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_70),
.Y(n_4246)
);

CKINVDCx5p33_ASAP7_75t_R g4247 ( 
.A(n_1367),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_2126),
.Y(n_4248)
);

CKINVDCx5p33_ASAP7_75t_R g4249 ( 
.A(n_984),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_38),
.Y(n_4250)
);

HB1xp67_ASAP7_75t_L g4251 ( 
.A(n_3416),
.Y(n_4251)
);

BUFx6f_ASAP7_75t_L g4252 ( 
.A(n_3353),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_3380),
.Y(n_4253)
);

INVx1_ASAP7_75t_SL g4254 ( 
.A(n_3132),
.Y(n_4254)
);

BUFx6f_ASAP7_75t_L g4255 ( 
.A(n_2697),
.Y(n_4255)
);

BUFx8_ASAP7_75t_SL g4256 ( 
.A(n_457),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_870),
.Y(n_4257)
);

CKINVDCx20_ASAP7_75t_R g4258 ( 
.A(n_625),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_683),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_547),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_246),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_866),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_2761),
.Y(n_4263)
);

CKINVDCx5p33_ASAP7_75t_R g4264 ( 
.A(n_3362),
.Y(n_4264)
);

CKINVDCx5p33_ASAP7_75t_R g4265 ( 
.A(n_3418),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_2487),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_1816),
.Y(n_4267)
);

CKINVDCx20_ASAP7_75t_R g4268 ( 
.A(n_1430),
.Y(n_4268)
);

BUFx3_ASAP7_75t_L g4269 ( 
.A(n_3430),
.Y(n_4269)
);

CKINVDCx5p33_ASAP7_75t_R g4270 ( 
.A(n_3255),
.Y(n_4270)
);

CKINVDCx5p33_ASAP7_75t_R g4271 ( 
.A(n_2933),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_681),
.Y(n_4272)
);

CKINVDCx5p33_ASAP7_75t_R g4273 ( 
.A(n_2912),
.Y(n_4273)
);

CKINVDCx14_ASAP7_75t_R g4274 ( 
.A(n_2604),
.Y(n_4274)
);

HB1xp67_ASAP7_75t_L g4275 ( 
.A(n_581),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_1529),
.Y(n_4276)
);

CKINVDCx5p33_ASAP7_75t_R g4277 ( 
.A(n_3234),
.Y(n_4277)
);

CKINVDCx5p33_ASAP7_75t_R g4278 ( 
.A(n_273),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_2950),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_2236),
.Y(n_4280)
);

CKINVDCx5p33_ASAP7_75t_R g4281 ( 
.A(n_1285),
.Y(n_4281)
);

BUFx6f_ASAP7_75t_L g4282 ( 
.A(n_3319),
.Y(n_4282)
);

CKINVDCx5p33_ASAP7_75t_R g4283 ( 
.A(n_1805),
.Y(n_4283)
);

CKINVDCx5p33_ASAP7_75t_R g4284 ( 
.A(n_1368),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3323),
.Y(n_4285)
);

CKINVDCx5p33_ASAP7_75t_R g4286 ( 
.A(n_3032),
.Y(n_4286)
);

CKINVDCx5p33_ASAP7_75t_R g4287 ( 
.A(n_2944),
.Y(n_4287)
);

BUFx10_ASAP7_75t_L g4288 ( 
.A(n_953),
.Y(n_4288)
);

INVx1_ASAP7_75t_SL g4289 ( 
.A(n_168),
.Y(n_4289)
);

CKINVDCx5p33_ASAP7_75t_R g4290 ( 
.A(n_511),
.Y(n_4290)
);

CKINVDCx5p33_ASAP7_75t_R g4291 ( 
.A(n_3133),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_2906),
.Y(n_4292)
);

CKINVDCx5p33_ASAP7_75t_R g4293 ( 
.A(n_2371),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_1932),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_2691),
.Y(n_4295)
);

CKINVDCx5p33_ASAP7_75t_R g4296 ( 
.A(n_2041),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_3290),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_1505),
.Y(n_4298)
);

CKINVDCx5p33_ASAP7_75t_R g4299 ( 
.A(n_2048),
.Y(n_4299)
);

CKINVDCx5p33_ASAP7_75t_R g4300 ( 
.A(n_2826),
.Y(n_4300)
);

CKINVDCx5p33_ASAP7_75t_R g4301 ( 
.A(n_1409),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_2208),
.Y(n_4302)
);

CKINVDCx5p33_ASAP7_75t_R g4303 ( 
.A(n_3414),
.Y(n_4303)
);

BUFx6f_ASAP7_75t_L g4304 ( 
.A(n_1230),
.Y(n_4304)
);

CKINVDCx5p33_ASAP7_75t_R g4305 ( 
.A(n_451),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_3299),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_477),
.Y(n_4307)
);

CKINVDCx5p33_ASAP7_75t_R g4308 ( 
.A(n_1352),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_1209),
.Y(n_4309)
);

CKINVDCx5p33_ASAP7_75t_R g4310 ( 
.A(n_1064),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_3236),
.Y(n_4311)
);

CKINVDCx5p33_ASAP7_75t_R g4312 ( 
.A(n_2796),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_2893),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_457),
.Y(n_4314)
);

CKINVDCx5p33_ASAP7_75t_R g4315 ( 
.A(n_1077),
.Y(n_4315)
);

INVx2_ASAP7_75t_SL g4316 ( 
.A(n_1671),
.Y(n_4316)
);

CKINVDCx5p33_ASAP7_75t_R g4317 ( 
.A(n_3216),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3277),
.Y(n_4318)
);

CKINVDCx5p33_ASAP7_75t_R g4319 ( 
.A(n_2876),
.Y(n_4319)
);

CKINVDCx5p33_ASAP7_75t_R g4320 ( 
.A(n_1234),
.Y(n_4320)
);

CKINVDCx5p33_ASAP7_75t_R g4321 ( 
.A(n_1253),
.Y(n_4321)
);

CKINVDCx5p33_ASAP7_75t_R g4322 ( 
.A(n_2897),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_1072),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_1553),
.Y(n_4324)
);

CKINVDCx5p33_ASAP7_75t_R g4325 ( 
.A(n_2922),
.Y(n_4325)
);

CKINVDCx20_ASAP7_75t_R g4326 ( 
.A(n_2189),
.Y(n_4326)
);

CKINVDCx5p33_ASAP7_75t_R g4327 ( 
.A(n_2563),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_2258),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_2520),
.Y(n_4329)
);

BUFx8_ASAP7_75t_SL g4330 ( 
.A(n_2250),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_503),
.Y(n_4331)
);

CKINVDCx5p33_ASAP7_75t_R g4332 ( 
.A(n_1044),
.Y(n_4332)
);

BUFx10_ASAP7_75t_L g4333 ( 
.A(n_3266),
.Y(n_4333)
);

CKINVDCx5p33_ASAP7_75t_R g4334 ( 
.A(n_1894),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_953),
.Y(n_4335)
);

CKINVDCx5p33_ASAP7_75t_R g4336 ( 
.A(n_2315),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_2274),
.Y(n_4337)
);

CKINVDCx20_ASAP7_75t_R g4338 ( 
.A(n_612),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_2150),
.Y(n_4339)
);

CKINVDCx5p33_ASAP7_75t_R g4340 ( 
.A(n_1958),
.Y(n_4340)
);

BUFx5_ASAP7_75t_L g4341 ( 
.A(n_3126),
.Y(n_4341)
);

CKINVDCx5p33_ASAP7_75t_R g4342 ( 
.A(n_346),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_1953),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_2729),
.Y(n_4344)
);

CKINVDCx5p33_ASAP7_75t_R g4345 ( 
.A(n_380),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_224),
.Y(n_4346)
);

CKINVDCx5p33_ASAP7_75t_R g4347 ( 
.A(n_2309),
.Y(n_4347)
);

INVx1_ASAP7_75t_SL g4348 ( 
.A(n_1510),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_3309),
.Y(n_4349)
);

BUFx10_ASAP7_75t_L g4350 ( 
.A(n_682),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_2702),
.Y(n_4351)
);

CKINVDCx20_ASAP7_75t_R g4352 ( 
.A(n_935),
.Y(n_4352)
);

BUFx3_ASAP7_75t_L g4353 ( 
.A(n_36),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3400),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3054),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_2855),
.Y(n_4356)
);

CKINVDCx5p33_ASAP7_75t_R g4357 ( 
.A(n_3411),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_3072),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_479),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_2635),
.Y(n_4360)
);

CKINVDCx5p33_ASAP7_75t_R g4361 ( 
.A(n_2142),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_1720),
.Y(n_4362)
);

CKINVDCx5p33_ASAP7_75t_R g4363 ( 
.A(n_2328),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_1350),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_1549),
.Y(n_4365)
);

INVx1_ASAP7_75t_SL g4366 ( 
.A(n_1432),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_434),
.Y(n_4367)
);

CKINVDCx5p33_ASAP7_75t_R g4368 ( 
.A(n_3348),
.Y(n_4368)
);

CKINVDCx5p33_ASAP7_75t_R g4369 ( 
.A(n_2442),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_1215),
.Y(n_4370)
);

BUFx10_ASAP7_75t_L g4371 ( 
.A(n_713),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_1278),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_427),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_1995),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_1348),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_2999),
.Y(n_4376)
);

CKINVDCx5p33_ASAP7_75t_R g4377 ( 
.A(n_433),
.Y(n_4377)
);

INVxp67_ASAP7_75t_SL g4378 ( 
.A(n_1169),
.Y(n_4378)
);

CKINVDCx5p33_ASAP7_75t_R g4379 ( 
.A(n_1570),
.Y(n_4379)
);

BUFx2_ASAP7_75t_L g4380 ( 
.A(n_1109),
.Y(n_4380)
);

CKINVDCx5p33_ASAP7_75t_R g4381 ( 
.A(n_2657),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_2511),
.Y(n_4382)
);

CKINVDCx20_ASAP7_75t_R g4383 ( 
.A(n_1402),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_635),
.Y(n_4384)
);

BUFx2_ASAP7_75t_L g4385 ( 
.A(n_2250),
.Y(n_4385)
);

INVx3_ASAP7_75t_L g4386 ( 
.A(n_364),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_1891),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_3325),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_2185),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_733),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_3419),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_3350),
.Y(n_4392)
);

INVx1_ASAP7_75t_SL g4393 ( 
.A(n_1088),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_1600),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_448),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_1866),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_1279),
.Y(n_4397)
);

CKINVDCx5p33_ASAP7_75t_R g4398 ( 
.A(n_2389),
.Y(n_4398)
);

HB1xp67_ASAP7_75t_L g4399 ( 
.A(n_547),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_747),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_3352),
.Y(n_4401)
);

INVxp67_ASAP7_75t_L g4402 ( 
.A(n_1684),
.Y(n_4402)
);

CKINVDCx5p33_ASAP7_75t_R g4403 ( 
.A(n_2354),
.Y(n_4403)
);

CKINVDCx20_ASAP7_75t_R g4404 ( 
.A(n_1197),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_1832),
.Y(n_4405)
);

CKINVDCx20_ASAP7_75t_R g4406 ( 
.A(n_1921),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_763),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_1518),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_3357),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_3300),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_2125),
.Y(n_4411)
);

CKINVDCx20_ASAP7_75t_R g4412 ( 
.A(n_1163),
.Y(n_4412)
);

CKINVDCx16_ASAP7_75t_R g4413 ( 
.A(n_1421),
.Y(n_4413)
);

CKINVDCx5p33_ASAP7_75t_R g4414 ( 
.A(n_2147),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_3354),
.Y(n_4415)
);

INVx1_ASAP7_75t_SL g4416 ( 
.A(n_455),
.Y(n_4416)
);

INVx1_ASAP7_75t_SL g4417 ( 
.A(n_3322),
.Y(n_4417)
);

CKINVDCx20_ASAP7_75t_R g4418 ( 
.A(n_2807),
.Y(n_4418)
);

CKINVDCx5p33_ASAP7_75t_R g4419 ( 
.A(n_3405),
.Y(n_4419)
);

CKINVDCx5p33_ASAP7_75t_R g4420 ( 
.A(n_1727),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3240),
.Y(n_4421)
);

CKINVDCx5p33_ASAP7_75t_R g4422 ( 
.A(n_121),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_20),
.Y(n_4423)
);

CKINVDCx5p33_ASAP7_75t_R g4424 ( 
.A(n_2588),
.Y(n_4424)
);

INVx1_ASAP7_75t_SL g4425 ( 
.A(n_1352),
.Y(n_4425)
);

CKINVDCx5p33_ASAP7_75t_R g4426 ( 
.A(n_1095),
.Y(n_4426)
);

CKINVDCx5p33_ASAP7_75t_R g4427 ( 
.A(n_3313),
.Y(n_4427)
);

CKINVDCx5p33_ASAP7_75t_R g4428 ( 
.A(n_1573),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_2887),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_3398),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_1579),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3324),
.Y(n_4432)
);

INVx1_ASAP7_75t_SL g4433 ( 
.A(n_2640),
.Y(n_4433)
);

BUFx2_ASAP7_75t_L g4434 ( 
.A(n_3058),
.Y(n_4434)
);

CKINVDCx5p33_ASAP7_75t_R g4435 ( 
.A(n_3064),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_1208),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3386),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_3376),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_299),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_1358),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_1483),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_717),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_3252),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_939),
.Y(n_4444)
);

CKINVDCx5p33_ASAP7_75t_R g4445 ( 
.A(n_1644),
.Y(n_4445)
);

BUFx3_ASAP7_75t_L g4446 ( 
.A(n_2538),
.Y(n_4446)
);

BUFx2_ASAP7_75t_L g4447 ( 
.A(n_3360),
.Y(n_4447)
);

BUFx10_ASAP7_75t_L g4448 ( 
.A(n_595),
.Y(n_4448)
);

CKINVDCx16_ASAP7_75t_R g4449 ( 
.A(n_2085),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_2048),
.Y(n_4450)
);

CKINVDCx5p33_ASAP7_75t_R g4451 ( 
.A(n_136),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_3272),
.Y(n_4452)
);

CKINVDCx20_ASAP7_75t_R g4453 ( 
.A(n_3172),
.Y(n_4453)
);

CKINVDCx5p33_ASAP7_75t_R g4454 ( 
.A(n_3245),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_2881),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_1963),
.Y(n_4456)
);

INVx2_ASAP7_75t_SL g4457 ( 
.A(n_790),
.Y(n_4457)
);

BUFx10_ASAP7_75t_L g4458 ( 
.A(n_1903),
.Y(n_4458)
);

CKINVDCx5p33_ASAP7_75t_R g4459 ( 
.A(n_1454),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_1246),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_3338),
.Y(n_4461)
);

BUFx3_ASAP7_75t_L g4462 ( 
.A(n_1663),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_237),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_2166),
.Y(n_4464)
);

CKINVDCx20_ASAP7_75t_R g4465 ( 
.A(n_1085),
.Y(n_4465)
);

CKINVDCx5p33_ASAP7_75t_R g4466 ( 
.A(n_2633),
.Y(n_4466)
);

CKINVDCx5p33_ASAP7_75t_R g4467 ( 
.A(n_2916),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_67),
.Y(n_4468)
);

CKINVDCx5p33_ASAP7_75t_R g4469 ( 
.A(n_1693),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_2184),
.Y(n_4470)
);

BUFx8_ASAP7_75t_SL g4471 ( 
.A(n_126),
.Y(n_4471)
);

BUFx6f_ASAP7_75t_L g4472 ( 
.A(n_1086),
.Y(n_4472)
);

CKINVDCx5p33_ASAP7_75t_R g4473 ( 
.A(n_1311),
.Y(n_4473)
);

BUFx10_ASAP7_75t_L g4474 ( 
.A(n_88),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_2107),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_711),
.Y(n_4476)
);

CKINVDCx5p33_ASAP7_75t_R g4477 ( 
.A(n_1270),
.Y(n_4477)
);

CKINVDCx5p33_ASAP7_75t_R g4478 ( 
.A(n_2979),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_3359),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_1762),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_934),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_3084),
.Y(n_4482)
);

BUFx10_ASAP7_75t_L g4483 ( 
.A(n_176),
.Y(n_4483)
);

HB1xp67_ASAP7_75t_L g4484 ( 
.A(n_505),
.Y(n_4484)
);

CKINVDCx5p33_ASAP7_75t_R g4485 ( 
.A(n_332),
.Y(n_4485)
);

BUFx3_ASAP7_75t_L g4486 ( 
.A(n_3240),
.Y(n_4486)
);

CKINVDCx5p33_ASAP7_75t_R g4487 ( 
.A(n_1300),
.Y(n_4487)
);

CKINVDCx20_ASAP7_75t_R g4488 ( 
.A(n_1434),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_3301),
.Y(n_4489)
);

CKINVDCx5p33_ASAP7_75t_R g4490 ( 
.A(n_1667),
.Y(n_4490)
);

CKINVDCx20_ASAP7_75t_R g4491 ( 
.A(n_2808),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_469),
.Y(n_4492)
);

CKINVDCx5p33_ASAP7_75t_R g4493 ( 
.A(n_1575),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_983),
.Y(n_4494)
);

CKINVDCx5p33_ASAP7_75t_R g4495 ( 
.A(n_2223),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_118),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_2899),
.Y(n_4497)
);

BUFx3_ASAP7_75t_L g4498 ( 
.A(n_3361),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3253),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_2543),
.Y(n_4500)
);

INVx2_ASAP7_75t_L g4501 ( 
.A(n_676),
.Y(n_4501)
);

BUFx10_ASAP7_75t_L g4502 ( 
.A(n_2312),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_2553),
.Y(n_4503)
);

BUFx3_ASAP7_75t_L g4504 ( 
.A(n_3381),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_2358),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_2613),
.Y(n_4506)
);

INVx1_ASAP7_75t_SL g4507 ( 
.A(n_2131),
.Y(n_4507)
);

CKINVDCx5p33_ASAP7_75t_R g4508 ( 
.A(n_2918),
.Y(n_4508)
);

CKINVDCx14_ASAP7_75t_R g4509 ( 
.A(n_1671),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3342),
.Y(n_4510)
);

CKINVDCx5p33_ASAP7_75t_R g4511 ( 
.A(n_1262),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_3297),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_1353),
.Y(n_4513)
);

CKINVDCx5p33_ASAP7_75t_R g4514 ( 
.A(n_2479),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_1641),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_1494),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_1701),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_2013),
.Y(n_4518)
);

INVxp67_ASAP7_75t_L g4519 ( 
.A(n_3156),
.Y(n_4519)
);

CKINVDCx5p33_ASAP7_75t_R g4520 ( 
.A(n_1732),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3216),
.Y(n_4521)
);

CKINVDCx20_ASAP7_75t_R g4522 ( 
.A(n_3369),
.Y(n_4522)
);

BUFx3_ASAP7_75t_L g4523 ( 
.A(n_2762),
.Y(n_4523)
);

CKINVDCx5p33_ASAP7_75t_R g4524 ( 
.A(n_1369),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_802),
.Y(n_4525)
);

CKINVDCx5p33_ASAP7_75t_R g4526 ( 
.A(n_1515),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_3385),
.Y(n_4527)
);

CKINVDCx5p33_ASAP7_75t_R g4528 ( 
.A(n_2388),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_2668),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_1910),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_2004),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_1605),
.Y(n_4532)
);

CKINVDCx5p33_ASAP7_75t_R g4533 ( 
.A(n_1058),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_2918),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_2593),
.Y(n_4535)
);

CKINVDCx5p33_ASAP7_75t_R g4536 ( 
.A(n_1971),
.Y(n_4536)
);

CKINVDCx5p33_ASAP7_75t_R g4537 ( 
.A(n_1507),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_194),
.Y(n_4538)
);

CKINVDCx5p33_ASAP7_75t_R g4539 ( 
.A(n_1019),
.Y(n_4539)
);

CKINVDCx5p33_ASAP7_75t_R g4540 ( 
.A(n_2307),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_3275),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_1501),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_1931),
.Y(n_4543)
);

CKINVDCx5p33_ASAP7_75t_R g4544 ( 
.A(n_1540),
.Y(n_4544)
);

CKINVDCx5p33_ASAP7_75t_R g4545 ( 
.A(n_1185),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_3402),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_2771),
.Y(n_4547)
);

CKINVDCx5p33_ASAP7_75t_R g4548 ( 
.A(n_1770),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_714),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_2782),
.Y(n_4550)
);

CKINVDCx20_ASAP7_75t_R g4551 ( 
.A(n_706),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_2364),
.Y(n_4552)
);

CKINVDCx5p33_ASAP7_75t_R g4553 ( 
.A(n_1806),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_3436),
.Y(n_4554)
);

CKINVDCx5p33_ASAP7_75t_R g4555 ( 
.A(n_943),
.Y(n_4555)
);

BUFx3_ASAP7_75t_L g4556 ( 
.A(n_2940),
.Y(n_4556)
);

CKINVDCx5p33_ASAP7_75t_R g4557 ( 
.A(n_1091),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_523),
.Y(n_4558)
);

CKINVDCx20_ASAP7_75t_R g4559 ( 
.A(n_107),
.Y(n_4559)
);

CKINVDCx5p33_ASAP7_75t_R g4560 ( 
.A(n_2170),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3417),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_831),
.Y(n_4562)
);

BUFx3_ASAP7_75t_L g4563 ( 
.A(n_812),
.Y(n_4563)
);

CKINVDCx20_ASAP7_75t_R g4564 ( 
.A(n_3022),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_3028),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_1255),
.Y(n_4566)
);

BUFx3_ASAP7_75t_L g4567 ( 
.A(n_2986),
.Y(n_4567)
);

CKINVDCx5p33_ASAP7_75t_R g4568 ( 
.A(n_2727),
.Y(n_4568)
);

CKINVDCx5p33_ASAP7_75t_R g4569 ( 
.A(n_278),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_1693),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_3310),
.Y(n_4571)
);

CKINVDCx5p33_ASAP7_75t_R g4572 ( 
.A(n_2347),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_1410),
.Y(n_4573)
);

CKINVDCx5p33_ASAP7_75t_R g4574 ( 
.A(n_2551),
.Y(n_4574)
);

CKINVDCx5p33_ASAP7_75t_R g4575 ( 
.A(n_1599),
.Y(n_4575)
);

CKINVDCx5p33_ASAP7_75t_R g4576 ( 
.A(n_306),
.Y(n_4576)
);

CKINVDCx5p33_ASAP7_75t_R g4577 ( 
.A(n_956),
.Y(n_4577)
);

CKINVDCx5p33_ASAP7_75t_R g4578 ( 
.A(n_1725),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_3420),
.Y(n_4579)
);

CKINVDCx5p33_ASAP7_75t_R g4580 ( 
.A(n_2593),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_3332),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_599),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_3018),
.Y(n_4583)
);

CKINVDCx5p33_ASAP7_75t_R g4584 ( 
.A(n_563),
.Y(n_4584)
);

CKINVDCx5p33_ASAP7_75t_R g4585 ( 
.A(n_2956),
.Y(n_4585)
);

CKINVDCx5p33_ASAP7_75t_R g4586 ( 
.A(n_1327),
.Y(n_4586)
);

CKINVDCx5p33_ASAP7_75t_R g4587 ( 
.A(n_84),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_619),
.Y(n_4588)
);

BUFx3_ASAP7_75t_L g4589 ( 
.A(n_668),
.Y(n_4589)
);

INVx1_ASAP7_75t_SL g4590 ( 
.A(n_1296),
.Y(n_4590)
);

CKINVDCx20_ASAP7_75t_R g4591 ( 
.A(n_657),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_1723),
.Y(n_4592)
);

CKINVDCx5p33_ASAP7_75t_R g4593 ( 
.A(n_82),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_2921),
.Y(n_4594)
);

HB1xp67_ASAP7_75t_L g4595 ( 
.A(n_1445),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_752),
.Y(n_4596)
);

INVx1_ASAP7_75t_SL g4597 ( 
.A(n_3357),
.Y(n_4597)
);

BUFx3_ASAP7_75t_L g4598 ( 
.A(n_3303),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_1655),
.Y(n_4599)
);

CKINVDCx5p33_ASAP7_75t_R g4600 ( 
.A(n_3037),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_760),
.Y(n_4601)
);

CKINVDCx5p33_ASAP7_75t_R g4602 ( 
.A(n_1629),
.Y(n_4602)
);

INVx2_ASAP7_75t_SL g4603 ( 
.A(n_3088),
.Y(n_4603)
);

CKINVDCx20_ASAP7_75t_R g4604 ( 
.A(n_557),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_1554),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_3377),
.Y(n_4606)
);

CKINVDCx5p33_ASAP7_75t_R g4607 ( 
.A(n_1286),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_186),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_1354),
.Y(n_4609)
);

CKINVDCx5p33_ASAP7_75t_R g4610 ( 
.A(n_3242),
.Y(n_4610)
);

CKINVDCx5p33_ASAP7_75t_R g4611 ( 
.A(n_2353),
.Y(n_4611)
);

CKINVDCx5p33_ASAP7_75t_R g4612 ( 
.A(n_3333),
.Y(n_4612)
);

CKINVDCx20_ASAP7_75t_R g4613 ( 
.A(n_3387),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_2504),
.Y(n_4614)
);

CKINVDCx5p33_ASAP7_75t_R g4615 ( 
.A(n_488),
.Y(n_4615)
);

CKINVDCx5p33_ASAP7_75t_R g4616 ( 
.A(n_7),
.Y(n_4616)
);

CKINVDCx5p33_ASAP7_75t_R g4617 ( 
.A(n_1832),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_2742),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_561),
.Y(n_4619)
);

BUFx10_ASAP7_75t_L g4620 ( 
.A(n_2346),
.Y(n_4620)
);

BUFx6f_ASAP7_75t_L g4621 ( 
.A(n_1661),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_2720),
.Y(n_4622)
);

CKINVDCx5p33_ASAP7_75t_R g4623 ( 
.A(n_3359),
.Y(n_4623)
);

CKINVDCx5p33_ASAP7_75t_R g4624 ( 
.A(n_1350),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_300),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_3401),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_3091),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_2932),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_2966),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_1765),
.Y(n_4630)
);

CKINVDCx5p33_ASAP7_75t_R g4631 ( 
.A(n_1027),
.Y(n_4631)
);

CKINVDCx5p33_ASAP7_75t_R g4632 ( 
.A(n_1481),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_1389),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_3366),
.Y(n_4634)
);

CKINVDCx5p33_ASAP7_75t_R g4635 ( 
.A(n_3194),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_2287),
.Y(n_4636)
);

BUFx5_ASAP7_75t_L g4637 ( 
.A(n_2894),
.Y(n_4637)
);

CKINVDCx20_ASAP7_75t_R g4638 ( 
.A(n_1854),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_489),
.Y(n_4639)
);

CKINVDCx20_ASAP7_75t_R g4640 ( 
.A(n_483),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_2597),
.Y(n_4641)
);

CKINVDCx16_ASAP7_75t_R g4642 ( 
.A(n_2034),
.Y(n_4642)
);

CKINVDCx5p33_ASAP7_75t_R g4643 ( 
.A(n_2699),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_1987),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_472),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_1858),
.Y(n_4646)
);

INVx2_ASAP7_75t_L g4647 ( 
.A(n_577),
.Y(n_4647)
);

CKINVDCx5p33_ASAP7_75t_R g4648 ( 
.A(n_2236),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_2423),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_3457),
.Y(n_4650)
);

BUFx6f_ASAP7_75t_L g4651 ( 
.A(n_2318),
.Y(n_4651)
);

CKINVDCx5p33_ASAP7_75t_R g4652 ( 
.A(n_1735),
.Y(n_4652)
);

BUFx3_ASAP7_75t_L g4653 ( 
.A(n_1306),
.Y(n_4653)
);

BUFx2_ASAP7_75t_SL g4654 ( 
.A(n_2780),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_3232),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_326),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_2578),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_2017),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_553),
.Y(n_4659)
);

CKINVDCx5p33_ASAP7_75t_R g4660 ( 
.A(n_3412),
.Y(n_4660)
);

BUFx10_ASAP7_75t_L g4661 ( 
.A(n_1310),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_1283),
.Y(n_4662)
);

CKINVDCx5p33_ASAP7_75t_R g4663 ( 
.A(n_865),
.Y(n_4663)
);

CKINVDCx5p33_ASAP7_75t_R g4664 ( 
.A(n_3362),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_975),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_3091),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_3343),
.Y(n_4667)
);

CKINVDCx20_ASAP7_75t_R g4668 ( 
.A(n_1055),
.Y(n_4668)
);

CKINVDCx5p33_ASAP7_75t_R g4669 ( 
.A(n_1182),
.Y(n_4669)
);

CKINVDCx5p33_ASAP7_75t_R g4670 ( 
.A(n_2177),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_3280),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_2650),
.Y(n_4672)
);

CKINVDCx20_ASAP7_75t_R g4673 ( 
.A(n_3394),
.Y(n_4673)
);

CKINVDCx20_ASAP7_75t_R g4674 ( 
.A(n_1853),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_3445),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_995),
.Y(n_4676)
);

CKINVDCx5p33_ASAP7_75t_R g4677 ( 
.A(n_1429),
.Y(n_4677)
);

BUFx10_ASAP7_75t_L g4678 ( 
.A(n_2011),
.Y(n_4678)
);

BUFx3_ASAP7_75t_L g4679 ( 
.A(n_1554),
.Y(n_4679)
);

CKINVDCx5p33_ASAP7_75t_R g4680 ( 
.A(n_3433),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_1437),
.Y(n_4681)
);

CKINVDCx16_ASAP7_75t_R g4682 ( 
.A(n_997),
.Y(n_4682)
);

BUFx5_ASAP7_75t_L g4683 ( 
.A(n_3384),
.Y(n_4683)
);

CKINVDCx20_ASAP7_75t_R g4684 ( 
.A(n_2997),
.Y(n_4684)
);

CKINVDCx5p33_ASAP7_75t_R g4685 ( 
.A(n_1037),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_1910),
.Y(n_4686)
);

CKINVDCx5p33_ASAP7_75t_R g4687 ( 
.A(n_3358),
.Y(n_4687)
);

CKINVDCx5p33_ASAP7_75t_R g4688 ( 
.A(n_3238),
.Y(n_4688)
);

CKINVDCx5p33_ASAP7_75t_R g4689 ( 
.A(n_1464),
.Y(n_4689)
);

BUFx10_ASAP7_75t_L g4690 ( 
.A(n_2900),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_1842),
.Y(n_4691)
);

BUFx6f_ASAP7_75t_L g4692 ( 
.A(n_842),
.Y(n_4692)
);

CKINVDCx20_ASAP7_75t_R g4693 ( 
.A(n_1566),
.Y(n_4693)
);

CKINVDCx5p33_ASAP7_75t_R g4694 ( 
.A(n_2987),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_846),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_642),
.Y(n_4696)
);

INVx1_ASAP7_75t_SL g4697 ( 
.A(n_1464),
.Y(n_4697)
);

CKINVDCx5p33_ASAP7_75t_R g4698 ( 
.A(n_259),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_3337),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_228),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_1799),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_1844),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_3311),
.Y(n_4703)
);

CKINVDCx5p33_ASAP7_75t_R g4704 ( 
.A(n_2225),
.Y(n_4704)
);

CKINVDCx5p33_ASAP7_75t_R g4705 ( 
.A(n_2848),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_1908),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_2121),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_2612),
.Y(n_4708)
);

CKINVDCx5p33_ASAP7_75t_R g4709 ( 
.A(n_1458),
.Y(n_4709)
);

CKINVDCx20_ASAP7_75t_R g4710 ( 
.A(n_3375),
.Y(n_4710)
);

CKINVDCx5p33_ASAP7_75t_R g4711 ( 
.A(n_824),
.Y(n_4711)
);

BUFx6f_ASAP7_75t_L g4712 ( 
.A(n_940),
.Y(n_4712)
);

CKINVDCx20_ASAP7_75t_R g4713 ( 
.A(n_2514),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_16),
.Y(n_4714)
);

BUFx3_ASAP7_75t_L g4715 ( 
.A(n_568),
.Y(n_4715)
);

CKINVDCx5p33_ASAP7_75t_R g4716 ( 
.A(n_314),
.Y(n_4716)
);

CKINVDCx5p33_ASAP7_75t_R g4717 ( 
.A(n_3254),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_737),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_2164),
.Y(n_4719)
);

CKINVDCx16_ASAP7_75t_R g4720 ( 
.A(n_603),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_3212),
.Y(n_4721)
);

CKINVDCx5p33_ASAP7_75t_R g4722 ( 
.A(n_2704),
.Y(n_4722)
);

CKINVDCx5p33_ASAP7_75t_R g4723 ( 
.A(n_2680),
.Y(n_4723)
);

CKINVDCx5p33_ASAP7_75t_R g4724 ( 
.A(n_3222),
.Y(n_4724)
);

CKINVDCx16_ASAP7_75t_R g4725 ( 
.A(n_2327),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_960),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_270),
.Y(n_4727)
);

CKINVDCx5p33_ASAP7_75t_R g4728 ( 
.A(n_3269),
.Y(n_4728)
);

CKINVDCx5p33_ASAP7_75t_R g4729 ( 
.A(n_2733),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_624),
.Y(n_4730)
);

CKINVDCx5p33_ASAP7_75t_R g4731 ( 
.A(n_3408),
.Y(n_4731)
);

BUFx3_ASAP7_75t_L g4732 ( 
.A(n_869),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_326),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_573),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_3140),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_15),
.Y(n_4736)
);

BUFx6f_ASAP7_75t_L g4737 ( 
.A(n_3287),
.Y(n_4737)
);

CKINVDCx20_ASAP7_75t_R g4738 ( 
.A(n_3291),
.Y(n_4738)
);

BUFx3_ASAP7_75t_L g4739 ( 
.A(n_3307),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_2707),
.Y(n_4740)
);

CKINVDCx5p33_ASAP7_75t_R g4741 ( 
.A(n_2755),
.Y(n_4741)
);

CKINVDCx5p33_ASAP7_75t_R g4742 ( 
.A(n_1846),
.Y(n_4742)
);

CKINVDCx5p33_ASAP7_75t_R g4743 ( 
.A(n_3465),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_3286),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_3036),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_2517),
.Y(n_4746)
);

CKINVDCx5p33_ASAP7_75t_R g4747 ( 
.A(n_1768),
.Y(n_4747)
);

CKINVDCx5p33_ASAP7_75t_R g4748 ( 
.A(n_1143),
.Y(n_4748)
);

INVx1_ASAP7_75t_SL g4749 ( 
.A(n_3372),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_1242),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_2304),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_1421),
.Y(n_4752)
);

CKINVDCx5p33_ASAP7_75t_R g4753 ( 
.A(n_1237),
.Y(n_4753)
);

CKINVDCx5p33_ASAP7_75t_R g4754 ( 
.A(n_1240),
.Y(n_4754)
);

CKINVDCx5p33_ASAP7_75t_R g4755 ( 
.A(n_3335),
.Y(n_4755)
);

CKINVDCx5p33_ASAP7_75t_R g4756 ( 
.A(n_3304),
.Y(n_4756)
);

CKINVDCx5p33_ASAP7_75t_R g4757 ( 
.A(n_1623),
.Y(n_4757)
);

CKINVDCx5p33_ASAP7_75t_R g4758 ( 
.A(n_2728),
.Y(n_4758)
);

CKINVDCx5p33_ASAP7_75t_R g4759 ( 
.A(n_1559),
.Y(n_4759)
);

BUFx2_ASAP7_75t_L g4760 ( 
.A(n_2809),
.Y(n_4760)
);

CKINVDCx20_ASAP7_75t_R g4761 ( 
.A(n_3245),
.Y(n_4761)
);

CKINVDCx5p33_ASAP7_75t_R g4762 ( 
.A(n_3289),
.Y(n_4762)
);

CKINVDCx5p33_ASAP7_75t_R g4763 ( 
.A(n_2688),
.Y(n_4763)
);

CKINVDCx5p33_ASAP7_75t_R g4764 ( 
.A(n_3421),
.Y(n_4764)
);

BUFx6f_ASAP7_75t_L g4765 ( 
.A(n_3396),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_1344),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_87),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_3126),
.Y(n_4768)
);

CKINVDCx5p33_ASAP7_75t_R g4769 ( 
.A(n_3247),
.Y(n_4769)
);

CKINVDCx5p33_ASAP7_75t_R g4770 ( 
.A(n_2130),
.Y(n_4770)
);

HB1xp67_ASAP7_75t_L g4771 ( 
.A(n_1398),
.Y(n_4771)
);

CKINVDCx16_ASAP7_75t_R g4772 ( 
.A(n_1507),
.Y(n_4772)
);

BUFx8_ASAP7_75t_SL g4773 ( 
.A(n_1857),
.Y(n_4773)
);

INVx2_ASAP7_75t_SL g4774 ( 
.A(n_2612),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_251),
.Y(n_4775)
);

BUFx3_ASAP7_75t_L g4776 ( 
.A(n_1934),
.Y(n_4776)
);

CKINVDCx5p33_ASAP7_75t_R g4777 ( 
.A(n_2603),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_1882),
.Y(n_4778)
);

BUFx2_ASAP7_75t_SL g4779 ( 
.A(n_2749),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_2049),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_1044),
.Y(n_4781)
);

INVx1_ASAP7_75t_SL g4782 ( 
.A(n_141),
.Y(n_4782)
);

CKINVDCx20_ASAP7_75t_R g4783 ( 
.A(n_1612),
.Y(n_4783)
);

INVx1_ASAP7_75t_SL g4784 ( 
.A(n_2311),
.Y(n_4784)
);

CKINVDCx14_ASAP7_75t_R g4785 ( 
.A(n_3183),
.Y(n_4785)
);

INVx1_ASAP7_75t_SL g4786 ( 
.A(n_2278),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_3372),
.Y(n_4787)
);

CKINVDCx5p33_ASAP7_75t_R g4788 ( 
.A(n_3246),
.Y(n_4788)
);

INVx1_ASAP7_75t_SL g4789 ( 
.A(n_3230),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_2280),
.Y(n_4790)
);

BUFx10_ASAP7_75t_L g4791 ( 
.A(n_49),
.Y(n_4791)
);

CKINVDCx20_ASAP7_75t_R g4792 ( 
.A(n_899),
.Y(n_4792)
);

CKINVDCx20_ASAP7_75t_R g4793 ( 
.A(n_3228),
.Y(n_4793)
);

BUFx2_ASAP7_75t_L g4794 ( 
.A(n_882),
.Y(n_4794)
);

CKINVDCx20_ASAP7_75t_R g4795 ( 
.A(n_781),
.Y(n_4795)
);

INVx1_ASAP7_75t_SL g4796 ( 
.A(n_2965),
.Y(n_4796)
);

CKINVDCx16_ASAP7_75t_R g4797 ( 
.A(n_1262),
.Y(n_4797)
);

INVx1_ASAP7_75t_SL g4798 ( 
.A(n_131),
.Y(n_4798)
);

CKINVDCx20_ASAP7_75t_R g4799 ( 
.A(n_141),
.Y(n_4799)
);

CKINVDCx5p33_ASAP7_75t_R g4800 ( 
.A(n_2657),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_3391),
.Y(n_4801)
);

CKINVDCx5p33_ASAP7_75t_R g4802 ( 
.A(n_2346),
.Y(n_4802)
);

CKINVDCx20_ASAP7_75t_R g4803 ( 
.A(n_1422),
.Y(n_4803)
);

CKINVDCx5p33_ASAP7_75t_R g4804 ( 
.A(n_2815),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_2205),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_219),
.Y(n_4806)
);

BUFx6f_ASAP7_75t_L g4807 ( 
.A(n_3367),
.Y(n_4807)
);

BUFx3_ASAP7_75t_L g4808 ( 
.A(n_2201),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_2311),
.Y(n_4809)
);

INVx2_ASAP7_75t_L g4810 ( 
.A(n_3167),
.Y(n_4810)
);

CKINVDCx5p33_ASAP7_75t_R g4811 ( 
.A(n_3224),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_3295),
.Y(n_4812)
);

BUFx6f_ASAP7_75t_L g4813 ( 
.A(n_24),
.Y(n_4813)
);

CKINVDCx5p33_ASAP7_75t_R g4814 ( 
.A(n_2360),
.Y(n_4814)
);

CKINVDCx5p33_ASAP7_75t_R g4815 ( 
.A(n_3273),
.Y(n_4815)
);

CKINVDCx20_ASAP7_75t_R g4816 ( 
.A(n_2061),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_1923),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_688),
.Y(n_4818)
);

CKINVDCx20_ASAP7_75t_R g4819 ( 
.A(n_902),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_1975),
.Y(n_4820)
);

CKINVDCx16_ASAP7_75t_R g4821 ( 
.A(n_2274),
.Y(n_4821)
);

INVx2_ASAP7_75t_SL g4822 ( 
.A(n_473),
.Y(n_4822)
);

CKINVDCx20_ASAP7_75t_R g4823 ( 
.A(n_696),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_7),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_2504),
.Y(n_4825)
);

BUFx10_ASAP7_75t_L g4826 ( 
.A(n_3297),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_525),
.Y(n_4827)
);

CKINVDCx5p33_ASAP7_75t_R g4828 ( 
.A(n_3223),
.Y(n_4828)
);

BUFx6f_ASAP7_75t_L g4829 ( 
.A(n_2232),
.Y(n_4829)
);

CKINVDCx5p33_ASAP7_75t_R g4830 ( 
.A(n_3407),
.Y(n_4830)
);

INVx1_ASAP7_75t_SL g4831 ( 
.A(n_2764),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_1925),
.Y(n_4832)
);

CKINVDCx20_ASAP7_75t_R g4833 ( 
.A(n_3261),
.Y(n_4833)
);

CKINVDCx5p33_ASAP7_75t_R g4834 ( 
.A(n_595),
.Y(n_4834)
);

CKINVDCx5p33_ASAP7_75t_R g4835 ( 
.A(n_2517),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_485),
.Y(n_4836)
);

CKINVDCx5p33_ASAP7_75t_R g4837 ( 
.A(n_3085),
.Y(n_4837)
);

CKINVDCx5p33_ASAP7_75t_R g4838 ( 
.A(n_3417),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_511),
.Y(n_4839)
);

CKINVDCx20_ASAP7_75t_R g4840 ( 
.A(n_3119),
.Y(n_4840)
);

CKINVDCx5p33_ASAP7_75t_R g4841 ( 
.A(n_1585),
.Y(n_4841)
);

CKINVDCx5p33_ASAP7_75t_R g4842 ( 
.A(n_3194),
.Y(n_4842)
);

CKINVDCx5p33_ASAP7_75t_R g4843 ( 
.A(n_837),
.Y(n_4843)
);

CKINVDCx5p33_ASAP7_75t_R g4844 ( 
.A(n_2307),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_1485),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_1110),
.Y(n_4846)
);

CKINVDCx5p33_ASAP7_75t_R g4847 ( 
.A(n_2729),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_1256),
.Y(n_4848)
);

CKINVDCx16_ASAP7_75t_R g4849 ( 
.A(n_1187),
.Y(n_4849)
);

BUFx10_ASAP7_75t_L g4850 ( 
.A(n_2081),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_802),
.Y(n_4851)
);

CKINVDCx5p33_ASAP7_75t_R g4852 ( 
.A(n_1366),
.Y(n_4852)
);

CKINVDCx5p33_ASAP7_75t_R g4853 ( 
.A(n_1919),
.Y(n_4853)
);

CKINVDCx20_ASAP7_75t_R g4854 ( 
.A(n_1310),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_2551),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_2384),
.Y(n_4856)
);

INVx1_ASAP7_75t_SL g4857 ( 
.A(n_2198),
.Y(n_4857)
);

CKINVDCx5p33_ASAP7_75t_R g4858 ( 
.A(n_2413),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_1400),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_1637),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_2818),
.Y(n_4861)
);

BUFx3_ASAP7_75t_L g4862 ( 
.A(n_2072),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_3232),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_3062),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_864),
.Y(n_4865)
);

CKINVDCx5p33_ASAP7_75t_R g4866 ( 
.A(n_2705),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_1564),
.Y(n_4867)
);

CKINVDCx5p33_ASAP7_75t_R g4868 ( 
.A(n_3424),
.Y(n_4868)
);

CKINVDCx5p33_ASAP7_75t_R g4869 ( 
.A(n_2579),
.Y(n_4869)
);

CKINVDCx5p33_ASAP7_75t_R g4870 ( 
.A(n_1167),
.Y(n_4870)
);

CKINVDCx20_ASAP7_75t_R g4871 ( 
.A(n_1266),
.Y(n_4871)
);

CKINVDCx5p33_ASAP7_75t_R g4872 ( 
.A(n_2505),
.Y(n_4872)
);

BUFx3_ASAP7_75t_L g4873 ( 
.A(n_3804),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_4256),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_3713),
.B(n_0),
.Y(n_4875)
);

INVx1_ASAP7_75t_SL g4876 ( 
.A(n_4471),
.Y(n_4876)
);

CKINVDCx5p33_ASAP7_75t_R g4877 ( 
.A(n_3794),
.Y(n_4877)
);

CKINVDCx20_ASAP7_75t_R g4878 ( 
.A(n_3776),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_3571),
.Y(n_4879)
);

BUFx3_ASAP7_75t_L g4880 ( 
.A(n_3999),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_3571),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_3571),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_4028),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_4220),
.Y(n_4884)
);

CKINVDCx16_ASAP7_75t_R g4885 ( 
.A(n_4124),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_3571),
.Y(n_4886)
);

BUFx6f_ASAP7_75t_L g4887 ( 
.A(n_3847),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_3571),
.Y(n_4888)
);

CKINVDCx5p33_ASAP7_75t_R g4889 ( 
.A(n_4330),
.Y(n_4889)
);

CKINVDCx14_ASAP7_75t_R g4890 ( 
.A(n_3953),
.Y(n_4890)
);

CKINVDCx5p33_ASAP7_75t_R g4891 ( 
.A(n_4773),
.Y(n_4891)
);

INVx2_ASAP7_75t_L g4892 ( 
.A(n_3762),
.Y(n_4892)
);

INVx1_ASAP7_75t_SL g4893 ( 
.A(n_3701),
.Y(n_4893)
);

BUFx10_ASAP7_75t_L g4894 ( 
.A(n_4275),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_3762),
.Y(n_4895)
);

CKINVDCx5p33_ASAP7_75t_R g4896 ( 
.A(n_4720),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_3762),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_3762),
.Y(n_4898)
);

INVxp67_ASAP7_75t_L g4899 ( 
.A(n_3873),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_3762),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4102),
.Y(n_4901)
);

CKINVDCx5p33_ASAP7_75t_R g4902 ( 
.A(n_4012),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4102),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4102),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4102),
.Y(n_4905)
);

CKINVDCx5p33_ASAP7_75t_R g4906 ( 
.A(n_4274),
.Y(n_4906)
);

CKINVDCx5p33_ASAP7_75t_R g4907 ( 
.A(n_4509),
.Y(n_4907)
);

CKINVDCx5p33_ASAP7_75t_R g4908 ( 
.A(n_4785),
.Y(n_4908)
);

NOR2xp67_ASAP7_75t_L g4909 ( 
.A(n_3825),
.B(n_0),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4102),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4341),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4341),
.Y(n_4912)
);

CKINVDCx16_ASAP7_75t_R g4913 ( 
.A(n_3574),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4341),
.Y(n_4914)
);

CKINVDCx5p33_ASAP7_75t_R g4915 ( 
.A(n_3696),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_3736),
.Y(n_4916)
);

CKINVDCx16_ASAP7_75t_R g4917 ( 
.A(n_3914),
.Y(n_4917)
);

CKINVDCx5p33_ASAP7_75t_R g4918 ( 
.A(n_4108),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4341),
.Y(n_4919)
);

CKINVDCx5p33_ASAP7_75t_R g4920 ( 
.A(n_4110),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_4127),
.Y(n_4921)
);

BUFx10_ASAP7_75t_L g4922 ( 
.A(n_4399),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_4413),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4341),
.Y(n_4924)
);

CKINVDCx5p33_ASAP7_75t_R g4925 ( 
.A(n_4449),
.Y(n_4925)
);

CKINVDCx20_ASAP7_75t_R g4926 ( 
.A(n_4642),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4637),
.Y(n_4927)
);

HB1xp67_ASAP7_75t_L g4928 ( 
.A(n_4484),
.Y(n_4928)
);

CKINVDCx5p33_ASAP7_75t_R g4929 ( 
.A(n_4682),
.Y(n_4929)
);

INVx2_ASAP7_75t_SL g4930 ( 
.A(n_3524),
.Y(n_4930)
);

CKINVDCx20_ASAP7_75t_R g4931 ( 
.A(n_4725),
.Y(n_4931)
);

CKINVDCx5p33_ASAP7_75t_R g4932 ( 
.A(n_4772),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4637),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4637),
.Y(n_4934)
);

CKINVDCx16_ASAP7_75t_R g4935 ( 
.A(n_4797),
.Y(n_4935)
);

HB1xp67_ASAP7_75t_L g4936 ( 
.A(n_4582),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4637),
.Y(n_4937)
);

CKINVDCx16_ASAP7_75t_R g4938 ( 
.A(n_4821),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4637),
.Y(n_4939)
);

INVx1_ASAP7_75t_SL g4940 ( 
.A(n_3542),
.Y(n_4940)
);

INVxp67_ASAP7_75t_SL g4941 ( 
.A(n_3951),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4683),
.Y(n_4942)
);

OR2x2_ASAP7_75t_L g4943 ( 
.A(n_4416),
.B(n_0),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4683),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4683),
.Y(n_4945)
);

BUFx6f_ASAP7_75t_L g4946 ( 
.A(n_3847),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4683),
.Y(n_4947)
);

CKINVDCx16_ASAP7_75t_R g4948 ( 
.A(n_4849),
.Y(n_4948)
);

BUFx6f_ASAP7_75t_L g4949 ( 
.A(n_3847),
.Y(n_4949)
);

INVx3_ASAP7_75t_L g4950 ( 
.A(n_3492),
.Y(n_4950)
);

CKINVDCx16_ASAP7_75t_R g4951 ( 
.A(n_3524),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_3483),
.Y(n_4952)
);

CKINVDCx5p33_ASAP7_75t_R g4953 ( 
.A(n_3486),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4683),
.Y(n_4954)
);

CKINVDCx20_ASAP7_75t_R g4955 ( 
.A(n_3490),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_3951),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_3487),
.Y(n_4957)
);

BUFx3_ASAP7_75t_L g4958 ( 
.A(n_4353),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4386),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4386),
.Y(n_4960)
);

NOR2xp67_ASAP7_75t_L g4961 ( 
.A(n_3825),
.B(n_1),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_3502),
.Y(n_4962)
);

INVx3_ASAP7_75t_L g4963 ( 
.A(n_3492),
.Y(n_4963)
);

CKINVDCx16_ASAP7_75t_R g4964 ( 
.A(n_3567),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_3515),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_3538),
.Y(n_4966)
);

NOR2xp67_ASAP7_75t_L g4967 ( 
.A(n_4402),
.B(n_1),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_3613),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_3641),
.Y(n_4969)
);

INVx1_ASAP7_75t_SL g4970 ( 
.A(n_3666),
.Y(n_4970)
);

BUFx3_ASAP7_75t_L g4971 ( 
.A(n_4563),
.Y(n_4971)
);

CKINVDCx16_ASAP7_75t_R g4972 ( 
.A(n_3567),
.Y(n_4972)
);

CKINVDCx5p33_ASAP7_75t_R g4973 ( 
.A(n_3493),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4865),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_3648),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_3651),
.Y(n_4976)
);

CKINVDCx5p33_ASAP7_75t_R g4977 ( 
.A(n_3497),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_3504),
.Y(n_4978)
);

BUFx6f_ASAP7_75t_L g4979 ( 
.A(n_4013),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_3702),
.Y(n_4980)
);

NOR2xp67_ASAP7_75t_L g4981 ( 
.A(n_4519),
.B(n_1),
.Y(n_4981)
);

CKINVDCx5p33_ASAP7_75t_R g4982 ( 
.A(n_3507),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_3790),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_3793),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_3816),
.Y(n_4985)
);

INVx2_ASAP7_75t_SL g4986 ( 
.A(n_3729),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_3834),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_3850),
.Y(n_4988)
);

CKINVDCx5p33_ASAP7_75t_R g4989 ( 
.A(n_3512),
.Y(n_4989)
);

CKINVDCx5p33_ASAP7_75t_R g4990 ( 
.A(n_3530),
.Y(n_4990)
);

BUFx3_ASAP7_75t_L g4991 ( 
.A(n_4589),
.Y(n_4991)
);

CKINVDCx5p33_ASAP7_75t_R g4992 ( 
.A(n_3539),
.Y(n_4992)
);

CKINVDCx5p33_ASAP7_75t_R g4993 ( 
.A(n_3540),
.Y(n_4993)
);

CKINVDCx5p33_ASAP7_75t_R g4994 ( 
.A(n_3549),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_3882),
.Y(n_4995)
);

CKINVDCx5p33_ASAP7_75t_R g4996 ( 
.A(n_3555),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_3885),
.Y(n_4997)
);

CKINVDCx20_ASAP7_75t_R g4998 ( 
.A(n_3553),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_3938),
.Y(n_4999)
);

CKINVDCx5p33_ASAP7_75t_R g5000 ( 
.A(n_3561),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_3947),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_3966),
.Y(n_5002)
);

INVx2_ASAP7_75t_SL g5003 ( 
.A(n_3729),
.Y(n_5003)
);

BUFx2_ASAP7_75t_L g5004 ( 
.A(n_3674),
.Y(n_5004)
);

CKINVDCx20_ASAP7_75t_R g5005 ( 
.A(n_3591),
.Y(n_5005)
);

BUFx6f_ASAP7_75t_L g5006 ( 
.A(n_4013),
.Y(n_5006)
);

BUFx2_ASAP7_75t_L g5007 ( 
.A(n_4202),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_3990),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_3995),
.Y(n_5009)
);

CKINVDCx20_ASAP7_75t_R g5010 ( 
.A(n_3604),
.Y(n_5010)
);

CKINVDCx20_ASAP7_75t_R g5011 ( 
.A(n_3617),
.Y(n_5011)
);

CKINVDCx20_ASAP7_75t_R g5012 ( 
.A(n_3631),
.Y(n_5012)
);

NOR2xp67_ASAP7_75t_L g5013 ( 
.A(n_3671),
.B(n_2),
.Y(n_5013)
);

CKINVDCx5p33_ASAP7_75t_R g5014 ( 
.A(n_3563),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4002),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4045),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4060),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4099),
.Y(n_5018)
);

CKINVDCx20_ASAP7_75t_R g5019 ( 
.A(n_3639),
.Y(n_5019)
);

CKINVDCx5p33_ASAP7_75t_R g5020 ( 
.A(n_3573),
.Y(n_5020)
);

CKINVDCx5p33_ASAP7_75t_R g5021 ( 
.A(n_3580),
.Y(n_5021)
);

CKINVDCx20_ASAP7_75t_R g5022 ( 
.A(n_3655),
.Y(n_5022)
);

CKINVDCx20_ASAP7_75t_R g5023 ( 
.A(n_3656),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4105),
.Y(n_5024)
);

BUFx3_ASAP7_75t_L g5025 ( 
.A(n_4715),
.Y(n_5025)
);

CKINVDCx5p33_ASAP7_75t_R g5026 ( 
.A(n_3583),
.Y(n_5026)
);

CKINVDCx20_ASAP7_75t_R g5027 ( 
.A(n_3710),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4115),
.Y(n_5028)
);

BUFx2_ASAP7_75t_L g5029 ( 
.A(n_4380),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_3594),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4137),
.Y(n_5031)
);

CKINVDCx5p33_ASAP7_75t_R g5032 ( 
.A(n_3600),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4153),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4174),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4210),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_3607),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4257),
.Y(n_5037)
);

OR2x2_ASAP7_75t_L g5038 ( 
.A(n_4782),
.B(n_2),
.Y(n_5038)
);

INVxp33_ASAP7_75t_SL g5039 ( 
.A(n_3719),
.Y(n_5039)
);

BUFx6f_ASAP7_75t_L g5040 ( 
.A(n_4013),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4260),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_4262),
.Y(n_5042)
);

BUFx3_ASAP7_75t_L g5043 ( 
.A(n_4732),
.Y(n_5043)
);

INVx2_ASAP7_75t_L g5044 ( 
.A(n_4272),
.Y(n_5044)
);

CKINVDCx5p33_ASAP7_75t_R g5045 ( 
.A(n_3608),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4307),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4314),
.Y(n_5047)
);

BUFx3_ASAP7_75t_L g5048 ( 
.A(n_3597),
.Y(n_5048)
);

NOR2xp67_ASAP7_75t_L g5049 ( 
.A(n_3805),
.B(n_2),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_3621),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4346),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4359),
.Y(n_5052)
);

CKINVDCx5p33_ASAP7_75t_R g5053 ( 
.A(n_3630),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4367),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_3632),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4384),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4395),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4400),
.Y(n_5058)
);

CKINVDCx20_ASAP7_75t_R g5059 ( 
.A(n_3745),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_3638),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4407),
.Y(n_5061)
);

CKINVDCx5p33_ASAP7_75t_R g5062 ( 
.A(n_3646),
.Y(n_5062)
);

BUFx10_ASAP7_75t_L g5063 ( 
.A(n_3654),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_3659),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4423),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4439),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4468),
.Y(n_5067)
);

BUFx3_ASAP7_75t_L g5068 ( 
.A(n_3612),
.Y(n_5068)
);

CKINVDCx20_ASAP7_75t_R g5069 ( 
.A(n_3747),
.Y(n_5069)
);

INVx1_ASAP7_75t_SL g5070 ( 
.A(n_4385),
.Y(n_5070)
);

BUFx6f_ASAP7_75t_L g5071 ( 
.A(n_4138),
.Y(n_5071)
);

BUFx3_ASAP7_75t_L g5072 ( 
.A(n_3727),
.Y(n_5072)
);

CKINVDCx5p33_ASAP7_75t_R g5073 ( 
.A(n_3675),
.Y(n_5073)
);

CKINVDCx5p33_ASAP7_75t_R g5074 ( 
.A(n_3679),
.Y(n_5074)
);

CKINVDCx5p33_ASAP7_75t_R g5075 ( 
.A(n_3685),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4476),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4496),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_3686),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4525),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4549),
.Y(n_5080)
);

INVxp67_ASAP7_75t_L g5081 ( 
.A(n_4434),
.Y(n_5081)
);

CKINVDCx5p33_ASAP7_75t_R g5082 ( 
.A(n_3687),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_3698),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4619),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_3705),
.Y(n_5085)
);

CKINVDCx5p33_ASAP7_75t_R g5086 ( 
.A(n_3708),
.Y(n_5086)
);

INVx2_ASAP7_75t_L g5087 ( 
.A(n_4625),
.Y(n_5087)
);

CKINVDCx5p33_ASAP7_75t_R g5088 ( 
.A(n_3715),
.Y(n_5088)
);

CKINVDCx5p33_ASAP7_75t_R g5089 ( 
.A(n_3731),
.Y(n_5089)
);

CKINVDCx5p33_ASAP7_75t_R g5090 ( 
.A(n_3739),
.Y(n_5090)
);

CKINVDCx5p33_ASAP7_75t_R g5091 ( 
.A(n_3758),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4700),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4714),
.Y(n_5093)
);

NOR2xp67_ASAP7_75t_L g5094 ( 
.A(n_3829),
.B(n_3),
.Y(n_5094)
);

INVxp67_ASAP7_75t_L g5095 ( 
.A(n_4447),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4730),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4734),
.Y(n_5097)
);

CKINVDCx5p33_ASAP7_75t_R g5098 ( 
.A(n_3767),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4736),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_3773),
.Y(n_5100)
);

BUFx3_ASAP7_75t_L g5101 ( 
.A(n_3874),
.Y(n_5101)
);

CKINVDCx5p33_ASAP7_75t_R g5102 ( 
.A(n_3795),
.Y(n_5102)
);

CKINVDCx5p33_ASAP7_75t_R g5103 ( 
.A(n_3801),
.Y(n_5103)
);

CKINVDCx5p33_ASAP7_75t_R g5104 ( 
.A(n_3803),
.Y(n_5104)
);

OR2x2_ASAP7_75t_L g5105 ( 
.A(n_3576),
.B(n_3),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4767),
.Y(n_5106)
);

CKINVDCx5p33_ASAP7_75t_R g5107 ( 
.A(n_3806),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4824),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4836),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4839),
.Y(n_5110)
);

CKINVDCx16_ASAP7_75t_R g5111 ( 
.A(n_3798),
.Y(n_5111)
);

CKINVDCx20_ASAP7_75t_R g5112 ( 
.A(n_3827),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_3833),
.Y(n_5113)
);

CKINVDCx5p33_ASAP7_75t_R g5114 ( 
.A(n_3839),
.Y(n_5114)
);

CKINVDCx5p33_ASAP7_75t_R g5115 ( 
.A(n_3840),
.Y(n_5115)
);

BUFx2_ASAP7_75t_L g5116 ( 
.A(n_4628),
.Y(n_5116)
);

INVx1_ASAP7_75t_SL g5117 ( 
.A(n_4760),
.Y(n_5117)
);

CKINVDCx5p33_ASAP7_75t_R g5118 ( 
.A(n_3848),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4851),
.Y(n_5119)
);

CKINVDCx5p33_ASAP7_75t_R g5120 ( 
.A(n_3863),
.Y(n_5120)
);

CKINVDCx5p33_ASAP7_75t_R g5121 ( 
.A(n_3869),
.Y(n_5121)
);

CKINVDCx5p33_ASAP7_75t_R g5122 ( 
.A(n_3871),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_3525),
.Y(n_5123)
);

CKINVDCx5p33_ASAP7_75t_R g5124 ( 
.A(n_3878),
.Y(n_5124)
);

CKINVDCx20_ASAP7_75t_R g5125 ( 
.A(n_3830),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_3720),
.Y(n_5126)
);

CKINVDCx5p33_ASAP7_75t_R g5127 ( 
.A(n_3879),
.Y(n_5127)
);

CKINVDCx20_ASAP7_75t_R g5128 ( 
.A(n_3888),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4138),
.Y(n_5129)
);

CKINVDCx20_ASAP7_75t_R g5130 ( 
.A(n_3907),
.Y(n_5130)
);

CKINVDCx5p33_ASAP7_75t_R g5131 ( 
.A(n_3880),
.Y(n_5131)
);

CKINVDCx5p33_ASAP7_75t_R g5132 ( 
.A(n_3887),
.Y(n_5132)
);

INVx2_ASAP7_75t_L g5133 ( 
.A(n_3904),
.Y(n_5133)
);

BUFx3_ASAP7_75t_L g5134 ( 
.A(n_3883),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4138),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4692),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_3893),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4692),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_4010),
.Y(n_5139)
);

INVx1_ASAP7_75t_SL g5140 ( 
.A(n_4794),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4692),
.Y(n_5141)
);

CKINVDCx5p33_ASAP7_75t_R g5142 ( 
.A(n_3908),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4813),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4813),
.Y(n_5144)
);

CKINVDCx5p33_ASAP7_75t_R g5145 ( 
.A(n_3910),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4813),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4250),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4331),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_4501),
.Y(n_5149)
);

BUFx3_ASAP7_75t_L g5150 ( 
.A(n_3930),
.Y(n_5150)
);

OR2x2_ASAP7_75t_L g5151 ( 
.A(n_4178),
.B(n_3),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_3921),
.Y(n_5152)
);

INVx2_ASAP7_75t_L g5153 ( 
.A(n_4588),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_3927),
.Y(n_5154)
);

NOR2xp33_ASAP7_75t_L g5155 ( 
.A(n_3855),
.B(n_4),
.Y(n_5155)
);

CKINVDCx5p33_ASAP7_75t_R g5156 ( 
.A(n_3939),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4596),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_4601),
.Y(n_5158)
);

CKINVDCx20_ASAP7_75t_R g5159 ( 
.A(n_3913),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4647),
.Y(n_5160)
);

CKINVDCx5p33_ASAP7_75t_R g5161 ( 
.A(n_3942),
.Y(n_5161)
);

BUFx6f_ASAP7_75t_L g5162 ( 
.A(n_3492),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4656),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4806),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_3529),
.Y(n_5165)
);

CKINVDCx5p33_ASAP7_75t_R g5166 ( 
.A(n_3943),
.Y(n_5166)
);

CKINVDCx20_ASAP7_75t_R g5167 ( 
.A(n_3959),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_3529),
.Y(n_5168)
);

CKINVDCx5p33_ASAP7_75t_R g5169 ( 
.A(n_3948),
.Y(n_5169)
);

INVx1_ASAP7_75t_SL g5170 ( 
.A(n_3593),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_3529),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_3578),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_3964),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_3578),
.Y(n_5174)
);

CKINVDCx20_ASAP7_75t_R g5175 ( 
.A(n_3965),
.Y(n_5175)
);

HB1xp67_ASAP7_75t_L g5176 ( 
.A(n_3857),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_3578),
.Y(n_5177)
);

CKINVDCx5p33_ASAP7_75t_R g5178 ( 
.A(n_3968),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_3985),
.Y(n_5179)
);

INVx2_ASAP7_75t_L g5180 ( 
.A(n_3590),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_3986),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_3590),
.Y(n_5182)
);

CKINVDCx20_ASAP7_75t_R g5183 ( 
.A(n_3980),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_3590),
.Y(n_5184)
);

CKINVDCx5p33_ASAP7_75t_R g5185 ( 
.A(n_3997),
.Y(n_5185)
);

CKINVDCx20_ASAP7_75t_R g5186 ( 
.A(n_4017),
.Y(n_5186)
);

CKINVDCx20_ASAP7_75t_R g5187 ( 
.A(n_4024),
.Y(n_5187)
);

CKINVDCx5p33_ASAP7_75t_R g5188 ( 
.A(n_4007),
.Y(n_5188)
);

BUFx6f_ASAP7_75t_L g5189 ( 
.A(n_3609),
.Y(n_5189)
);

INVxp33_ASAP7_75t_L g5190 ( 
.A(n_4098),
.Y(n_5190)
);

INVx2_ASAP7_75t_SL g5191 ( 
.A(n_3798),
.Y(n_5191)
);

CKINVDCx5p33_ASAP7_75t_R g5192 ( 
.A(n_4034),
.Y(n_5192)
);

INVxp67_ASAP7_75t_L g5193 ( 
.A(n_4177),
.Y(n_5193)
);

CKINVDCx20_ASAP7_75t_R g5194 ( 
.A(n_4032),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_3609),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_3609),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_4046),
.Y(n_5197)
);

CKINVDCx5p33_ASAP7_75t_R g5198 ( 
.A(n_4067),
.Y(n_5198)
);

CKINVDCx5p33_ASAP7_75t_R g5199 ( 
.A(n_4075),
.Y(n_5199)
);

BUFx2_ASAP7_75t_L g5200 ( 
.A(n_4078),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_4087),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_3619),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_3619),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_3619),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_3815),
.Y(n_5205)
);

INVxp33_ASAP7_75t_L g5206 ( 
.A(n_4196),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_3815),
.Y(n_5207)
);

CKINVDCx5p33_ASAP7_75t_R g5208 ( 
.A(n_4096),
.Y(n_5208)
);

CKINVDCx5p33_ASAP7_75t_R g5209 ( 
.A(n_4101),
.Y(n_5209)
);

NOR2xp67_ASAP7_75t_L g5210 ( 
.A(n_4251),
.B(n_4),
.Y(n_5210)
);

INVxp67_ASAP7_75t_L g5211 ( 
.A(n_4595),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_4104),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_3815),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_3905),
.Y(n_5214)
);

CKINVDCx5p33_ASAP7_75t_R g5215 ( 
.A(n_4131),
.Y(n_5215)
);

CKINVDCx5p33_ASAP7_75t_R g5216 ( 
.A(n_4132),
.Y(n_5216)
);

CKINVDCx5p33_ASAP7_75t_R g5217 ( 
.A(n_4136),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_3905),
.Y(n_5218)
);

BUFx3_ASAP7_75t_L g5219 ( 
.A(n_4214),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_3905),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_3928),
.Y(n_5221)
);

CKINVDCx5p33_ASAP7_75t_R g5222 ( 
.A(n_4140),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_3928),
.Y(n_5223)
);

CKINVDCx5p33_ASAP7_75t_R g5224 ( 
.A(n_4147),
.Y(n_5224)
);

CKINVDCx20_ASAP7_75t_R g5225 ( 
.A(n_4056),
.Y(n_5225)
);

INVxp67_ASAP7_75t_L g5226 ( 
.A(n_4633),
.Y(n_5226)
);

BUFx2_ASAP7_75t_L g5227 ( 
.A(n_4165),
.Y(n_5227)
);

CKINVDCx5p33_ASAP7_75t_R g5228 ( 
.A(n_4167),
.Y(n_5228)
);

INVx1_ASAP7_75t_SL g5229 ( 
.A(n_4171),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_4172),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_3928),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_4173),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_3941),
.Y(n_5233)
);

INVx1_ASAP7_75t_SL g5234 ( 
.A(n_4591),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_3941),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_3941),
.Y(n_5236)
);

INVxp67_ASAP7_75t_SL g5237 ( 
.A(n_4771),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_3957),
.Y(n_5238)
);

CKINVDCx5p33_ASAP7_75t_R g5239 ( 
.A(n_4181),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_3957),
.Y(n_5240)
);

INVx1_ASAP7_75t_SL g5241 ( 
.A(n_3605),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_3957),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_3978),
.Y(n_5243)
);

BUFx6f_ASAP7_75t_L g5244 ( 
.A(n_3978),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_3978),
.Y(n_5245)
);

CKINVDCx5p33_ASAP7_75t_R g5246 ( 
.A(n_4198),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4035),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_4035),
.Y(n_5248)
);

CKINVDCx5p33_ASAP7_75t_R g5249 ( 
.A(n_4199),
.Y(n_5249)
);

CKINVDCx5p33_ASAP7_75t_R g5250 ( 
.A(n_4226),
.Y(n_5250)
);

BUFx6f_ASAP7_75t_L g5251 ( 
.A(n_4035),
.Y(n_5251)
);

CKINVDCx5p33_ASAP7_75t_R g5252 ( 
.A(n_4230),
.Y(n_5252)
);

CKINVDCx5p33_ASAP7_75t_R g5253 ( 
.A(n_4237),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4063),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_4246),
.Y(n_5255)
);

INVxp67_ASAP7_75t_L g5256 ( 
.A(n_3865),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_4063),
.Y(n_5257)
);

CKINVDCx5p33_ASAP7_75t_R g5258 ( 
.A(n_4259),
.Y(n_5258)
);

BUFx2_ASAP7_75t_L g5259 ( 
.A(n_4261),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_4063),
.Y(n_5260)
);

CKINVDCx5p33_ASAP7_75t_R g5261 ( 
.A(n_4278),
.Y(n_5261)
);

CKINVDCx5p33_ASAP7_75t_R g5262 ( 
.A(n_4290),
.Y(n_5262)
);

CKINVDCx16_ASAP7_75t_R g5263 ( 
.A(n_3865),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_4064),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_4064),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_4064),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_4109),
.Y(n_5267)
);

BUFx2_ASAP7_75t_SL g5268 ( 
.A(n_4350),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_4109),
.Y(n_5269)
);

BUFx3_ASAP7_75t_L g5270 ( 
.A(n_4241),
.Y(n_5270)
);

CKINVDCx5p33_ASAP7_75t_R g5271 ( 
.A(n_4305),
.Y(n_5271)
);

CKINVDCx5p33_ASAP7_75t_R g5272 ( 
.A(n_4342),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_4109),
.Y(n_5273)
);

OR2x2_ASAP7_75t_L g5274 ( 
.A(n_4289),
.B(n_4),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_4146),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_4345),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_4146),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4146),
.Y(n_5278)
);

CKINVDCx5p33_ASAP7_75t_R g5279 ( 
.A(n_4373),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4161),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4161),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4161),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4190),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4190),
.Y(n_5284)
);

BUFx2_ASAP7_75t_SL g5285 ( 
.A(n_4350),
.Y(n_5285)
);

CKINVDCx20_ASAP7_75t_R g5286 ( 
.A(n_4084),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_4190),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_4252),
.Y(n_5288)
);

CKINVDCx20_ASAP7_75t_R g5289 ( 
.A(n_4113),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_4252),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_4252),
.Y(n_5291)
);

INVxp67_ASAP7_75t_L g5292 ( 
.A(n_4791),
.Y(n_5292)
);

CKINVDCx20_ASAP7_75t_R g5293 ( 
.A(n_4123),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_4377),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4255),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4255),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_4255),
.Y(n_5297)
);

OR2x2_ASAP7_75t_L g5298 ( 
.A(n_4798),
.B(n_5),
.Y(n_5298)
);

CKINVDCx5p33_ASAP7_75t_R g5299 ( 
.A(n_4390),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_4422),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4280),
.Y(n_5301)
);

CKINVDCx5p33_ASAP7_75t_R g5302 ( 
.A(n_4442),
.Y(n_5302)
);

CKINVDCx20_ASAP7_75t_R g5303 ( 
.A(n_4133),
.Y(n_5303)
);

INVx1_ASAP7_75t_SL g5304 ( 
.A(n_3764),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4280),
.Y(n_5305)
);

CKINVDCx14_ASAP7_75t_R g5306 ( 
.A(n_4371),
.Y(n_5306)
);

CKINVDCx5p33_ASAP7_75t_R g5307 ( 
.A(n_4451),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_4879),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4882),
.Y(n_5309)
);

CKINVDCx5p33_ASAP7_75t_R g5310 ( 
.A(n_4877),
.Y(n_5310)
);

CKINVDCx20_ASAP7_75t_R g5311 ( 
.A(n_4955),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_5171),
.Y(n_5312)
);

CKINVDCx5p33_ASAP7_75t_R g5313 ( 
.A(n_4883),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_4886),
.Y(n_5314)
);

HB1xp67_ASAP7_75t_L g5315 ( 
.A(n_4915),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_5180),
.Y(n_5316)
);

INVxp67_ASAP7_75t_SL g5317 ( 
.A(n_5048),
.Y(n_5317)
);

CKINVDCx16_ASAP7_75t_R g5318 ( 
.A(n_4878),
.Y(n_5318)
);

INVxp67_ASAP7_75t_SL g5319 ( 
.A(n_5068),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4888),
.Y(n_5320)
);

HB1xp67_ASAP7_75t_L g5321 ( 
.A(n_4916),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5162),
.Y(n_5322)
);

INVxp67_ASAP7_75t_L g5323 ( 
.A(n_5268),
.Y(n_5323)
);

INVxp67_ASAP7_75t_L g5324 ( 
.A(n_5285),
.Y(n_5324)
);

INVx2_ASAP7_75t_L g5325 ( 
.A(n_5202),
.Y(n_5325)
);

INVx1_ASAP7_75t_SL g5326 ( 
.A(n_5170),
.Y(n_5326)
);

INVxp67_ASAP7_75t_SL g5327 ( 
.A(n_5072),
.Y(n_5327)
);

CKINVDCx20_ASAP7_75t_R g5328 ( 
.A(n_4998),
.Y(n_5328)
);

CKINVDCx20_ASAP7_75t_R g5329 ( 
.A(n_5005),
.Y(n_5329)
);

CKINVDCx5p33_ASAP7_75t_R g5330 ( 
.A(n_4884),
.Y(n_5330)
);

CKINVDCx5p33_ASAP7_75t_R g5331 ( 
.A(n_4889),
.Y(n_5331)
);

CKINVDCx5p33_ASAP7_75t_R g5332 ( 
.A(n_4891),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_5162),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5162),
.Y(n_5334)
);

CKINVDCx20_ASAP7_75t_R g5335 ( 
.A(n_5010),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_5189),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5189),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5189),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5244),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_4952),
.Y(n_5340)
);

BUFx6f_ASAP7_75t_SL g5341 ( 
.A(n_5063),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_5244),
.Y(n_5342)
);

CKINVDCx16_ASAP7_75t_R g5343 ( 
.A(n_4885),
.Y(n_5343)
);

CKINVDCx14_ASAP7_75t_R g5344 ( 
.A(n_4890),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5244),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5251),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5251),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5251),
.Y(n_5348)
);

INVxp67_ASAP7_75t_L g5349 ( 
.A(n_5200),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5129),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5135),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5136),
.Y(n_5352)
);

CKINVDCx5p33_ASAP7_75t_R g5353 ( 
.A(n_4953),
.Y(n_5353)
);

CKINVDCx20_ASAP7_75t_R g5354 ( 
.A(n_5011),
.Y(n_5354)
);

CKINVDCx5p33_ASAP7_75t_R g5355 ( 
.A(n_4957),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5138),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_5245),
.Y(n_5357)
);

CKINVDCx16_ASAP7_75t_R g5358 ( 
.A(n_4913),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5141),
.Y(n_5359)
);

INVxp67_ASAP7_75t_SL g5360 ( 
.A(n_5101),
.Y(n_5360)
);

CKINVDCx16_ASAP7_75t_R g5361 ( 
.A(n_4917),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5143),
.Y(n_5362)
);

INVxp33_ASAP7_75t_L g5363 ( 
.A(n_4928),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5144),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_4973),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_5146),
.Y(n_5366)
);

CKINVDCx5p33_ASAP7_75t_R g5367 ( 
.A(n_4977),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4887),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_4887),
.Y(n_5369)
);

INVxp33_ASAP7_75t_L g5370 ( 
.A(n_4936),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_4887),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_4946),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4946),
.Y(n_5373)
);

INVxp67_ASAP7_75t_SL g5374 ( 
.A(n_5134),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_4978),
.Y(n_5375)
);

CKINVDCx5p33_ASAP7_75t_R g5376 ( 
.A(n_4982),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_4946),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_4949),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_4989),
.Y(n_5379)
);

CKINVDCx5p33_ASAP7_75t_R g5380 ( 
.A(n_4990),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_5287),
.Y(n_5381)
);

INVxp67_ASAP7_75t_L g5382 ( 
.A(n_5227),
.Y(n_5382)
);

INVxp33_ASAP7_75t_L g5383 ( 
.A(n_5176),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_4949),
.Y(n_5384)
);

CKINVDCx5p33_ASAP7_75t_R g5385 ( 
.A(n_4992),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_4949),
.Y(n_5386)
);

BUFx3_ASAP7_75t_L g5387 ( 
.A(n_4873),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_4979),
.Y(n_5388)
);

CKINVDCx5p33_ASAP7_75t_R g5389 ( 
.A(n_4993),
.Y(n_5389)
);

CKINVDCx20_ASAP7_75t_R g5390 ( 
.A(n_5012),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_4979),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_4979),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_5006),
.Y(n_5393)
);

INVx1_ASAP7_75t_L g5394 ( 
.A(n_5006),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5006),
.Y(n_5395)
);

CKINVDCx20_ASAP7_75t_R g5396 ( 
.A(n_5019),
.Y(n_5396)
);

INVxp33_ASAP7_75t_SL g5397 ( 
.A(n_4874),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5040),
.Y(n_5398)
);

CKINVDCx20_ASAP7_75t_R g5399 ( 
.A(n_5022),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_4994),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_4996),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5040),
.Y(n_5402)
);

BUFx6f_ASAP7_75t_L g5403 ( 
.A(n_5040),
.Y(n_5403)
);

INVx2_ASAP7_75t_L g5404 ( 
.A(n_5071),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5071),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5071),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_4881),
.Y(n_5407)
);

HB1xp67_ASAP7_75t_L g5408 ( 
.A(n_4918),
.Y(n_5408)
);

CKINVDCx20_ASAP7_75t_R g5409 ( 
.A(n_5023),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_4941),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5165),
.Y(n_5411)
);

INVxp67_ASAP7_75t_SL g5412 ( 
.A(n_5150),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5168),
.Y(n_5413)
);

CKINVDCx20_ASAP7_75t_R g5414 ( 
.A(n_5027),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5172),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5174),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5177),
.Y(n_5417)
);

CKINVDCx20_ASAP7_75t_R g5418 ( 
.A(n_5059),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5182),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_5184),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5195),
.Y(n_5421)
);

INVxp67_ASAP7_75t_SL g5422 ( 
.A(n_5219),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5196),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5203),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_5000),
.Y(n_5425)
);

HB1xp67_ASAP7_75t_L g5426 ( 
.A(n_4920),
.Y(n_5426)
);

INVx3_ASAP7_75t_L g5427 ( 
.A(n_4950),
.Y(n_5427)
);

BUFx3_ASAP7_75t_L g5428 ( 
.A(n_4880),
.Y(n_5428)
);

CKINVDCx5p33_ASAP7_75t_R g5429 ( 
.A(n_5014),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_4950),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5204),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_5020),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5205),
.Y(n_5433)
);

INVxp33_ASAP7_75t_SL g5434 ( 
.A(n_4921),
.Y(n_5434)
);

INVxp67_ASAP7_75t_L g5435 ( 
.A(n_5259),
.Y(n_5435)
);

BUFx6f_ASAP7_75t_L g5436 ( 
.A(n_4963),
.Y(n_5436)
);

CKINVDCx20_ASAP7_75t_R g5437 ( 
.A(n_5069),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5207),
.Y(n_5438)
);

CKINVDCx20_ASAP7_75t_R g5439 ( 
.A(n_5112),
.Y(n_5439)
);

BUFx2_ASAP7_75t_L g5440 ( 
.A(n_4926),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5213),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5214),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5218),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5220),
.Y(n_5444)
);

CKINVDCx20_ASAP7_75t_R g5445 ( 
.A(n_5125),
.Y(n_5445)
);

CKINVDCx5p33_ASAP7_75t_R g5446 ( 
.A(n_5021),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5221),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5223),
.Y(n_5448)
);

CKINVDCx20_ASAP7_75t_R g5449 ( 
.A(n_5128),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5231),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_4963),
.Y(n_5451)
);

CKINVDCx20_ASAP7_75t_R g5452 ( 
.A(n_5130),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5233),
.Y(n_5453)
);

INVxp33_ASAP7_75t_SL g5454 ( 
.A(n_4923),
.Y(n_5454)
);

CKINVDCx5p33_ASAP7_75t_R g5455 ( 
.A(n_5026),
.Y(n_5455)
);

INVxp67_ASAP7_75t_SL g5456 ( 
.A(n_5270),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_5235),
.Y(n_5457)
);

CKINVDCx20_ASAP7_75t_R g5458 ( 
.A(n_5159),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5236),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5238),
.Y(n_5460)
);

CKINVDCx5p33_ASAP7_75t_R g5461 ( 
.A(n_5030),
.Y(n_5461)
);

INVxp67_ASAP7_75t_SL g5462 ( 
.A(n_4958),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_5032),
.Y(n_5463)
);

INVxp33_ASAP7_75t_L g5464 ( 
.A(n_5190),
.Y(n_5464)
);

INVxp67_ASAP7_75t_SL g5465 ( 
.A(n_4971),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_5036),
.Y(n_5466)
);

CKINVDCx5p33_ASAP7_75t_R g5467 ( 
.A(n_5045),
.Y(n_5467)
);

CKINVDCx5p33_ASAP7_75t_R g5468 ( 
.A(n_5050),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5240),
.Y(n_5469)
);

CKINVDCx5p33_ASAP7_75t_R g5470 ( 
.A(n_5053),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5242),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5243),
.Y(n_5472)
);

INVxp67_ASAP7_75t_L g5473 ( 
.A(n_5004),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5247),
.Y(n_5474)
);

INVxp33_ASAP7_75t_L g5475 ( 
.A(n_5206),
.Y(n_5475)
);

CKINVDCx20_ASAP7_75t_R g5476 ( 
.A(n_5167),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_5055),
.Y(n_5477)
);

CKINVDCx5p33_ASAP7_75t_R g5478 ( 
.A(n_5060),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5248),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5254),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5257),
.Y(n_5481)
);

CKINVDCx5p33_ASAP7_75t_R g5482 ( 
.A(n_5062),
.Y(n_5482)
);

CKINVDCx20_ASAP7_75t_R g5483 ( 
.A(n_5175),
.Y(n_5483)
);

CKINVDCx20_ASAP7_75t_R g5484 ( 
.A(n_5183),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5260),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5264),
.Y(n_5486)
);

CKINVDCx5p33_ASAP7_75t_R g5487 ( 
.A(n_5064),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5265),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5266),
.Y(n_5489)
);

CKINVDCx20_ASAP7_75t_R g5490 ( 
.A(n_5186),
.Y(n_5490)
);

CKINVDCx14_ASAP7_75t_R g5491 ( 
.A(n_5306),
.Y(n_5491)
);

BUFx3_ASAP7_75t_L g5492 ( 
.A(n_4991),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_5267),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5269),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5273),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5275),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5277),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5278),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5280),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_5281),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5282),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5283),
.Y(n_5502)
);

CKINVDCx5p33_ASAP7_75t_R g5503 ( 
.A(n_5073),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_5284),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_5288),
.Y(n_5505)
);

CKINVDCx5p33_ASAP7_75t_R g5506 ( 
.A(n_5074),
.Y(n_5506)
);

CKINVDCx20_ASAP7_75t_R g5507 ( 
.A(n_5187),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5290),
.Y(n_5508)
);

CKINVDCx5p33_ASAP7_75t_R g5509 ( 
.A(n_5075),
.Y(n_5509)
);

CKINVDCx20_ASAP7_75t_R g5510 ( 
.A(n_5194),
.Y(n_5510)
);

INVxp67_ASAP7_75t_SL g5511 ( 
.A(n_5025),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5291),
.Y(n_5512)
);

CKINVDCx5p33_ASAP7_75t_R g5513 ( 
.A(n_5078),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5295),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5296),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5297),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5301),
.Y(n_5517)
);

HB1xp67_ASAP7_75t_L g5518 ( 
.A(n_4925),
.Y(n_5518)
);

CKINVDCx5p33_ASAP7_75t_R g5519 ( 
.A(n_5082),
.Y(n_5519)
);

BUFx2_ASAP7_75t_L g5520 ( 
.A(n_4931),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5305),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_4892),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_4956),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_4959),
.Y(n_5524)
);

CKINVDCx5p33_ASAP7_75t_R g5525 ( 
.A(n_5083),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_4960),
.Y(n_5526)
);

CKINVDCx20_ASAP7_75t_R g5527 ( 
.A(n_5225),
.Y(n_5527)
);

CKINVDCx20_ASAP7_75t_R g5528 ( 
.A(n_5286),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4895),
.Y(n_5529)
);

INVxp33_ASAP7_75t_SL g5530 ( 
.A(n_4929),
.Y(n_5530)
);

CKINVDCx5p33_ASAP7_75t_R g5531 ( 
.A(n_5085),
.Y(n_5531)
);

BUFx2_ASAP7_75t_SL g5532 ( 
.A(n_5063),
.Y(n_5532)
);

CKINVDCx5p33_ASAP7_75t_R g5533 ( 
.A(n_5086),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_4897),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_4898),
.Y(n_5535)
);

CKINVDCx5p33_ASAP7_75t_R g5536 ( 
.A(n_5088),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_4900),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_4901),
.Y(n_5538)
);

INVxp67_ASAP7_75t_L g5539 ( 
.A(n_5007),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_4903),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_4905),
.Y(n_5541)
);

CKINVDCx5p33_ASAP7_75t_R g5542 ( 
.A(n_5089),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_4904),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_4910),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_4911),
.Y(n_5545)
);

CKINVDCx5p33_ASAP7_75t_R g5546 ( 
.A(n_5090),
.Y(n_5546)
);

CKINVDCx5p33_ASAP7_75t_R g5547 ( 
.A(n_5091),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_4912),
.Y(n_5548)
);

CKINVDCx5p33_ASAP7_75t_R g5549 ( 
.A(n_5098),
.Y(n_5549)
);

CKINVDCx5p33_ASAP7_75t_R g5550 ( 
.A(n_5100),
.Y(n_5550)
);

CKINVDCx20_ASAP7_75t_R g5551 ( 
.A(n_5289),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_4914),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4919),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_4924),
.Y(n_5554)
);

CKINVDCx5p33_ASAP7_75t_R g5555 ( 
.A(n_5102),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_4927),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4933),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_5103),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_4934),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4937),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_4939),
.Y(n_5561)
);

CKINVDCx5p33_ASAP7_75t_R g5562 ( 
.A(n_5104),
.Y(n_5562)
);

CKINVDCx16_ASAP7_75t_R g5563 ( 
.A(n_4935),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_5001),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_4942),
.Y(n_5565)
);

INVxp67_ASAP7_75t_L g5566 ( 
.A(n_5029),
.Y(n_5566)
);

HB1xp67_ASAP7_75t_L g5567 ( 
.A(n_4932),
.Y(n_5567)
);

CKINVDCx5p33_ASAP7_75t_R g5568 ( 
.A(n_5107),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_4944),
.Y(n_5569)
);

CKINVDCx5p33_ASAP7_75t_R g5570 ( 
.A(n_5113),
.Y(n_5570)
);

INVxp67_ASAP7_75t_L g5571 ( 
.A(n_5116),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_4945),
.Y(n_5572)
);

CKINVDCx20_ASAP7_75t_R g5573 ( 
.A(n_5293),
.Y(n_5573)
);

INVxp67_ASAP7_75t_SL g5574 ( 
.A(n_5043),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_4947),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_4954),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_4962),
.Y(n_5577)
);

INVxp67_ASAP7_75t_SL g5578 ( 
.A(n_5013),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_4965),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_5041),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_4966),
.Y(n_5581)
);

CKINVDCx5p33_ASAP7_75t_R g5582 ( 
.A(n_5114),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_4968),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_4969),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_4974),
.Y(n_5585)
);

CKINVDCx5p33_ASAP7_75t_R g5586 ( 
.A(n_5115),
.Y(n_5586)
);

INVxp67_ASAP7_75t_SL g5587 ( 
.A(n_5049),
.Y(n_5587)
);

CKINVDCx16_ASAP7_75t_R g5588 ( 
.A(n_4938),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_4975),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_4976),
.Y(n_5590)
);

HB1xp67_ASAP7_75t_L g5591 ( 
.A(n_4896),
.Y(n_5591)
);

CKINVDCx16_ASAP7_75t_R g5592 ( 
.A(n_4948),
.Y(n_5592)
);

CKINVDCx20_ASAP7_75t_R g5593 ( 
.A(n_5303),
.Y(n_5593)
);

INVxp33_ASAP7_75t_SL g5594 ( 
.A(n_4902),
.Y(n_5594)
);

CKINVDCx5p33_ASAP7_75t_R g5595 ( 
.A(n_5118),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_4980),
.Y(n_5596)
);

INVx1_ASAP7_75t_SL g5597 ( 
.A(n_5229),
.Y(n_5597)
);

CKINVDCx5p33_ASAP7_75t_R g5598 ( 
.A(n_5120),
.Y(n_5598)
);

INVxp67_ASAP7_75t_SL g5599 ( 
.A(n_5094),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_4983),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_4984),
.Y(n_5601)
);

INVxp33_ASAP7_75t_SL g5602 ( 
.A(n_4906),
.Y(n_5602)
);

CKINVDCx5p33_ASAP7_75t_R g5603 ( 
.A(n_5121),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_4985),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_4987),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_4988),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_4995),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_4997),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_4999),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_5002),
.Y(n_5610)
);

HB1xp67_ASAP7_75t_L g5611 ( 
.A(n_5122),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5008),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5009),
.Y(n_5613)
);

CKINVDCx20_ASAP7_75t_R g5614 ( 
.A(n_4907),
.Y(n_5614)
);

CKINVDCx5p33_ASAP7_75t_R g5615 ( 
.A(n_5124),
.Y(n_5615)
);

INVxp33_ASAP7_75t_SL g5616 ( 
.A(n_4908),
.Y(n_5616)
);

CKINVDCx5p33_ASAP7_75t_R g5617 ( 
.A(n_5127),
.Y(n_5617)
);

CKINVDCx20_ASAP7_75t_R g5618 ( 
.A(n_5234),
.Y(n_5618)
);

INVxp33_ASAP7_75t_L g5619 ( 
.A(n_5155),
.Y(n_5619)
);

INVxp67_ASAP7_75t_SL g5620 ( 
.A(n_5210),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5015),
.Y(n_5621)
);

CKINVDCx5p33_ASAP7_75t_R g5622 ( 
.A(n_5131),
.Y(n_5622)
);

CKINVDCx5p33_ASAP7_75t_R g5623 ( 
.A(n_5132),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_5137),
.Y(n_5624)
);

HB1xp67_ASAP7_75t_L g5625 ( 
.A(n_5142),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5016),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5017),
.Y(n_5627)
);

INVxp67_ASAP7_75t_SL g5628 ( 
.A(n_4909),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5018),
.Y(n_5629)
);

INVxp67_ASAP7_75t_SL g5630 ( 
.A(n_4961),
.Y(n_5630)
);

BUFx3_ASAP7_75t_L g5631 ( 
.A(n_5024),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5028),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5042),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5031),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5033),
.Y(n_5635)
);

INVx4_ASAP7_75t_R g5636 ( 
.A(n_4876),
.Y(n_5636)
);

CKINVDCx20_ASAP7_75t_R g5637 ( 
.A(n_5241),
.Y(n_5637)
);

CKINVDCx20_ASAP7_75t_R g5638 ( 
.A(n_5304),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5034),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5035),
.Y(n_5640)
);

CKINVDCx5p33_ASAP7_75t_R g5641 ( 
.A(n_5145),
.Y(n_5641)
);

INVx2_ASAP7_75t_L g5642 ( 
.A(n_5044),
.Y(n_5642)
);

CKINVDCx16_ASAP7_75t_R g5643 ( 
.A(n_4951),
.Y(n_5643)
);

INVxp67_ASAP7_75t_SL g5644 ( 
.A(n_5256),
.Y(n_5644)
);

INVxp67_ASAP7_75t_SL g5645 ( 
.A(n_5292),
.Y(n_5645)
);

BUFx3_ASAP7_75t_L g5646 ( 
.A(n_5037),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5046),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5047),
.Y(n_5648)
);

INVxp67_ASAP7_75t_L g5649 ( 
.A(n_4930),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_5051),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5052),
.Y(n_5651)
);

CKINVDCx5p33_ASAP7_75t_R g5652 ( 
.A(n_5152),
.Y(n_5652)
);

CKINVDCx20_ASAP7_75t_R g5653 ( 
.A(n_5154),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5054),
.Y(n_5654)
);

BUFx2_ASAP7_75t_SL g5655 ( 
.A(n_4986),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5056),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5057),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5058),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5061),
.Y(n_5659)
);

CKINVDCx5p33_ASAP7_75t_R g5660 ( 
.A(n_5156),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_5077),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5065),
.Y(n_5662)
);

CKINVDCx5p33_ASAP7_75t_R g5663 ( 
.A(n_5161),
.Y(n_5663)
);

CKINVDCx5p33_ASAP7_75t_R g5664 ( 
.A(n_5166),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5066),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5087),
.Y(n_5666)
);

CKINVDCx20_ASAP7_75t_R g5667 ( 
.A(n_5169),
.Y(n_5667)
);

INVx2_ASAP7_75t_L g5668 ( 
.A(n_5123),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5067),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5076),
.Y(n_5670)
);

INVxp33_ASAP7_75t_L g5671 ( 
.A(n_4943),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5079),
.Y(n_5672)
);

CKINVDCx5p33_ASAP7_75t_R g5673 ( 
.A(n_5173),
.Y(n_5673)
);

CKINVDCx5p33_ASAP7_75t_R g5674 ( 
.A(n_5178),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5080),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5084),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5092),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_4894),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5093),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5096),
.Y(n_5680)
);

CKINVDCx20_ASAP7_75t_R g5681 ( 
.A(n_5179),
.Y(n_5681)
);

INVxp33_ASAP7_75t_L g5682 ( 
.A(n_5038),
.Y(n_5682)
);

CKINVDCx5p33_ASAP7_75t_R g5683 ( 
.A(n_5181),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5097),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5099),
.Y(n_5685)
);

CKINVDCx5p33_ASAP7_75t_R g5686 ( 
.A(n_5185),
.Y(n_5686)
);

CKINVDCx20_ASAP7_75t_R g5687 ( 
.A(n_5188),
.Y(n_5687)
);

CKINVDCx5p33_ASAP7_75t_R g5688 ( 
.A(n_5192),
.Y(n_5688)
);

CKINVDCx16_ASAP7_75t_R g5689 ( 
.A(n_4964),
.Y(n_5689)
);

INVxp33_ASAP7_75t_SL g5690 ( 
.A(n_5197),
.Y(n_5690)
);

BUFx3_ASAP7_75t_L g5691 ( 
.A(n_5106),
.Y(n_5691)
);

CKINVDCx5p33_ASAP7_75t_R g5692 ( 
.A(n_5198),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5108),
.Y(n_5693)
);

INVxp33_ASAP7_75t_SL g5694 ( 
.A(n_5199),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5109),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5110),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5119),
.Y(n_5697)
);

BUFx2_ASAP7_75t_L g5698 ( 
.A(n_5201),
.Y(n_5698)
);

INVxp33_ASAP7_75t_SL g5699 ( 
.A(n_5208),
.Y(n_5699)
);

CKINVDCx20_ASAP7_75t_R g5700 ( 
.A(n_5209),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_5126),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5133),
.Y(n_5702)
);

CKINVDCx5p33_ASAP7_75t_R g5703 ( 
.A(n_5212),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5139),
.Y(n_5704)
);

BUFx2_ASAP7_75t_SL g5705 ( 
.A(n_5003),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5153),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5164),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5147),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5148),
.Y(n_5709)
);

CKINVDCx20_ASAP7_75t_R g5710 ( 
.A(n_5215),
.Y(n_5710)
);

CKINVDCx16_ASAP7_75t_R g5711 ( 
.A(n_4972),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5149),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5157),
.Y(n_5713)
);

BUFx6f_ASAP7_75t_L g5714 ( 
.A(n_5158),
.Y(n_5714)
);

CKINVDCx20_ASAP7_75t_R g5715 ( 
.A(n_5216),
.Y(n_5715)
);

INVxp67_ASAP7_75t_SL g5716 ( 
.A(n_5193),
.Y(n_5716)
);

INVxp33_ASAP7_75t_SL g5717 ( 
.A(n_5217),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5160),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5163),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5237),
.Y(n_5720)
);

CKINVDCx20_ASAP7_75t_R g5721 ( 
.A(n_5222),
.Y(n_5721)
);

INVxp67_ASAP7_75t_SL g5722 ( 
.A(n_5211),
.Y(n_5722)
);

CKINVDCx14_ASAP7_75t_R g5723 ( 
.A(n_4875),
.Y(n_5723)
);

INVxp67_ASAP7_75t_SL g5724 ( 
.A(n_5226),
.Y(n_5724)
);

CKINVDCx20_ASAP7_75t_R g5725 ( 
.A(n_5224),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_4967),
.Y(n_5726)
);

CKINVDCx5p33_ASAP7_75t_R g5727 ( 
.A(n_5228),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_5307),
.Y(n_5728)
);

INVxp67_ASAP7_75t_SL g5729 ( 
.A(n_4899),
.Y(n_5729)
);

CKINVDCx20_ASAP7_75t_R g5730 ( 
.A(n_5230),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_4981),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5232),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5239),
.Y(n_5733)
);

INVxp67_ASAP7_75t_L g5734 ( 
.A(n_5191),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5246),
.Y(n_5735)
);

CKINVDCx20_ASAP7_75t_R g5736 ( 
.A(n_5249),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_5250),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5252),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_5253),
.Y(n_5739)
);

CKINVDCx5p33_ASAP7_75t_R g5740 ( 
.A(n_5255),
.Y(n_5740)
);

BUFx2_ASAP7_75t_L g5741 ( 
.A(n_5258),
.Y(n_5741)
);

CKINVDCx20_ASAP7_75t_R g5742 ( 
.A(n_5261),
.Y(n_5742)
);

CKINVDCx20_ASAP7_75t_R g5743 ( 
.A(n_5262),
.Y(n_5743)
);

CKINVDCx20_ASAP7_75t_R g5744 ( 
.A(n_5271),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5272),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5276),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5279),
.Y(n_5747)
);

CKINVDCx5p33_ASAP7_75t_R g5748 ( 
.A(n_5294),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5299),
.Y(n_5749)
);

CKINVDCx5p33_ASAP7_75t_R g5750 ( 
.A(n_5300),
.Y(n_5750)
);

CKINVDCx5p33_ASAP7_75t_R g5751 ( 
.A(n_5302),
.Y(n_5751)
);

INVxp67_ASAP7_75t_SL g5752 ( 
.A(n_5081),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_5105),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5095),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_4894),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_4922),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_4922),
.Y(n_5757)
);

CKINVDCx20_ASAP7_75t_R g5758 ( 
.A(n_5111),
.Y(n_5758)
);

CKINVDCx5p33_ASAP7_75t_R g5759 ( 
.A(n_5263),
.Y(n_5759)
);

BUFx3_ASAP7_75t_L g5760 ( 
.A(n_5151),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5298),
.Y(n_5761)
);

CKINVDCx20_ASAP7_75t_R g5762 ( 
.A(n_4940),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5274),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5039),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_4970),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5070),
.Y(n_5766)
);

INVxp67_ASAP7_75t_SL g5767 ( 
.A(n_4893),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5117),
.Y(n_5768)
);

CKINVDCx20_ASAP7_75t_R g5769 ( 
.A(n_5140),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_4879),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_4879),
.Y(n_5771)
);

BUFx2_ASAP7_75t_SL g5772 ( 
.A(n_4878),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_4879),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_4879),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_4879),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_4879),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_4879),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_4879),
.Y(n_5778)
);

CKINVDCx5p33_ASAP7_75t_R g5779 ( 
.A(n_4877),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_4879),
.Y(n_5780)
);

BUFx2_ASAP7_75t_L g5781 ( 
.A(n_4926),
.Y(n_5781)
);

INVxp33_ASAP7_75t_SL g5782 ( 
.A(n_4874),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_4879),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_4879),
.Y(n_5784)
);

CKINVDCx20_ASAP7_75t_R g5785 ( 
.A(n_4955),
.Y(n_5785)
);

INVxp67_ASAP7_75t_SL g5786 ( 
.A(n_5048),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_4879),
.Y(n_5787)
);

CKINVDCx20_ASAP7_75t_R g5788 ( 
.A(n_4955),
.Y(n_5788)
);

CKINVDCx5p33_ASAP7_75t_R g5789 ( 
.A(n_4877),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_4879),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_4879),
.Y(n_5791)
);

CKINVDCx14_ASAP7_75t_R g5792 ( 
.A(n_4890),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_4879),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_4879),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_4879),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_4879),
.Y(n_5796)
);

CKINVDCx14_ASAP7_75t_R g5797 ( 
.A(n_4890),
.Y(n_5797)
);

BUFx6f_ASAP7_75t_L g5798 ( 
.A(n_4887),
.Y(n_5798)
);

CKINVDCx16_ASAP7_75t_R g5799 ( 
.A(n_4878),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_4877),
.Y(n_5800)
);

CKINVDCx20_ASAP7_75t_R g5801 ( 
.A(n_4955),
.Y(n_5801)
);

CKINVDCx5p33_ASAP7_75t_R g5802 ( 
.A(n_4877),
.Y(n_5802)
);

CKINVDCx5p33_ASAP7_75t_R g5803 ( 
.A(n_4877),
.Y(n_5803)
);

INVx2_ASAP7_75t_L g5804 ( 
.A(n_5171),
.Y(n_5804)
);

CKINVDCx5p33_ASAP7_75t_R g5805 ( 
.A(n_4877),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_4877),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_4879),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_4879),
.Y(n_5808)
);

CKINVDCx20_ASAP7_75t_R g5809 ( 
.A(n_4955),
.Y(n_5809)
);

CKINVDCx5p33_ASAP7_75t_R g5810 ( 
.A(n_4877),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_4879),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_4879),
.Y(n_5812)
);

CKINVDCx5p33_ASAP7_75t_R g5813 ( 
.A(n_4877),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_4879),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_4877),
.Y(n_5815)
);

INVx5_ASAP7_75t_L g5816 ( 
.A(n_5343),
.Y(n_5816)
);

NOR2x1_ASAP7_75t_L g5817 ( 
.A(n_5732),
.B(n_4269),
.Y(n_5817)
);

BUFx3_ASAP7_75t_L g5818 ( 
.A(n_5387),
.Y(n_5818)
);

INVx4_ASAP7_75t_L g5819 ( 
.A(n_5340),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5631),
.Y(n_5820)
);

BUFx6f_ASAP7_75t_L g5821 ( 
.A(n_5403),
.Y(n_5821)
);

BUFx3_ASAP7_75t_L g5822 ( 
.A(n_5428),
.Y(n_5822)
);

CKINVDCx6p67_ASAP7_75t_R g5823 ( 
.A(n_5341),
.Y(n_5823)
);

NAND2xp5_ASAP7_75t_L g5824 ( 
.A(n_5628),
.B(n_4280),
.Y(n_5824)
);

CKINVDCx5p33_ASAP7_75t_R g5825 ( 
.A(n_5353),
.Y(n_5825)
);

INVx3_ASAP7_75t_L g5826 ( 
.A(n_5492),
.Y(n_5826)
);

BUFx6f_ASAP7_75t_L g5827 ( 
.A(n_5403),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5404),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5646),
.Y(n_5829)
);

NOR2xp33_ASAP7_75t_L g5830 ( 
.A(n_5733),
.B(n_4463),
.Y(n_5830)
);

OA21x2_ASAP7_75t_L g5831 ( 
.A1(n_5308),
.A2(n_3475),
.B(n_4058),
.Y(n_5831)
);

OAI21x1_ASAP7_75t_L g5832 ( 
.A1(n_5407),
.A2(n_3481),
.B(n_3477),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5691),
.Y(n_5833)
);

AOI22xp5_ASAP7_75t_L g5834 ( 
.A1(n_5349),
.A2(n_5435),
.B1(n_5382),
.B2(n_5752),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5577),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5668),
.Y(n_5836)
);

NOR2xp33_ASAP7_75t_L g5837 ( 
.A(n_5735),
.B(n_4485),
.Y(n_5837)
);

HB1xp67_ASAP7_75t_L g5838 ( 
.A(n_5326),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5579),
.Y(n_5839)
);

INVxp67_ASAP7_75t_L g5840 ( 
.A(n_5767),
.Y(n_5840)
);

BUFx2_ASAP7_75t_L g5841 ( 
.A(n_5762),
.Y(n_5841)
);

INVx2_ASAP7_75t_L g5842 ( 
.A(n_5436),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5581),
.Y(n_5843)
);

INVx2_ASAP7_75t_L g5844 ( 
.A(n_5436),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_5436),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5451),
.Y(n_5846)
);

OAI21x1_ASAP7_75t_L g5847 ( 
.A1(n_5522),
.A2(n_3516),
.B(n_3503),
.Y(n_5847)
);

CKINVDCx5p33_ASAP7_75t_R g5848 ( 
.A(n_5355),
.Y(n_5848)
);

OA21x2_ASAP7_75t_L g5849 ( 
.A1(n_5309),
.A2(n_4378),
.B(n_3915),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5451),
.Y(n_5850)
);

BUFx6f_ASAP7_75t_L g5851 ( 
.A(n_5403),
.Y(n_5851)
);

OAI22xp5_ASAP7_75t_L g5852 ( 
.A1(n_5619),
.A2(n_3476),
.B1(n_4538),
.B2(n_4492),
.Y(n_5852)
);

BUFx6f_ASAP7_75t_L g5853 ( 
.A(n_5798),
.Y(n_5853)
);

NAND2xp5_ASAP7_75t_L g5854 ( 
.A(n_5630),
.B(n_4282),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5583),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5464),
.B(n_4371),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5584),
.Y(n_5857)
);

INVx5_ASAP7_75t_L g5858 ( 
.A(n_5358),
.Y(n_5858)
);

BUFx3_ASAP7_75t_L g5859 ( 
.A(n_5451),
.Y(n_5859)
);

BUFx2_ASAP7_75t_L g5860 ( 
.A(n_5769),
.Y(n_5860)
);

OA21x2_ASAP7_75t_L g5861 ( 
.A1(n_5314),
.A2(n_3471),
.B(n_3470),
.Y(n_5861)
);

AND2x4_ASAP7_75t_L g5862 ( 
.A(n_5462),
.B(n_4396),
.Y(n_5862)
);

HB1xp67_ASAP7_75t_L g5863 ( 
.A(n_5597),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5585),
.Y(n_5864)
);

AOI22xp5_ASAP7_75t_L g5865 ( 
.A1(n_5729),
.A2(n_3601),
.B1(n_3629),
.B2(n_3564),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5312),
.Y(n_5866)
);

INVx6_ASAP7_75t_L g5867 ( 
.A(n_5361),
.Y(n_5867)
);

BUFx6f_ASAP7_75t_L g5868 ( 
.A(n_5798),
.Y(n_5868)
);

AND2x4_ASAP7_75t_L g5869 ( 
.A(n_5465),
.B(n_4446),
.Y(n_5869)
);

BUFx6f_ASAP7_75t_L g5870 ( 
.A(n_5798),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5589),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5590),
.Y(n_5872)
);

INVxp33_ASAP7_75t_SL g5873 ( 
.A(n_5532),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5596),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5600),
.Y(n_5875)
);

INVx4_ASAP7_75t_L g5876 ( 
.A(n_5365),
.Y(n_5876)
);

INVx5_ASAP7_75t_L g5877 ( 
.A(n_5563),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5601),
.Y(n_5878)
);

BUFx3_ASAP7_75t_L g5879 ( 
.A(n_5653),
.Y(n_5879)
);

CKINVDCx6p67_ASAP7_75t_R g5880 ( 
.A(n_5341),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5604),
.Y(n_5881)
);

AOI22xp5_ASAP7_75t_L g5882 ( 
.A1(n_5738),
.A2(n_3709),
.B1(n_3778),
.B2(n_3691),
.Y(n_5882)
);

AND2x2_ASAP7_75t_SL g5883 ( 
.A(n_5588),
.B(n_4282),
.Y(n_5883)
);

INVx6_ASAP7_75t_L g5884 ( 
.A(n_5592),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5605),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5606),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5607),
.Y(n_5887)
);

AOI22xp5_ASAP7_75t_L g5888 ( 
.A1(n_5745),
.A2(n_3845),
.B1(n_3849),
.B2(n_3844),
.Y(n_5888)
);

BUFx6f_ASAP7_75t_L g5889 ( 
.A(n_5714),
.Y(n_5889)
);

INVx3_ASAP7_75t_L g5890 ( 
.A(n_5427),
.Y(n_5890)
);

NOR2xp33_ASAP7_75t_L g5891 ( 
.A(n_5746),
.B(n_4558),
.Y(n_5891)
);

OAI22xp5_ASAP7_75t_L g5892 ( 
.A1(n_5761),
.A2(n_4569),
.B1(n_4576),
.B2(n_4562),
.Y(n_5892)
);

BUFx6f_ASAP7_75t_L g5893 ( 
.A(n_5714),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5316),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5608),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5609),
.Y(n_5896)
);

CKINVDCx5p33_ASAP7_75t_R g5897 ( 
.A(n_5367),
.Y(n_5897)
);

BUFx3_ASAP7_75t_L g5898 ( 
.A(n_5667),
.Y(n_5898)
);

INVx2_ASAP7_75t_SL g5899 ( 
.A(n_5760),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5610),
.Y(n_5900)
);

BUFx6f_ASAP7_75t_L g5901 ( 
.A(n_5714),
.Y(n_5901)
);

INVx2_ASAP7_75t_L g5902 ( 
.A(n_5325),
.Y(n_5902)
);

AND2x6_ASAP7_75t_L g5903 ( 
.A(n_5747),
.B(n_4462),
.Y(n_5903)
);

AND2x4_ASAP7_75t_L g5904 ( 
.A(n_5511),
.B(n_4486),
.Y(n_5904)
);

BUFx6f_ASAP7_75t_L g5905 ( 
.A(n_5430),
.Y(n_5905)
);

INVx2_ASAP7_75t_L g5906 ( 
.A(n_5357),
.Y(n_5906)
);

AND2x4_ASAP7_75t_L g5907 ( 
.A(n_5574),
.B(n_4498),
.Y(n_5907)
);

INVx3_ASAP7_75t_L g5908 ( 
.A(n_5427),
.Y(n_5908)
);

AND2x4_ASAP7_75t_L g5909 ( 
.A(n_5317),
.B(n_4504),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5612),
.Y(n_5910)
);

AND2x6_ASAP7_75t_L g5911 ( 
.A(n_5749),
.B(n_4523),
.Y(n_5911)
);

BUFx6f_ASAP7_75t_L g5912 ( 
.A(n_5381),
.Y(n_5912)
);

AND2x4_ASAP7_75t_L g5913 ( 
.A(n_5319),
.B(n_4556),
.Y(n_5913)
);

BUFx3_ASAP7_75t_L g5914 ( 
.A(n_5681),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5804),
.Y(n_5915)
);

BUFx6f_ASAP7_75t_L g5916 ( 
.A(n_5564),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5613),
.Y(n_5917)
);

INVx3_ASAP7_75t_L g5918 ( 
.A(n_5541),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5621),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5626),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5627),
.Y(n_5921)
);

INVx3_ASAP7_75t_L g5922 ( 
.A(n_5322),
.Y(n_5922)
);

BUFx6f_ASAP7_75t_L g5923 ( 
.A(n_5580),
.Y(n_5923)
);

BUFx6f_ASAP7_75t_L g5924 ( 
.A(n_5633),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5578),
.B(n_4282),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5629),
.Y(n_5926)
);

INVx2_ASAP7_75t_L g5927 ( 
.A(n_5642),
.Y(n_5927)
);

INVx3_ASAP7_75t_L g5928 ( 
.A(n_5333),
.Y(n_5928)
);

CKINVDCx16_ASAP7_75t_R g5929 ( 
.A(n_5643),
.Y(n_5929)
);

AND2x4_ASAP7_75t_L g5930 ( 
.A(n_5327),
.B(n_4567),
.Y(n_5930)
);

INVx3_ASAP7_75t_L g5931 ( 
.A(n_5334),
.Y(n_5931)
);

AND2x2_ASAP7_75t_SL g5932 ( 
.A(n_5698),
.B(n_4304),
.Y(n_5932)
);

BUFx6f_ASAP7_75t_L g5933 ( 
.A(n_5661),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5632),
.Y(n_5934)
);

BUFx6f_ASAP7_75t_L g5935 ( 
.A(n_5666),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5514),
.Y(n_5936)
);

BUFx2_ASAP7_75t_L g5937 ( 
.A(n_5618),
.Y(n_5937)
);

AND2x2_ASAP7_75t_L g5938 ( 
.A(n_5475),
.B(n_4448),
.Y(n_5938)
);

INVx3_ASAP7_75t_L g5939 ( 
.A(n_5336),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5634),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5350),
.Y(n_5941)
);

OAI22xp5_ASAP7_75t_L g5942 ( 
.A1(n_5763),
.A2(n_4587),
.B1(n_4593),
.B2(n_4584),
.Y(n_5942)
);

INVx6_ASAP7_75t_L g5943 ( 
.A(n_5689),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5635),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5351),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5352),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5639),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5356),
.Y(n_5948)
);

INVx1_ASAP7_75t_L g5949 ( 
.A(n_5640),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_5375),
.Y(n_5950)
);

OAI22xp5_ASAP7_75t_L g5951 ( 
.A1(n_5753),
.A2(n_4615),
.B1(n_4616),
.B2(n_4608),
.Y(n_5951)
);

BUFx3_ASAP7_75t_L g5952 ( 
.A(n_5687),
.Y(n_5952)
);

INVx2_ASAP7_75t_L g5953 ( 
.A(n_5359),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5647),
.Y(n_5954)
);

BUFx6f_ASAP7_75t_L g5955 ( 
.A(n_5337),
.Y(n_5955)
);

NAND2xp5_ASAP7_75t_L g5956 ( 
.A(n_5587),
.B(n_4304),
.Y(n_5956)
);

BUFx6f_ASAP7_75t_L g5957 ( 
.A(n_5338),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_SL g5958 ( 
.A(n_5765),
.B(n_4304),
.Y(n_5958)
);

INVx6_ASAP7_75t_L g5959 ( 
.A(n_5711),
.Y(n_5959)
);

INVx2_ASAP7_75t_L g5960 ( 
.A(n_5362),
.Y(n_5960)
);

NOR2xp33_ASAP7_75t_L g5961 ( 
.A(n_5728),
.B(n_4639),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5364),
.Y(n_5962)
);

BUFx2_ASAP7_75t_L g5963 ( 
.A(n_5637),
.Y(n_5963)
);

OA21x2_ASAP7_75t_L g5964 ( 
.A1(n_5320),
.A2(n_3480),
.B(n_3479),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5648),
.Y(n_5965)
);

BUFx12f_ASAP7_75t_L g5966 ( 
.A(n_5759),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5650),
.Y(n_5967)
);

INVx2_ASAP7_75t_L g5968 ( 
.A(n_5366),
.Y(n_5968)
);

INVx3_ASAP7_75t_L g5969 ( 
.A(n_5339),
.Y(n_5969)
);

BUFx6f_ASAP7_75t_L g5970 ( 
.A(n_5342),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5701),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_SL g5972 ( 
.A(n_5766),
.B(n_4387),
.Y(n_5972)
);

INVx2_ASAP7_75t_L g5973 ( 
.A(n_5702),
.Y(n_5973)
);

INVx6_ASAP7_75t_L g5974 ( 
.A(n_5318),
.Y(n_5974)
);

AND2x4_ASAP7_75t_L g5975 ( 
.A(n_5360),
.B(n_4598),
.Y(n_5975)
);

CKINVDCx8_ASAP7_75t_R g5976 ( 
.A(n_5772),
.Y(n_5976)
);

BUFx12f_ASAP7_75t_L g5977 ( 
.A(n_5376),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_5704),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_L g5979 ( 
.A(n_5599),
.B(n_5620),
.Y(n_5979)
);

OA21x2_ASAP7_75t_L g5980 ( 
.A1(n_5770),
.A2(n_3498),
.B(n_3482),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5651),
.Y(n_5981)
);

BUFx6f_ASAP7_75t_L g5982 ( 
.A(n_5345),
.Y(n_5982)
);

AND2x6_ASAP7_75t_L g5983 ( 
.A(n_5726),
.B(n_4653),
.Y(n_5983)
);

OA21x2_ASAP7_75t_L g5984 ( 
.A1(n_5771),
.A2(n_3505),
.B(n_3500),
.Y(n_5984)
);

INVx3_ASAP7_75t_L g5985 ( 
.A(n_5346),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5654),
.Y(n_5986)
);

AND2x4_ASAP7_75t_SL g5987 ( 
.A(n_5638),
.B(n_3541),
.Y(n_5987)
);

BUFx6f_ASAP7_75t_L g5988 ( 
.A(n_5347),
.Y(n_5988)
);

BUFx6f_ASAP7_75t_L g5989 ( 
.A(n_5348),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5656),
.Y(n_5990)
);

AOI22xp5_ASAP7_75t_L g5991 ( 
.A1(n_5764),
.A2(n_4130),
.B1(n_4201),
.B2(n_4014),
.Y(n_5991)
);

BUFx3_ASAP7_75t_L g5992 ( 
.A(n_5700),
.Y(n_5992)
);

INVx3_ASAP7_75t_L g5993 ( 
.A(n_5368),
.Y(n_5993)
);

AND2x4_ASAP7_75t_L g5994 ( 
.A(n_5374),
.B(n_4679),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5657),
.Y(n_5995)
);

BUFx6f_ASAP7_75t_L g5996 ( 
.A(n_5369),
.Y(n_5996)
);

BUFx6f_ASAP7_75t_L g5997 ( 
.A(n_5371),
.Y(n_5997)
);

AOI22xp5_ASAP7_75t_L g5998 ( 
.A1(n_5720),
.A2(n_4254),
.B1(n_4348),
.B2(n_4208),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5706),
.Y(n_5999)
);

OAI22xp5_ASAP7_75t_SL g6000 ( 
.A1(n_5758),
.A2(n_3903),
.B1(n_4052),
.B2(n_3748),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5658),
.Y(n_6001)
);

BUFx6f_ASAP7_75t_L g6002 ( 
.A(n_5372),
.Y(n_6002)
);

INVx2_ASAP7_75t_L g6003 ( 
.A(n_5707),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5659),
.Y(n_6004)
);

BUFx6f_ASAP7_75t_L g6005 ( 
.A(n_5373),
.Y(n_6005)
);

NAND2x1p5_ASAP7_75t_L g6006 ( 
.A(n_5741),
.B(n_4739),
.Y(n_6006)
);

NOR2xp33_ASAP7_75t_L g6007 ( 
.A(n_5410),
.B(n_4645),
.Y(n_6007)
);

OAI22xp5_ASAP7_75t_L g6008 ( 
.A1(n_5671),
.A2(n_4663),
.B1(n_4695),
.B2(n_4659),
.Y(n_6008)
);

INVx2_ASAP7_75t_L g6009 ( 
.A(n_5411),
.Y(n_6009)
);

HB1xp67_ASAP7_75t_L g6010 ( 
.A(n_5723),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5662),
.Y(n_6011)
);

BUFx6f_ASAP7_75t_L g6012 ( 
.A(n_5377),
.Y(n_6012)
);

OAI22xp5_ASAP7_75t_L g6013 ( 
.A1(n_5682),
.A2(n_4698),
.B1(n_4711),
.B2(n_4696),
.Y(n_6013)
);

BUFx2_ASAP7_75t_L g6014 ( 
.A(n_5768),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5665),
.Y(n_6015)
);

OAI21x1_ASAP7_75t_L g6016 ( 
.A1(n_5773),
.A2(n_3626),
.B(n_3592),
.Y(n_6016)
);

OA21x2_ASAP7_75t_L g6017 ( 
.A1(n_5774),
.A2(n_3510),
.B(n_3508),
.Y(n_6017)
);

AND2x6_ASAP7_75t_L g6018 ( 
.A(n_5731),
.B(n_4776),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5669),
.Y(n_6019)
);

AOI22xp5_ASAP7_75t_L g6020 ( 
.A1(n_5716),
.A2(n_4393),
.B1(n_4417),
.B2(n_4366),
.Y(n_6020)
);

AOI22xp5_ASAP7_75t_L g6021 ( 
.A1(n_5722),
.A2(n_4433),
.B1(n_4507),
.B2(n_4425),
.Y(n_6021)
);

BUFx6f_ASAP7_75t_L g6022 ( 
.A(n_5378),
.Y(n_6022)
);

NAND2xp5_ASAP7_75t_SL g6023 ( 
.A(n_5323),
.B(n_4387),
.Y(n_6023)
);

BUFx6f_ASAP7_75t_L g6024 ( 
.A(n_5384),
.Y(n_6024)
);

NOR2xp33_ASAP7_75t_L g6025 ( 
.A(n_5690),
.B(n_4716),
.Y(n_6025)
);

INVx2_ASAP7_75t_L g6026 ( 
.A(n_5413),
.Y(n_6026)
);

AND2x6_ASAP7_75t_L g6027 ( 
.A(n_5754),
.B(n_4808),
.Y(n_6027)
);

INVxp67_ASAP7_75t_L g6028 ( 
.A(n_5655),
.Y(n_6028)
);

AND2x4_ASAP7_75t_L g6029 ( 
.A(n_5412),
.B(n_4862),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5415),
.Y(n_6030)
);

AND2x2_ASAP7_75t_L g6031 ( 
.A(n_5705),
.B(n_4448),
.Y(n_6031)
);

AOI22xp5_ASAP7_75t_L g6032 ( 
.A1(n_5724),
.A2(n_5645),
.B1(n_5644),
.B2(n_5694),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5670),
.Y(n_6033)
);

OAI22xp5_ASAP7_75t_L g6034 ( 
.A1(n_5324),
.A2(n_4727),
.B1(n_4733),
.B2(n_4718),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5775),
.B(n_4387),
.Y(n_6035)
);

INVx5_ASAP7_75t_L g6036 ( 
.A(n_5678),
.Y(n_6036)
);

AND2x2_ASAP7_75t_L g6037 ( 
.A(n_5383),
.B(n_4474),
.Y(n_6037)
);

HB1xp67_ASAP7_75t_L g6038 ( 
.A(n_5473),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5491),
.B(n_4474),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5672),
.Y(n_6040)
);

BUFx6f_ASAP7_75t_L g6041 ( 
.A(n_5386),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5675),
.Y(n_6042)
);

AOI22xp5_ASAP7_75t_L g6043 ( 
.A1(n_5699),
.A2(n_4597),
.B1(n_4697),
.B2(n_4590),
.Y(n_6043)
);

BUFx2_ASAP7_75t_L g6044 ( 
.A(n_5710),
.Y(n_6044)
);

INVx2_ASAP7_75t_L g6045 ( 
.A(n_5416),
.Y(n_6045)
);

INVx3_ASAP7_75t_L g6046 ( 
.A(n_5388),
.Y(n_6046)
);

OA21x2_ASAP7_75t_L g6047 ( 
.A1(n_5776),
.A2(n_3517),
.B(n_3511),
.Y(n_6047)
);

NOR2xp33_ASAP7_75t_L g6048 ( 
.A(n_5717),
.B(n_4775),
.Y(n_6048)
);

BUFx6f_ASAP7_75t_L g6049 ( 
.A(n_5391),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5676),
.Y(n_6050)
);

BUFx6f_ASAP7_75t_L g6051 ( 
.A(n_5392),
.Y(n_6051)
);

BUFx2_ASAP7_75t_L g6052 ( 
.A(n_5715),
.Y(n_6052)
);

INVx2_ASAP7_75t_SL g6053 ( 
.A(n_5591),
.Y(n_6053)
);

INVx2_ASAP7_75t_L g6054 ( 
.A(n_5417),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5677),
.Y(n_6055)
);

XOR2xp5_ASAP7_75t_L g6056 ( 
.A(n_5311),
.B(n_4168),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5679),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5419),
.Y(n_6058)
);

BUFx6f_ASAP7_75t_L g6059 ( 
.A(n_5393),
.Y(n_6059)
);

BUFx6f_ASAP7_75t_L g6060 ( 
.A(n_5394),
.Y(n_6060)
);

BUFx6f_ASAP7_75t_L g6061 ( 
.A(n_5395),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5680),
.Y(n_6062)
);

OAI22xp5_ASAP7_75t_L g6063 ( 
.A1(n_5539),
.A2(n_4827),
.B1(n_4834),
.B2(n_4818),
.Y(n_6063)
);

AND2x4_ASAP7_75t_L g6064 ( 
.A(n_5422),
.B(n_3496),
.Y(n_6064)
);

AND2x6_ASAP7_75t_L g6065 ( 
.A(n_5755),
.B(n_4749),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5363),
.B(n_4483),
.Y(n_6066)
);

INVx3_ASAP7_75t_L g6067 ( 
.A(n_5398),
.Y(n_6067)
);

OAI21x1_ASAP7_75t_L g6068 ( 
.A1(n_5777),
.A2(n_3714),
.B(n_3667),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5684),
.Y(n_6069)
);

AND2x6_ASAP7_75t_L g6070 ( 
.A(n_5756),
.B(n_4768),
.Y(n_6070)
);

AND2x2_ASAP7_75t_L g6071 ( 
.A(n_5370),
.B(n_4483),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5685),
.Y(n_6072)
);

BUFx2_ASAP7_75t_L g6073 ( 
.A(n_5721),
.Y(n_6073)
);

BUFx6f_ASAP7_75t_L g6074 ( 
.A(n_5402),
.Y(n_6074)
);

AOI22xp5_ASAP7_75t_L g6075 ( 
.A1(n_5611),
.A2(n_4786),
.B1(n_4789),
.B2(n_4784),
.Y(n_6075)
);

INVx2_ASAP7_75t_L g6076 ( 
.A(n_5420),
.Y(n_6076)
);

BUFx6f_ASAP7_75t_L g6077 ( 
.A(n_5405),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5693),
.Y(n_6078)
);

INVx3_ASAP7_75t_L g6079 ( 
.A(n_5406),
.Y(n_6079)
);

CKINVDCx5p33_ASAP7_75t_R g6080 ( 
.A(n_5379),
.Y(n_6080)
);

BUFx6f_ASAP7_75t_L g6081 ( 
.A(n_5695),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5456),
.B(n_5786),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5696),
.Y(n_6083)
);

BUFx3_ASAP7_75t_L g6084 ( 
.A(n_5725),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5697),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5778),
.Y(n_6086)
);

NOR2x1_ASAP7_75t_L g6087 ( 
.A(n_5780),
.B(n_3843),
.Y(n_6087)
);

BUFx6f_ASAP7_75t_L g6088 ( 
.A(n_5708),
.Y(n_6088)
);

NOR2xp33_ASAP7_75t_L g6089 ( 
.A(n_5380),
.B(n_4843),
.Y(n_6089)
);

AND2x4_ASAP7_75t_L g6090 ( 
.A(n_5523),
.B(n_3717),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5783),
.Y(n_6091)
);

AND2x2_ASAP7_75t_SL g6092 ( 
.A(n_5440),
.B(n_5520),
.Y(n_6092)
);

BUFx6f_ASAP7_75t_L g6093 ( 
.A(n_5709),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5784),
.Y(n_6094)
);

BUFx6f_ASAP7_75t_L g6095 ( 
.A(n_5712),
.Y(n_6095)
);

AND2x4_ASAP7_75t_L g6096 ( 
.A(n_5524),
.B(n_4457),
.Y(n_6096)
);

AND2x2_ASAP7_75t_L g6097 ( 
.A(n_5344),
.B(n_4791),
.Y(n_6097)
);

INVx2_ASAP7_75t_L g6098 ( 
.A(n_5421),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5423),
.Y(n_6099)
);

INVx2_ASAP7_75t_L g6100 ( 
.A(n_5424),
.Y(n_6100)
);

AND2x4_ASAP7_75t_L g6101 ( 
.A(n_5526),
.B(n_5787),
.Y(n_6101)
);

OAI22xp5_ASAP7_75t_SL g6102 ( 
.A1(n_5730),
.A2(n_4235),
.B1(n_4258),
.B2(n_4106),
.Y(n_6102)
);

CKINVDCx5p33_ASAP7_75t_R g6103 ( 
.A(n_5385),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5790),
.Y(n_6104)
);

INVx6_ASAP7_75t_L g6105 ( 
.A(n_5799),
.Y(n_6105)
);

OA21x2_ASAP7_75t_L g6106 ( 
.A1(n_5791),
.A2(n_3531),
.B(n_3523),
.Y(n_6106)
);

BUFx6f_ASAP7_75t_L g6107 ( 
.A(n_5713),
.Y(n_6107)
);

CKINVDCx16_ASAP7_75t_R g6108 ( 
.A(n_5328),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5793),
.Y(n_6109)
);

BUFx6f_ASAP7_75t_L g6110 ( 
.A(n_5718),
.Y(n_6110)
);

BUFx3_ASAP7_75t_L g6111 ( 
.A(n_5736),
.Y(n_6111)
);

BUFx2_ASAP7_75t_L g6112 ( 
.A(n_5742),
.Y(n_6112)
);

BUFx6f_ASAP7_75t_L g6113 ( 
.A(n_5719),
.Y(n_6113)
);

AOI22xp5_ASAP7_75t_L g6114 ( 
.A1(n_5625),
.A2(n_4831),
.B1(n_4857),
.B2(n_4796),
.Y(n_6114)
);

BUFx3_ASAP7_75t_L g6115 ( 
.A(n_5743),
.Y(n_6115)
);

INVx1_ASAP7_75t_SL g6116 ( 
.A(n_5329),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5431),
.Y(n_6117)
);

INVx6_ASAP7_75t_L g6118 ( 
.A(n_5397),
.Y(n_6118)
);

XNOR2xp5_ASAP7_75t_L g6119 ( 
.A(n_5335),
.B(n_4338),
.Y(n_6119)
);

AND2x2_ASAP7_75t_L g6120 ( 
.A(n_5792),
.B(n_3541),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5433),
.Y(n_6121)
);

INVx4_ASAP7_75t_L g6122 ( 
.A(n_5389),
.Y(n_6122)
);

AND2x2_ASAP7_75t_L g6123 ( 
.A(n_5797),
.B(n_3595),
.Y(n_6123)
);

INVx3_ASAP7_75t_L g6124 ( 
.A(n_5794),
.Y(n_6124)
);

BUFx6f_ASAP7_75t_L g6125 ( 
.A(n_5438),
.Y(n_6125)
);

INVx2_ASAP7_75t_L g6126 ( 
.A(n_5441),
.Y(n_6126)
);

AND2x2_ASAP7_75t_L g6127 ( 
.A(n_5649),
.B(n_3595),
.Y(n_6127)
);

INVxp67_ASAP7_75t_L g6128 ( 
.A(n_5757),
.Y(n_6128)
);

AND2x4_ASAP7_75t_L g6129 ( 
.A(n_5795),
.B(n_4822),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_5442),
.Y(n_6130)
);

CKINVDCx11_ASAP7_75t_R g6131 ( 
.A(n_5354),
.Y(n_6131)
);

AOI22xp5_ASAP7_75t_L g6132 ( 
.A1(n_5566),
.A2(n_3467),
.B1(n_3468),
.B2(n_3466),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5796),
.Y(n_6133)
);

BUFx6f_ASAP7_75t_L g6134 ( 
.A(n_5443),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_5444),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_5807),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5808),
.Y(n_6137)
);

NOR2xp33_ASAP7_75t_L g6138 ( 
.A(n_5400),
.B(n_3585),
.Y(n_6138)
);

AND2x4_ASAP7_75t_L g6139 ( 
.A(n_5811),
.B(n_3620),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5812),
.Y(n_6140)
);

BUFx6f_ASAP7_75t_L g6141 ( 
.A(n_5447),
.Y(n_6141)
);

INVx2_ASAP7_75t_L g6142 ( 
.A(n_5448),
.Y(n_6142)
);

NAND2xp5_ASAP7_75t_L g6143 ( 
.A(n_5814),
.B(n_4472),
.Y(n_6143)
);

BUFx6f_ASAP7_75t_L g6144 ( 
.A(n_5450),
.Y(n_6144)
);

BUFx2_ASAP7_75t_L g6145 ( 
.A(n_5744),
.Y(n_6145)
);

INVx2_ASAP7_75t_L g6146 ( 
.A(n_5453),
.Y(n_6146)
);

BUFx6f_ASAP7_75t_L g6147 ( 
.A(n_5457),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5529),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5534),
.Y(n_6149)
);

OAI21x1_ASAP7_75t_L g6150 ( 
.A1(n_5535),
.A2(n_5538),
.B(n_5537),
.Y(n_6150)
);

NOR2xp33_ASAP7_75t_L g6151 ( 
.A(n_5401),
.B(n_3676),
.Y(n_6151)
);

BUFx6f_ASAP7_75t_L g6152 ( 
.A(n_5459),
.Y(n_6152)
);

INVx5_ASAP7_75t_L g6153 ( 
.A(n_5781),
.Y(n_6153)
);

NOR2xp33_ASAP7_75t_L g6154 ( 
.A(n_5425),
.B(n_3706),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_5460),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5540),
.Y(n_6156)
);

BUFx12f_ASAP7_75t_L g6157 ( 
.A(n_5429),
.Y(n_6157)
);

CKINVDCx5p33_ASAP7_75t_R g6158 ( 
.A(n_5432),
.Y(n_6158)
);

AND2x4_ASAP7_75t_L g6159 ( 
.A(n_5543),
.B(n_3787),
.Y(n_6159)
);

AND2x2_ASAP7_75t_L g6160 ( 
.A(n_5734),
.B(n_3610),
.Y(n_6160)
);

INVx1_ASAP7_75t_L g6161 ( 
.A(n_5544),
.Y(n_6161)
);

OA21x2_ASAP7_75t_L g6162 ( 
.A1(n_5545),
.A2(n_3534),
.B(n_3532),
.Y(n_6162)
);

NOR2xp33_ASAP7_75t_L g6163 ( 
.A(n_5446),
.B(n_3846),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5548),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_5552),
.B(n_3891),
.Y(n_6165)
);

AND2x4_ASAP7_75t_L g6166 ( 
.A(n_5553),
.B(n_3963),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_5571),
.B(n_3610),
.Y(n_6167)
);

BUFx6f_ASAP7_75t_L g6168 ( 
.A(n_5469),
.Y(n_6168)
);

BUFx6f_ASAP7_75t_L g6169 ( 
.A(n_5471),
.Y(n_6169)
);

OA21x2_ASAP7_75t_L g6170 ( 
.A1(n_5554),
.A2(n_3536),
.B(n_3535),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_5472),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5556),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5557),
.Y(n_6173)
);

BUFx12f_ASAP7_75t_L g6174 ( 
.A(n_5455),
.Y(n_6174)
);

INVx3_ASAP7_75t_L g6175 ( 
.A(n_5559),
.Y(n_6175)
);

NOR2xp33_ASAP7_75t_L g6176 ( 
.A(n_5461),
.B(n_4044),
.Y(n_6176)
);

NOR2xp33_ASAP7_75t_L g6177 ( 
.A(n_5463),
.B(n_4111),
.Y(n_6177)
);

OA21x2_ASAP7_75t_L g6178 ( 
.A1(n_5560),
.A2(n_3558),
.B(n_3544),
.Y(n_6178)
);

OR2x6_ASAP7_75t_L g6179 ( 
.A(n_5315),
.B(n_4654),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_5561),
.Y(n_6180)
);

BUFx2_ASAP7_75t_L g6181 ( 
.A(n_5390),
.Y(n_6181)
);

AOI22xp5_ASAP7_75t_L g6182 ( 
.A1(n_5466),
.A2(n_3472),
.B1(n_3473),
.B2(n_3469),
.Y(n_6182)
);

BUFx12f_ASAP7_75t_L g6183 ( 
.A(n_5467),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5565),
.Y(n_6184)
);

INVx2_ASAP7_75t_L g6185 ( 
.A(n_5474),
.Y(n_6185)
);

AND2x2_ASAP7_75t_L g6186 ( 
.A(n_5468),
.B(n_3681),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_5569),
.B(n_5572),
.Y(n_6187)
);

BUFx3_ASAP7_75t_L g6188 ( 
.A(n_5575),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5576),
.Y(n_6189)
);

INVx2_ASAP7_75t_L g6190 ( 
.A(n_5479),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5480),
.Y(n_6191)
);

INVx2_ASAP7_75t_L g6192 ( 
.A(n_5481),
.Y(n_6192)
);

INVx6_ASAP7_75t_L g6193 ( 
.A(n_5782),
.Y(n_6193)
);

BUFx6f_ASAP7_75t_L g6194 ( 
.A(n_5485),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5486),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_L g6196 ( 
.A(n_5488),
.B(n_4472),
.Y(n_6196)
);

INVx2_ASAP7_75t_L g6197 ( 
.A(n_5489),
.Y(n_6197)
);

NOR2x1_ASAP7_75t_L g6198 ( 
.A(n_5493),
.B(n_4779),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_5494),
.Y(n_6199)
);

OA21x2_ASAP7_75t_L g6200 ( 
.A1(n_5495),
.A2(n_5497),
.B(n_5496),
.Y(n_6200)
);

INVx3_ASAP7_75t_L g6201 ( 
.A(n_5498),
.Y(n_6201)
);

INVx5_ASAP7_75t_L g6202 ( 
.A(n_5310),
.Y(n_6202)
);

AOI22xp5_ASAP7_75t_L g6203 ( 
.A1(n_5470),
.A2(n_3478),
.B1(n_3484),
.B2(n_3474),
.Y(n_6203)
);

OA21x2_ASAP7_75t_L g6204 ( 
.A1(n_5499),
.A2(n_3562),
.B(n_3560),
.Y(n_6204)
);

BUFx12f_ASAP7_75t_L g6205 ( 
.A(n_5477),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5500),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_5501),
.Y(n_6207)
);

AND2x2_ASAP7_75t_L g6208 ( 
.A(n_5478),
.B(n_3681),
.Y(n_6208)
);

INVx2_ASAP7_75t_L g6209 ( 
.A(n_5502),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_5504),
.Y(n_6210)
);

NAND2xp5_ASAP7_75t_L g6211 ( 
.A(n_5505),
.B(n_4472),
.Y(n_6211)
);

AND2x2_ASAP7_75t_L g6212 ( 
.A(n_5482),
.B(n_5487),
.Y(n_6212)
);

BUFx6f_ASAP7_75t_L g6213 ( 
.A(n_5508),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_5512),
.Y(n_6214)
);

CKINVDCx16_ASAP7_75t_R g6215 ( 
.A(n_5396),
.Y(n_6215)
);

INVx3_ASAP7_75t_L g6216 ( 
.A(n_5515),
.Y(n_6216)
);

INVx3_ASAP7_75t_L g6217 ( 
.A(n_5516),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_5503),
.Y(n_6218)
);

INVx2_ASAP7_75t_L g6219 ( 
.A(n_5517),
.Y(n_6219)
);

BUFx6f_ASAP7_75t_L g6220 ( 
.A(n_5521),
.Y(n_6220)
);

INVx3_ASAP7_75t_L g6221 ( 
.A(n_5506),
.Y(n_6221)
);

CKINVDCx5p33_ASAP7_75t_R g6222 ( 
.A(n_5509),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5321),
.Y(n_6223)
);

BUFx3_ASAP7_75t_L g6224 ( 
.A(n_5614),
.Y(n_6224)
);

INVx3_ASAP7_75t_L g6225 ( 
.A(n_5513),
.Y(n_6225)
);

INVx6_ASAP7_75t_L g6226 ( 
.A(n_5399),
.Y(n_6226)
);

BUFx6f_ASAP7_75t_L g6227 ( 
.A(n_5519),
.Y(n_6227)
);

AND2x6_ASAP7_75t_L g6228 ( 
.A(n_5594),
.B(n_4621),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_5525),
.Y(n_6229)
);

INVxp67_ASAP7_75t_L g6230 ( 
.A(n_5408),
.Y(n_6230)
);

AND2x4_ASAP7_75t_L g6231 ( 
.A(n_5426),
.B(n_4141),
.Y(n_6231)
);

OAI22x1_ASAP7_75t_R g6232 ( 
.A1(n_5409),
.A2(n_4559),
.B1(n_4604),
.B2(n_4551),
.Y(n_6232)
);

CKINVDCx20_ASAP7_75t_R g6233 ( 
.A(n_5414),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_5518),
.Y(n_6234)
);

OAI22x1_ASAP7_75t_SL g6235 ( 
.A1(n_5418),
.A2(n_4795),
.B1(n_4799),
.B2(n_4640),
.Y(n_6235)
);

NAND2xp5_ASAP7_75t_L g6236 ( 
.A(n_5531),
.B(n_5533),
.Y(n_6236)
);

BUFx6f_ASAP7_75t_L g6237 ( 
.A(n_5536),
.Y(n_6237)
);

INVx3_ASAP7_75t_L g6238 ( 
.A(n_5542),
.Y(n_6238)
);

INVx2_ASAP7_75t_L g6239 ( 
.A(n_5546),
.Y(n_6239)
);

HB1xp67_ASAP7_75t_L g6240 ( 
.A(n_5567),
.Y(n_6240)
);

NOR2xp33_ASAP7_75t_L g6241 ( 
.A(n_5547),
.B(n_4157),
.Y(n_6241)
);

AND2x2_ASAP7_75t_L g6242 ( 
.A(n_5549),
.B(n_3693),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5550),
.Y(n_6243)
);

OA21x2_ASAP7_75t_L g6244 ( 
.A1(n_5555),
.A2(n_3577),
.B(n_3566),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5558),
.Y(n_6245)
);

BUFx6f_ASAP7_75t_L g6246 ( 
.A(n_5562),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_5568),
.Y(n_6247)
);

HB1xp67_ASAP7_75t_L g6248 ( 
.A(n_5570),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_5582),
.B(n_4621),
.Y(n_6249)
);

AND2x2_ASAP7_75t_L g6250 ( 
.A(n_5586),
.B(n_3693),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5595),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5598),
.Y(n_6252)
);

BUFx6f_ASAP7_75t_L g6253 ( 
.A(n_5603),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_5615),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_5617),
.Y(n_6255)
);

NAND2xp5_ASAP7_75t_L g6256 ( 
.A(n_5622),
.B(n_4621),
.Y(n_6256)
);

INVx2_ASAP7_75t_L g6257 ( 
.A(n_5623),
.Y(n_6257)
);

INVx2_ASAP7_75t_L g6258 ( 
.A(n_5624),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_5641),
.B(n_4651),
.Y(n_6259)
);

INVxp33_ASAP7_75t_SL g6260 ( 
.A(n_5652),
.Y(n_6260)
);

BUFx6f_ASAP7_75t_L g6261 ( 
.A(n_5660),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_5663),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_5664),
.Y(n_6263)
);

INVx2_ASAP7_75t_L g6264 ( 
.A(n_5673),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5674),
.Y(n_6265)
);

AND2x4_ASAP7_75t_L g6266 ( 
.A(n_5683),
.B(n_4316),
.Y(n_6266)
);

CKINVDCx11_ASAP7_75t_R g6267 ( 
.A(n_5437),
.Y(n_6267)
);

INVx2_ASAP7_75t_L g6268 ( 
.A(n_5686),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5688),
.Y(n_6269)
);

AOI22xp5_ASAP7_75t_L g6270 ( 
.A1(n_5692),
.A2(n_3488),
.B1(n_3489),
.B2(n_3485),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5703),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_5727),
.Y(n_6272)
);

HB1xp67_ASAP7_75t_L g6273 ( 
.A(n_5737),
.Y(n_6273)
);

BUFx6f_ASAP7_75t_L g6274 ( 
.A(n_5739),
.Y(n_6274)
);

AND2x4_ASAP7_75t_L g6275 ( 
.A(n_5740),
.B(n_4603),
.Y(n_6275)
);

INVx1_ASAP7_75t_L g6276 ( 
.A(n_5748),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_5750),
.Y(n_6277)
);

AND2x6_ASAP7_75t_L g6278 ( 
.A(n_5602),
.B(n_4651),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_5751),
.Y(n_6279)
);

BUFx3_ASAP7_75t_L g6280 ( 
.A(n_5439),
.Y(n_6280)
);

CKINVDCx5p33_ASAP7_75t_R g6281 ( 
.A(n_5313),
.Y(n_6281)
);

AND2x6_ASAP7_75t_L g6282 ( 
.A(n_5616),
.B(n_4651),
.Y(n_6282)
);

INVx2_ASAP7_75t_L g6283 ( 
.A(n_5330),
.Y(n_6283)
);

INVx4_ASAP7_75t_L g6284 ( 
.A(n_5331),
.Y(n_6284)
);

AND2x4_ASAP7_75t_L g6285 ( 
.A(n_5445),
.B(n_4774),
.Y(n_6285)
);

INVx3_ASAP7_75t_L g6286 ( 
.A(n_5332),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_5779),
.B(n_3744),
.Y(n_6287)
);

INVx5_ASAP7_75t_L g6288 ( 
.A(n_5789),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_5434),
.Y(n_6289)
);

AND2x4_ASAP7_75t_L g6290 ( 
.A(n_5449),
.B(n_3586),
.Y(n_6290)
);

BUFx6f_ASAP7_75t_L g6291 ( 
.A(n_5800),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_5454),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_5802),
.Y(n_6293)
);

AND2x2_ASAP7_75t_L g6294 ( 
.A(n_5803),
.B(n_3744),
.Y(n_6294)
);

NAND2xp5_ASAP7_75t_L g6295 ( 
.A(n_5530),
.B(n_4712),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_5805),
.Y(n_6296)
);

OAI21x1_ASAP7_75t_L g6297 ( 
.A1(n_5806),
.A2(n_3775),
.B(n_3737),
.Y(n_6297)
);

INVx2_ASAP7_75t_L g6298 ( 
.A(n_5810),
.Y(n_6298)
);

AND2x4_ASAP7_75t_L g6299 ( 
.A(n_5452),
.B(n_3588),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5813),
.Y(n_6300)
);

INVxp67_ASAP7_75t_L g6301 ( 
.A(n_5815),
.Y(n_6301)
);

INVx2_ASAP7_75t_L g6302 ( 
.A(n_5458),
.Y(n_6302)
);

BUFx6f_ASAP7_75t_L g6303 ( 
.A(n_5636),
.Y(n_6303)
);

BUFx6f_ASAP7_75t_L g6304 ( 
.A(n_5476),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5483),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_5484),
.Y(n_6306)
);

AND2x6_ASAP7_75t_L g6307 ( 
.A(n_5490),
.B(n_4712),
.Y(n_6307)
);

INVx3_ASAP7_75t_L g6308 ( 
.A(n_5507),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5510),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_5809),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_5527),
.Y(n_6311)
);

NAND2xp5_ASAP7_75t_L g6312 ( 
.A(n_5528),
.B(n_4712),
.Y(n_6312)
);

CKINVDCx20_ASAP7_75t_R g6313 ( 
.A(n_5551),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_5801),
.Y(n_6314)
);

NOR2xp33_ASAP7_75t_L g6315 ( 
.A(n_5573),
.B(n_3491),
.Y(n_6315)
);

INVx3_ASAP7_75t_L g6316 ( 
.A(n_5593),
.Y(n_6316)
);

CKINVDCx5p33_ASAP7_75t_R g6317 ( 
.A(n_5785),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_5788),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_5767),
.B(n_3757),
.Y(n_6319)
);

NAND2xp5_ASAP7_75t_L g6320 ( 
.A(n_5628),
.B(n_4737),
.Y(n_6320)
);

NAND2xp5_ASAP7_75t_L g6321 ( 
.A(n_5628),
.B(n_4737),
.Y(n_6321)
);

BUFx6f_ASAP7_75t_L g6322 ( 
.A(n_5403),
.Y(n_6322)
);

NAND2xp5_ASAP7_75t_L g6323 ( 
.A(n_5628),
.B(n_4737),
.Y(n_6323)
);

OAI22xp5_ASAP7_75t_SL g6324 ( 
.A1(n_5762),
.A2(n_4823),
.B1(n_4234),
.B2(n_4268),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5631),
.Y(n_6325)
);

INVx4_ASAP7_75t_L g6326 ( 
.A(n_5340),
.Y(n_6326)
);

INVx5_ASAP7_75t_L g6327 ( 
.A(n_5343),
.Y(n_6327)
);

AND2x2_ASAP7_75t_L g6328 ( 
.A(n_5767),
.B(n_3757),
.Y(n_6328)
);

BUFx3_ASAP7_75t_L g6329 ( 
.A(n_5387),
.Y(n_6329)
);

CKINVDCx6p67_ASAP7_75t_R g6330 ( 
.A(n_5341),
.Y(n_6330)
);

AND2x4_ASAP7_75t_L g6331 ( 
.A(n_5387),
.B(n_3589),
.Y(n_6331)
);

AOI22xp5_ASAP7_75t_L g6332 ( 
.A1(n_5349),
.A2(n_3495),
.B1(n_3499),
.B2(n_3494),
.Y(n_6332)
);

CKINVDCx5p33_ASAP7_75t_R g6333 ( 
.A(n_5340),
.Y(n_6333)
);

INVx3_ASAP7_75t_L g6334 ( 
.A(n_5387),
.Y(n_6334)
);

INVx2_ASAP7_75t_L g6335 ( 
.A(n_5404),
.Y(n_6335)
);

HB1xp67_ASAP7_75t_L g6336 ( 
.A(n_5326),
.Y(n_6336)
);

NAND2xp5_ASAP7_75t_SL g6337 ( 
.A(n_5767),
.B(n_4765),
.Y(n_6337)
);

HB1xp67_ASAP7_75t_L g6338 ( 
.A(n_5326),
.Y(n_6338)
);

AND2x6_ASAP7_75t_L g6339 ( 
.A(n_5732),
.B(n_4765),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_5631),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_5631),
.Y(n_6341)
);

OA21x2_ASAP7_75t_L g6342 ( 
.A1(n_5308),
.A2(n_3623),
.B(n_3598),
.Y(n_6342)
);

INVx5_ASAP7_75t_L g6343 ( 
.A(n_5343),
.Y(n_6343)
);

AND2x4_ASAP7_75t_L g6344 ( 
.A(n_5387),
.B(n_3624),
.Y(n_6344)
);

HB1xp67_ASAP7_75t_L g6345 ( 
.A(n_5326),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_5628),
.B(n_4765),
.Y(n_6346)
);

AND2x6_ASAP7_75t_L g6347 ( 
.A(n_5732),
.B(n_4807),
.Y(n_6347)
);

NAND2xp5_ASAP7_75t_L g6348 ( 
.A(n_5628),
.B(n_4807),
.Y(n_6348)
);

BUFx6f_ASAP7_75t_L g6349 ( 
.A(n_5403),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_5404),
.Y(n_6350)
);

OAI21x1_ASAP7_75t_L g6351 ( 
.A1(n_5407),
.A2(n_3814),
.B(n_3811),
.Y(n_6351)
);

OAI22xp5_ASAP7_75t_L g6352 ( 
.A1(n_5619),
.A2(n_3506),
.B1(n_3509),
.B2(n_3501),
.Y(n_6352)
);

AND2x2_ASAP7_75t_L g6353 ( 
.A(n_5767),
.B(n_3810),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_5628),
.B(n_4807),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5631),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_5767),
.B(n_3810),
.Y(n_6356)
);

NAND2xp5_ASAP7_75t_L g6357 ( 
.A(n_5628),
.B(n_4829),
.Y(n_6357)
);

INVx4_ASAP7_75t_L g6358 ( 
.A(n_5340),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_5628),
.B(n_4829),
.Y(n_6359)
);

NAND2xp5_ASAP7_75t_L g6360 ( 
.A(n_5628),
.B(n_4829),
.Y(n_6360)
);

BUFx6f_ASAP7_75t_L g6361 ( 
.A(n_5403),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5631),
.Y(n_6362)
);

INVx2_ASAP7_75t_L g6363 ( 
.A(n_5404),
.Y(n_6363)
);

BUFx12f_ASAP7_75t_L g6364 ( 
.A(n_5759),
.Y(n_6364)
);

INVx5_ASAP7_75t_L g6365 ( 
.A(n_5343),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_5326),
.Y(n_6366)
);

HB1xp67_ASAP7_75t_L g6367 ( 
.A(n_5326),
.Y(n_6367)
);

INVx2_ASAP7_75t_SL g6368 ( 
.A(n_5760),
.Y(n_6368)
);

OAI21x1_ASAP7_75t_L g6369 ( 
.A1(n_5407),
.A2(n_3933),
.B(n_3902),
.Y(n_6369)
);

INVx3_ASAP7_75t_L g6370 ( 
.A(n_5387),
.Y(n_6370)
);

BUFx2_ASAP7_75t_L g6371 ( 
.A(n_5762),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_5628),
.B(n_3976),
.Y(n_6372)
);

AOI22xp5_ASAP7_75t_L g6373 ( 
.A1(n_5349),
.A2(n_3514),
.B1(n_3518),
.B2(n_3513),
.Y(n_6373)
);

AND2x4_ASAP7_75t_L g6374 ( 
.A(n_5387),
.B(n_3635),
.Y(n_6374)
);

BUFx2_ASAP7_75t_L g6375 ( 
.A(n_5762),
.Y(n_6375)
);

HB1xp67_ASAP7_75t_L g6376 ( 
.A(n_5326),
.Y(n_6376)
);

HB1xp67_ASAP7_75t_L g6377 ( 
.A(n_5326),
.Y(n_6377)
);

BUFx6f_ASAP7_75t_L g6378 ( 
.A(n_5403),
.Y(n_6378)
);

NOR2x1_ASAP7_75t_L g6379 ( 
.A(n_5732),
.B(n_3636),
.Y(n_6379)
);

OAI21x1_ASAP7_75t_L g6380 ( 
.A1(n_5407),
.A2(n_4027),
.B(n_4011),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_5631),
.Y(n_6381)
);

BUFx2_ASAP7_75t_L g6382 ( 
.A(n_5762),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_5404),
.Y(n_6383)
);

AOI22xp5_ASAP7_75t_L g6384 ( 
.A1(n_5349),
.A2(n_3520),
.B1(n_3521),
.B2(n_3519),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_5631),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_5628),
.B(n_4160),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_5628),
.B(n_4238),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5631),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_5404),
.Y(n_6389)
);

INVx6_ASAP7_75t_L g6390 ( 
.A(n_5387),
.Y(n_6390)
);

AND2x2_ASAP7_75t_L g6391 ( 
.A(n_5767),
.B(n_3918),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_5767),
.B(n_3918),
.Y(n_6392)
);

BUFx2_ASAP7_75t_L g6393 ( 
.A(n_5762),
.Y(n_6393)
);

BUFx6f_ASAP7_75t_L g6394 ( 
.A(n_5403),
.Y(n_6394)
);

INVx4_ASAP7_75t_L g6395 ( 
.A(n_5340),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6200),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_5927),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_5835),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_5839),
.Y(n_6399)
);

NOR2xp33_ASAP7_75t_L g6400 ( 
.A(n_5840),
.B(n_3522),
.Y(n_6400)
);

NAND2xp5_ASAP7_75t_L g6401 ( 
.A(n_6082),
.B(n_3526),
.Y(n_6401)
);

INVx2_ASAP7_75t_L g6402 ( 
.A(n_5836),
.Y(n_6402)
);

NAND2xp5_ASAP7_75t_L g6403 ( 
.A(n_6086),
.B(n_3527),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_6091),
.B(n_3528),
.Y(n_6404)
);

BUFx3_ASAP7_75t_L g6405 ( 
.A(n_6390),
.Y(n_6405)
);

INVxp67_ASAP7_75t_L g6406 ( 
.A(n_5838),
.Y(n_6406)
);

AND2x4_ASAP7_75t_L g6407 ( 
.A(n_5818),
.B(n_3637),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_6094),
.B(n_3533),
.Y(n_6408)
);

NAND2xp5_ASAP7_75t_SL g6409 ( 
.A(n_5932),
.B(n_3537),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5843),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_5866),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_L g6412 ( 
.A(n_6104),
.B(n_3543),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_5894),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_5855),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5857),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5864),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_5871),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_5902),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_6109),
.B(n_3545),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5872),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5874),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_5875),
.Y(n_6422)
);

BUFx6f_ASAP7_75t_L g6423 ( 
.A(n_6303),
.Y(n_6423)
);

XNOR2xp5_ASAP7_75t_L g6424 ( 
.A(n_6056),
.B(n_4211),
.Y(n_6424)
);

OA21x2_ASAP7_75t_L g6425 ( 
.A1(n_6150),
.A2(n_3644),
.B(n_3643),
.Y(n_6425)
);

INVx3_ASAP7_75t_L g6426 ( 
.A(n_5916),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_5878),
.Y(n_6427)
);

INVx3_ASAP7_75t_L g6428 ( 
.A(n_5923),
.Y(n_6428)
);

INVxp67_ASAP7_75t_L g6429 ( 
.A(n_5863),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_5881),
.Y(n_6430)
);

AND2x2_ASAP7_75t_L g6431 ( 
.A(n_6336),
.B(n_3923),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_5885),
.Y(n_6432)
);

AND2x2_ASAP7_75t_L g6433 ( 
.A(n_6338),
.B(n_6345),
.Y(n_6433)
);

INVx2_ASAP7_75t_L g6434 ( 
.A(n_5906),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_5915),
.Y(n_6435)
);

INVx1_ASAP7_75t_SL g6436 ( 
.A(n_6366),
.Y(n_6436)
);

INVx2_ASAP7_75t_L g6437 ( 
.A(n_5971),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_5973),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_5886),
.Y(n_6439)
);

BUFx6f_ASAP7_75t_L g6440 ( 
.A(n_6394),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_5978),
.Y(n_6441)
);

INVx2_ASAP7_75t_L g6442 ( 
.A(n_5999),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5887),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_6133),
.B(n_6136),
.Y(n_6444)
);

NAND3xp33_ASAP7_75t_L g6445 ( 
.A(n_5830),
.B(n_3547),
.C(n_3546),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_5895),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5896),
.Y(n_6447)
);

INVx3_ASAP7_75t_L g6448 ( 
.A(n_5924),
.Y(n_6448)
);

INVx2_ASAP7_75t_L g6449 ( 
.A(n_6003),
.Y(n_6449)
);

NOR2xp33_ASAP7_75t_L g6450 ( 
.A(n_5979),
.B(n_3548),
.Y(n_6450)
);

OAI22xp5_ASAP7_75t_L g6451 ( 
.A1(n_6032),
.A2(n_3551),
.B1(n_3552),
.B2(n_3550),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_5900),
.Y(n_6452)
);

INVx1_ASAP7_75t_SL g6453 ( 
.A(n_6367),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_5910),
.Y(n_6454)
);

BUFx6f_ASAP7_75t_L g6455 ( 
.A(n_5821),
.Y(n_6455)
);

OAI22xp5_ASAP7_75t_L g6456 ( 
.A1(n_5837),
.A2(n_3556),
.B1(n_3557),
.B2(n_3554),
.Y(n_6456)
);

INVx2_ASAP7_75t_L g6457 ( 
.A(n_5918),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_5917),
.Y(n_6458)
);

BUFx6f_ASAP7_75t_L g6459 ( 
.A(n_5827),
.Y(n_6459)
);

BUFx2_ASAP7_75t_L g6460 ( 
.A(n_6377),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_5936),
.Y(n_6461)
);

CKINVDCx5p33_ASAP7_75t_R g6462 ( 
.A(n_5825),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5919),
.Y(n_6463)
);

INVx2_ASAP7_75t_L g6464 ( 
.A(n_5941),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_5920),
.Y(n_6465)
);

BUFx2_ASAP7_75t_L g6466 ( 
.A(n_6376),
.Y(n_6466)
);

HB1xp67_ASAP7_75t_L g6467 ( 
.A(n_5856),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_5921),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_5926),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_5934),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_5945),
.Y(n_6471)
);

AND2x4_ASAP7_75t_L g6472 ( 
.A(n_5822),
.B(n_3645),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_5940),
.Y(n_6473)
);

OA21x2_ASAP7_75t_L g6474 ( 
.A1(n_6016),
.A2(n_3668),
.B(n_3658),
.Y(n_6474)
);

INVx2_ASAP7_75t_L g6475 ( 
.A(n_5946),
.Y(n_6475)
);

NAND2xp5_ASAP7_75t_L g6476 ( 
.A(n_6137),
.B(n_3559),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_5944),
.Y(n_6477)
);

INVx2_ASAP7_75t_L g6478 ( 
.A(n_5948),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_5947),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5949),
.Y(n_6480)
);

NAND2xp5_ASAP7_75t_L g6481 ( 
.A(n_6140),
.B(n_3565),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_5953),
.Y(n_6482)
);

INVx2_ASAP7_75t_L g6483 ( 
.A(n_5960),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_5954),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6148),
.B(n_3568),
.Y(n_6485)
);

HB1xp67_ASAP7_75t_L g6486 ( 
.A(n_5938),
.Y(n_6486)
);

HB1xp67_ASAP7_75t_L g6487 ( 
.A(n_6312),
.Y(n_6487)
);

INVx2_ASAP7_75t_SL g6488 ( 
.A(n_6031),
.Y(n_6488)
);

BUFx3_ASAP7_75t_L g6489 ( 
.A(n_6329),
.Y(n_6489)
);

INVx2_ASAP7_75t_L g6490 ( 
.A(n_5962),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_5965),
.Y(n_6491)
);

HB1xp67_ASAP7_75t_L g6492 ( 
.A(n_5841),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_5967),
.Y(n_6493)
);

INVx2_ASAP7_75t_L g6494 ( 
.A(n_5968),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_5981),
.Y(n_6495)
);

NAND2xp5_ASAP7_75t_SL g6496 ( 
.A(n_6319),
.B(n_3569),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_5986),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_5990),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_5995),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_6009),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6001),
.Y(n_6501)
);

INVx1_ASAP7_75t_L g6502 ( 
.A(n_6004),
.Y(n_6502)
);

BUFx6f_ASAP7_75t_L g6503 ( 
.A(n_5851),
.Y(n_6503)
);

INVx1_ASAP7_75t_SL g6504 ( 
.A(n_5860),
.Y(n_6504)
);

INVxp33_ASAP7_75t_SL g6505 ( 
.A(n_6119),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_6149),
.B(n_3570),
.Y(n_6506)
);

INVx3_ASAP7_75t_L g6507 ( 
.A(n_5933),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_6011),
.Y(n_6508)
);

INVx2_ASAP7_75t_L g6509 ( 
.A(n_6026),
.Y(n_6509)
);

INVx2_ASAP7_75t_L g6510 ( 
.A(n_6030),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6015),
.Y(n_6511)
);

OAI21x1_ASAP7_75t_L g6512 ( 
.A1(n_6068),
.A2(n_4329),
.B(n_4294),
.Y(n_6512)
);

BUFx6f_ASAP7_75t_L g6513 ( 
.A(n_5853),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_6019),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6033),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_6040),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_6042),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_6050),
.Y(n_6518)
);

BUFx6f_ASAP7_75t_L g6519 ( 
.A(n_5868),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6055),
.Y(n_6520)
);

INVx3_ASAP7_75t_L g6521 ( 
.A(n_5935),
.Y(n_6521)
);

AND2x2_ASAP7_75t_L g6522 ( 
.A(n_6328),
.B(n_3923),
.Y(n_6522)
);

INVx3_ASAP7_75t_L g6523 ( 
.A(n_5890),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6057),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6062),
.Y(n_6525)
);

HB1xp67_ASAP7_75t_L g6526 ( 
.A(n_6371),
.Y(n_6526)
);

OAI21x1_ASAP7_75t_L g6527 ( 
.A1(n_5832),
.A2(n_4360),
.B(n_4358),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_6069),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_6045),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_6054),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6072),
.Y(n_6531)
);

INVxp67_ASAP7_75t_L g6532 ( 
.A(n_6353),
.Y(n_6532)
);

AOI22xp5_ASAP7_75t_L g6533 ( 
.A1(n_5961),
.A2(n_4352),
.B1(n_4383),
.B2(n_4326),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_6078),
.Y(n_6534)
);

INVx1_ASAP7_75t_L g6535 ( 
.A(n_6083),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6085),
.Y(n_6536)
);

HB1xp67_ASAP7_75t_L g6537 ( 
.A(n_6375),
.Y(n_6537)
);

BUFx3_ASAP7_75t_L g6538 ( 
.A(n_6226),
.Y(n_6538)
);

BUFx6f_ASAP7_75t_L g6539 ( 
.A(n_5870),
.Y(n_6539)
);

INVx2_ASAP7_75t_L g6540 ( 
.A(n_6058),
.Y(n_6540)
);

INVx2_ASAP7_75t_L g6541 ( 
.A(n_6076),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6191),
.Y(n_6542)
);

INVx1_ASAP7_75t_L g6543 ( 
.A(n_6195),
.Y(n_6543)
);

AND2x4_ASAP7_75t_L g6544 ( 
.A(n_5826),
.B(n_3692),
.Y(n_6544)
);

INVx1_ASAP7_75t_L g6545 ( 
.A(n_6206),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6214),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_6156),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_L g6548 ( 
.A(n_6161),
.B(n_3572),
.Y(n_6548)
);

INVx3_ASAP7_75t_L g6549 ( 
.A(n_5908),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6164),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6356),
.B(n_3975),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_6172),
.B(n_3575),
.Y(n_6552)
);

AND2x2_ASAP7_75t_L g6553 ( 
.A(n_6391),
.B(n_3975),
.Y(n_6553)
);

INVx2_ASAP7_75t_L g6554 ( 
.A(n_6098),
.Y(n_6554)
);

INVx3_ASAP7_75t_L g6555 ( 
.A(n_5905),
.Y(n_6555)
);

INVx2_ASAP7_75t_L g6556 ( 
.A(n_6099),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6173),
.Y(n_6557)
);

BUFx3_ASAP7_75t_L g6558 ( 
.A(n_6304),
.Y(n_6558)
);

OAI21x1_ASAP7_75t_L g6559 ( 
.A1(n_5847),
.A2(n_6369),
.B(n_6351),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_6100),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_6117),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_6121),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6180),
.Y(n_6563)
);

HB1xp67_ASAP7_75t_L g6564 ( 
.A(n_6382),
.Y(n_6564)
);

INVx2_ASAP7_75t_L g6565 ( 
.A(n_6126),
.Y(n_6565)
);

AND2x4_ASAP7_75t_L g6566 ( 
.A(n_6334),
.B(n_3697),
.Y(n_6566)
);

HB1xp67_ASAP7_75t_L g6567 ( 
.A(n_6393),
.Y(n_6567)
);

INVx1_ASAP7_75t_L g6568 ( 
.A(n_6184),
.Y(n_6568)
);

BUFx6f_ASAP7_75t_L g6569 ( 
.A(n_6322),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6189),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6101),
.Y(n_6571)
);

CKINVDCx5p33_ASAP7_75t_R g6572 ( 
.A(n_5848),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6130),
.Y(n_6573)
);

NAND2xp5_ASAP7_75t_SL g6574 ( 
.A(n_6392),
.B(n_3579),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6135),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6014),
.B(n_3992),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_6124),
.B(n_3581),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6142),
.Y(n_6578)
);

BUFx6f_ASAP7_75t_L g6579 ( 
.A(n_6349),
.Y(n_6579)
);

NAND2xp5_ASAP7_75t_L g6580 ( 
.A(n_6175),
.B(n_3582),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_6146),
.Y(n_6581)
);

INVx2_ASAP7_75t_L g6582 ( 
.A(n_6155),
.Y(n_6582)
);

INVx2_ASAP7_75t_L g6583 ( 
.A(n_6171),
.Y(n_6583)
);

HB1xp67_ASAP7_75t_L g6584 ( 
.A(n_5937),
.Y(n_6584)
);

BUFx6f_ASAP7_75t_L g6585 ( 
.A(n_6361),
.Y(n_6585)
);

BUFx2_ASAP7_75t_L g6586 ( 
.A(n_5963),
.Y(n_6586)
);

AND2x2_ASAP7_75t_L g6587 ( 
.A(n_6037),
.B(n_3992),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6185),
.Y(n_6588)
);

BUFx6f_ASAP7_75t_L g6589 ( 
.A(n_6378),
.Y(n_6589)
);

HB1xp67_ASAP7_75t_L g6590 ( 
.A(n_6290),
.Y(n_6590)
);

BUFx6f_ASAP7_75t_L g6591 ( 
.A(n_5859),
.Y(n_6591)
);

BUFx6f_ASAP7_75t_L g6592 ( 
.A(n_5912),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6190),
.Y(n_6593)
);

NAND2xp5_ASAP7_75t_L g6594 ( 
.A(n_6187),
.B(n_3584),
.Y(n_6594)
);

AND2x4_ASAP7_75t_L g6595 ( 
.A(n_6370),
.B(n_3703),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6192),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6197),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_SL g6598 ( 
.A(n_5873),
.B(n_6260),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6199),
.Y(n_6599)
);

HB1xp67_ASAP7_75t_L g6600 ( 
.A(n_6299),
.Y(n_6600)
);

INVx2_ASAP7_75t_L g6601 ( 
.A(n_6207),
.Y(n_6601)
);

INVxp67_ASAP7_75t_L g6602 ( 
.A(n_6066),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6209),
.Y(n_6603)
);

NAND2xp5_ASAP7_75t_SL g6604 ( 
.A(n_5883),
.B(n_5891),
.Y(n_6604)
);

HB1xp67_ASAP7_75t_L g6605 ( 
.A(n_6038),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6210),
.Y(n_6606)
);

AND2x2_ASAP7_75t_L g6607 ( 
.A(n_6071),
.B(n_3993),
.Y(n_6607)
);

HB1xp67_ASAP7_75t_L g6608 ( 
.A(n_6285),
.Y(n_6608)
);

BUFx3_ASAP7_75t_L g6609 ( 
.A(n_6233),
.Y(n_6609)
);

AND2x4_ASAP7_75t_L g6610 ( 
.A(n_6331),
.B(n_3707),
.Y(n_6610)
);

INVxp67_ASAP7_75t_L g6611 ( 
.A(n_6127),
.Y(n_6611)
);

INVx1_ASAP7_75t_SL g6612 ( 
.A(n_5987),
.Y(n_6612)
);

BUFx2_ASAP7_75t_L g6613 ( 
.A(n_6307),
.Y(n_6613)
);

NAND2xp5_ASAP7_75t_L g6614 ( 
.A(n_5831),
.B(n_3587),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_6219),
.Y(n_6615)
);

HB1xp67_ASAP7_75t_L g6616 ( 
.A(n_6244),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_5828),
.Y(n_6617)
);

BUFx6f_ASAP7_75t_L g6618 ( 
.A(n_6081),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_6335),
.Y(n_6619)
);

INVx3_ASAP7_75t_L g6620 ( 
.A(n_5842),
.Y(n_6620)
);

NAND2xp5_ASAP7_75t_L g6621 ( 
.A(n_5849),
.B(n_3596),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6350),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_6363),
.Y(n_6623)
);

BUFx6f_ASAP7_75t_L g6624 ( 
.A(n_6188),
.Y(n_6624)
);

OAI22xp5_ASAP7_75t_SL g6625 ( 
.A1(n_6102),
.A2(n_4406),
.B1(n_4412),
.B2(n_4404),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_5899),
.B(n_3993),
.Y(n_6626)
);

OA21x2_ASAP7_75t_L g6627 ( 
.A1(n_6380),
.A2(n_3723),
.B(n_3721),
.Y(n_6627)
);

INVx3_ASAP7_75t_L g6628 ( 
.A(n_5844),
.Y(n_6628)
);

INVx2_ASAP7_75t_L g6629 ( 
.A(n_6383),
.Y(n_6629)
);

INVx2_ASAP7_75t_L g6630 ( 
.A(n_6389),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_5824),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_5922),
.Y(n_6632)
);

AND2x2_ASAP7_75t_L g6633 ( 
.A(n_6368),
.B(n_4009),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_5854),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6320),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6321),
.Y(n_6636)
);

INVx3_ASAP7_75t_L g6637 ( 
.A(n_5845),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6323),
.Y(n_6638)
);

INVx2_ASAP7_75t_L g6639 ( 
.A(n_5928),
.Y(n_6639)
);

BUFx6f_ASAP7_75t_L g6640 ( 
.A(n_5867),
.Y(n_6640)
);

INVx1_ASAP7_75t_SL g6641 ( 
.A(n_5884),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6346),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6348),
.Y(n_6643)
);

BUFx6f_ASAP7_75t_L g6644 ( 
.A(n_5955),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_6354),
.Y(n_6645)
);

NAND2xp33_ASAP7_75t_L g6646 ( 
.A(n_6228),
.B(n_3599),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6357),
.Y(n_6647)
);

NAND2xp33_ASAP7_75t_SL g6648 ( 
.A(n_6186),
.B(n_4418),
.Y(n_6648)
);

OAI21x1_ASAP7_75t_L g6649 ( 
.A1(n_6297),
.A2(n_4464),
.B(n_4440),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_6359),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_5931),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6360),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_L g6653 ( 
.A(n_6007),
.B(n_3602),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5925),
.Y(n_6654)
);

BUFx6f_ASAP7_75t_L g6655 ( 
.A(n_5957),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_5956),
.Y(n_6656)
);

INVxp67_ASAP7_75t_L g6657 ( 
.A(n_6160),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6201),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_6216),
.Y(n_6659)
);

HB1xp67_ASAP7_75t_L g6660 ( 
.A(n_6231),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6217),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_SL g6662 ( 
.A(n_6138),
.B(n_3603),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_5939),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6204),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_5861),
.Y(n_6665)
);

INVxp67_ASAP7_75t_L g6666 ( 
.A(n_6167),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_5964),
.Y(n_6667)
);

INVx2_ASAP7_75t_L g6668 ( 
.A(n_5969),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_5980),
.Y(n_6669)
);

INVx1_ASAP7_75t_L g6670 ( 
.A(n_5984),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6017),
.Y(n_6671)
);

INVx3_ASAP7_75t_L g6672 ( 
.A(n_5846),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6047),
.Y(n_6673)
);

NAND2xp5_ASAP7_75t_SL g6674 ( 
.A(n_6151),
.B(n_3606),
.Y(n_6674)
);

BUFx6f_ASAP7_75t_L g6675 ( 
.A(n_5970),
.Y(n_6675)
);

NAND2xp33_ASAP7_75t_SL g6676 ( 
.A(n_6208),
.B(n_4453),
.Y(n_6676)
);

NAND2xp5_ASAP7_75t_L g6677 ( 
.A(n_6249),
.B(n_3611),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6106),
.Y(n_6678)
);

BUFx6f_ASAP7_75t_L g6679 ( 
.A(n_5982),
.Y(n_6679)
);

AOI22xp5_ASAP7_75t_L g6680 ( 
.A1(n_6379),
.A2(n_4488),
.B1(n_4491),
.B2(n_4465),
.Y(n_6680)
);

HB1xp67_ASAP7_75t_L g6681 ( 
.A(n_6179),
.Y(n_6681)
);

BUFx6f_ASAP7_75t_L g6682 ( 
.A(n_5988),
.Y(n_6682)
);

OAI22xp5_ASAP7_75t_SL g6683 ( 
.A1(n_6324),
.A2(n_4564),
.B1(n_4613),
.B2(n_4522),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6162),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_5985),
.Y(n_6685)
);

BUFx6f_ASAP7_75t_L g6686 ( 
.A(n_5989),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6170),
.Y(n_6687)
);

INVx2_ASAP7_75t_L g6688 ( 
.A(n_5993),
.Y(n_6688)
);

INVx2_ASAP7_75t_L g6689 ( 
.A(n_6046),
.Y(n_6689)
);

INVx3_ASAP7_75t_L g6690 ( 
.A(n_5850),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6178),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6342),
.Y(n_6692)
);

INVx1_ASAP7_75t_SL g6693 ( 
.A(n_5943),
.Y(n_6693)
);

INVx1_ASAP7_75t_L g6694 ( 
.A(n_5820),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_5829),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_5833),
.Y(n_6696)
);

INVx2_ASAP7_75t_L g6697 ( 
.A(n_6067),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6325),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6340),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6079),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6088),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_6341),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6355),
.Y(n_6703)
);

BUFx6f_ASAP7_75t_L g6704 ( 
.A(n_5996),
.Y(n_6704)
);

INVx3_ASAP7_75t_L g6705 ( 
.A(n_6093),
.Y(n_6705)
);

NAND3xp33_ASAP7_75t_L g6706 ( 
.A(n_6154),
.B(n_3615),
.C(n_3614),
.Y(n_6706)
);

NAND2xp5_ASAP7_75t_L g6707 ( 
.A(n_6256),
.B(n_3616),
.Y(n_6707)
);

BUFx6f_ASAP7_75t_L g6708 ( 
.A(n_5997),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6362),
.Y(n_6709)
);

OAI22xp5_ASAP7_75t_SL g6710 ( 
.A1(n_6000),
.A2(n_4668),
.B1(n_4673),
.B2(n_4638),
.Y(n_6710)
);

INVx2_ASAP7_75t_L g6711 ( 
.A(n_6095),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6381),
.Y(n_6712)
);

BUFx6f_ASAP7_75t_L g6713 ( 
.A(n_6002),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_6107),
.Y(n_6714)
);

BUFx3_ASAP7_75t_L g6715 ( 
.A(n_6313),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6385),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6025),
.B(n_4009),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6110),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6388),
.Y(n_6719)
);

NAND2xp5_ASAP7_75t_SL g6720 ( 
.A(n_6163),
.B(n_3618),
.Y(n_6720)
);

NAND2xp5_ASAP7_75t_L g6721 ( 
.A(n_6259),
.B(n_6176),
.Y(n_6721)
);

INVx1_ASAP7_75t_L g6722 ( 
.A(n_6372),
.Y(n_6722)
);

NAND2xp5_ASAP7_75t_SL g6723 ( 
.A(n_6177),
.B(n_3622),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6241),
.B(n_3625),
.Y(n_6724)
);

INVx2_ASAP7_75t_L g6725 ( 
.A(n_6113),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6386),
.Y(n_6726)
);

AND2x4_ASAP7_75t_L g6727 ( 
.A(n_6344),
.B(n_3726),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6387),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6196),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6211),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6035),
.Y(n_6731)
);

INVxp67_ASAP7_75t_L g6732 ( 
.A(n_6315),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6143),
.Y(n_6733)
);

NAND2xp5_ASAP7_75t_SL g6734 ( 
.A(n_6048),
.B(n_3627),
.Y(n_6734)
);

BUFx6f_ASAP7_75t_L g6735 ( 
.A(n_6005),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_6374),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6125),
.Y(n_6737)
);

INVx2_ASAP7_75t_L g6738 ( 
.A(n_6134),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_SL g6739 ( 
.A(n_6028),
.B(n_6266),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6141),
.Y(n_6740)
);

INVx3_ASAP7_75t_L g6741 ( 
.A(n_5889),
.Y(n_6741)
);

BUFx6f_ASAP7_75t_L g6742 ( 
.A(n_6012),
.Y(n_6742)
);

INVx2_ASAP7_75t_L g6743 ( 
.A(n_6144),
.Y(n_6743)
);

BUFx6f_ASAP7_75t_L g6744 ( 
.A(n_6022),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6242),
.B(n_4065),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6147),
.Y(n_6746)
);

BUFx6f_ASAP7_75t_L g6747 ( 
.A(n_6024),
.Y(n_6747)
);

NAND2xp5_ASAP7_75t_L g6748 ( 
.A(n_6064),
.B(n_3628),
.Y(n_6748)
);

INVx3_ASAP7_75t_L g6749 ( 
.A(n_5893),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6152),
.Y(n_6750)
);

BUFx6f_ASAP7_75t_L g6751 ( 
.A(n_6041),
.Y(n_6751)
);

NOR2xp33_ASAP7_75t_L g6752 ( 
.A(n_6089),
.B(n_3633),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6168),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6169),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6194),
.Y(n_6755)
);

NAND2xp5_ASAP7_75t_L g6756 ( 
.A(n_6295),
.B(n_3634),
.Y(n_6756)
);

BUFx6f_ASAP7_75t_L g6757 ( 
.A(n_6049),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6213),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_6220),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_5901),
.Y(n_6760)
);

BUFx2_ASAP7_75t_L g6761 ( 
.A(n_6307),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_6051),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6059),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6090),
.Y(n_6764)
);

INVx3_ASAP7_75t_L g6765 ( 
.A(n_6060),
.Y(n_6765)
);

INVx3_ASAP7_75t_L g6766 ( 
.A(n_6061),
.Y(n_6766)
);

BUFx6f_ASAP7_75t_L g6767 ( 
.A(n_6074),
.Y(n_6767)
);

AND2x2_ASAP7_75t_L g6768 ( 
.A(n_6250),
.B(n_4065),
.Y(n_6768)
);

INVx2_ASAP7_75t_L g6769 ( 
.A(n_6077),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6096),
.Y(n_6770)
);

NAND2xp5_ASAP7_75t_L g6771 ( 
.A(n_5862),
.B(n_3640),
.Y(n_6771)
);

NAND2xp5_ASAP7_75t_L g6772 ( 
.A(n_5869),
.B(n_3642),
.Y(n_6772)
);

INVx3_ASAP7_75t_L g6773 ( 
.A(n_5904),
.Y(n_6773)
);

INVx2_ASAP7_75t_L g6774 ( 
.A(n_6129),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_5907),
.B(n_3647),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6053),
.B(n_6221),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_6139),
.Y(n_6777)
);

CKINVDCx5p33_ASAP7_75t_R g6778 ( 
.A(n_5897),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6225),
.B(n_4072),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_5909),
.Y(n_6780)
);

INVx3_ASAP7_75t_L g6781 ( 
.A(n_5913),
.Y(n_6781)
);

AND2x4_ASAP7_75t_L g6782 ( 
.A(n_5816),
.B(n_3728),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_6159),
.Y(n_6783)
);

INVx2_ASAP7_75t_L g6784 ( 
.A(n_6165),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_5930),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_5975),
.Y(n_6786)
);

HB1xp67_ASAP7_75t_L g6787 ( 
.A(n_6010),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_6166),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6238),
.B(n_4072),
.Y(n_6789)
);

INVx2_ASAP7_75t_L g6790 ( 
.A(n_5994),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6029),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_6198),
.Y(n_6792)
);

BUFx2_ASAP7_75t_L g6793 ( 
.A(n_6317),
.Y(n_6793)
);

AND2x2_ASAP7_75t_L g6794 ( 
.A(n_6212),
.B(n_4093),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6087),
.Y(n_6795)
);

INVx1_ASAP7_75t_L g6796 ( 
.A(n_6337),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_5958),
.Y(n_6797)
);

INVx2_ASAP7_75t_L g6798 ( 
.A(n_5972),
.Y(n_6798)
);

BUFx6f_ASAP7_75t_L g6799 ( 
.A(n_5959),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6023),
.Y(n_6800)
);

INVx3_ASAP7_75t_L g6801 ( 
.A(n_6275),
.Y(n_6801)
);

BUFx6f_ASAP7_75t_L g6802 ( 
.A(n_6280),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_5817),
.Y(n_6803)
);

INVx1_ASAP7_75t_L g6804 ( 
.A(n_6223),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_SL g6805 ( 
.A(n_6036),
.B(n_3649),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6234),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_L g6807 ( 
.A(n_5903),
.B(n_5911),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6128),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_5951),
.Y(n_6809)
);

AND2x6_ASAP7_75t_L g6810 ( 
.A(n_6229),
.B(n_3738),
.Y(n_6810)
);

BUFx6f_ASAP7_75t_L g6811 ( 
.A(n_5974),
.Y(n_6811)
);

INVx2_ASAP7_75t_L g6812 ( 
.A(n_6239),
.Y(n_6812)
);

INVx2_ASAP7_75t_L g6813 ( 
.A(n_6254),
.Y(n_6813)
);

INVx3_ASAP7_75t_L g6814 ( 
.A(n_5976),
.Y(n_6814)
);

OA21x2_ASAP7_75t_L g6815 ( 
.A1(n_5834),
.A2(n_3765),
.B(n_3756),
.Y(n_6815)
);

INVx2_ASAP7_75t_L g6816 ( 
.A(n_6257),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_5903),
.B(n_3650),
.Y(n_6817)
);

AND2x4_ASAP7_75t_L g6818 ( 
.A(n_5858),
.B(n_3766),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6240),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6034),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6332),
.Y(n_6821)
);

AND2x2_ASAP7_75t_L g6822 ( 
.A(n_6287),
.B(n_4093),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6373),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6384),
.Y(n_6824)
);

INVx2_ASAP7_75t_L g6825 ( 
.A(n_6258),
.Y(n_6825)
);

INVx3_ASAP7_75t_L g6826 ( 
.A(n_6105),
.Y(n_6826)
);

INVxp67_ASAP7_75t_L g6827 ( 
.A(n_6294),
.Y(n_6827)
);

INVx2_ASAP7_75t_L g6828 ( 
.A(n_6264),
.Y(n_6828)
);

BUFx6f_ASAP7_75t_L g6829 ( 
.A(n_5877),
.Y(n_6829)
);

INVx2_ASAP7_75t_L g6830 ( 
.A(n_6268),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6132),
.Y(n_6831)
);

BUFx2_ASAP7_75t_L g6832 ( 
.A(n_6065),
.Y(n_6832)
);

OR2x2_ASAP7_75t_L g6833 ( 
.A(n_6352),
.B(n_3652),
.Y(n_6833)
);

AND2x4_ASAP7_75t_L g6834 ( 
.A(n_6327),
.B(n_3777),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6182),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_5911),
.B(n_3653),
.Y(n_6836)
);

BUFx2_ASAP7_75t_L g6837 ( 
.A(n_6065),
.Y(n_6837)
);

INVx2_ASAP7_75t_L g6838 ( 
.A(n_6279),
.Y(n_6838)
);

AND2x4_ASAP7_75t_L g6839 ( 
.A(n_6343),
.B(n_3781),
.Y(n_6839)
);

NAND2xp5_ASAP7_75t_SL g6840 ( 
.A(n_6203),
.B(n_3657),
.Y(n_6840)
);

INVx2_ASAP7_75t_L g6841 ( 
.A(n_6339),
.Y(n_6841)
);

NAND2xp5_ASAP7_75t_SL g6842 ( 
.A(n_6270),
.B(n_3660),
.Y(n_6842)
);

BUFx2_ASAP7_75t_L g6843 ( 
.A(n_6070),
.Y(n_6843)
);

BUFx2_ASAP7_75t_L g6844 ( 
.A(n_6070),
.Y(n_6844)
);

BUFx2_ASAP7_75t_L g6845 ( 
.A(n_6181),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_5882),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_5888),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6339),
.Y(n_6848)
);

BUFx8_ASAP7_75t_L g6849 ( 
.A(n_6044),
.Y(n_6849)
);

BUFx6f_ASAP7_75t_L g6850 ( 
.A(n_6365),
.Y(n_6850)
);

INVx3_ASAP7_75t_L g6851 ( 
.A(n_6153),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6347),
.Y(n_6852)
);

BUFx6f_ASAP7_75t_L g6853 ( 
.A(n_6227),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6347),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6286),
.B(n_4125),
.Y(n_6855)
);

HB1xp67_ASAP7_75t_L g6856 ( 
.A(n_6116),
.Y(n_6856)
);

BUFx6f_ASAP7_75t_L g6857 ( 
.A(n_6237),
.Y(n_6857)
);

INVx2_ASAP7_75t_L g6858 ( 
.A(n_5983),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6228),
.B(n_3661),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_L g6860 ( 
.A(n_6278),
.B(n_6282),
.Y(n_6860)
);

AND2x6_ASAP7_75t_L g6861 ( 
.A(n_6243),
.B(n_3784),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6278),
.B(n_3662),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_5998),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_5865),
.Y(n_6864)
);

INVx2_ASAP7_75t_L g6865 ( 
.A(n_5983),
.Y(n_6865)
);

INVx2_ASAP7_75t_L g6866 ( 
.A(n_6018),
.Y(n_6866)
);

INVx1_ASAP7_75t_L g6867 ( 
.A(n_6020),
.Y(n_6867)
);

BUFx6f_ASAP7_75t_L g6868 ( 
.A(n_6246),
.Y(n_6868)
);

CKINVDCx8_ASAP7_75t_R g6869 ( 
.A(n_5929),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6021),
.Y(n_6870)
);

BUFx6f_ASAP7_75t_L g6871 ( 
.A(n_6253),
.Y(n_6871)
);

BUFx6f_ASAP7_75t_L g6872 ( 
.A(n_6261),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6006),
.Y(n_6873)
);

NAND2xp5_ASAP7_75t_L g6874 ( 
.A(n_6282),
.B(n_3663),
.Y(n_6874)
);

BUFx6f_ASAP7_75t_L g6875 ( 
.A(n_6274),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_5892),
.Y(n_6876)
);

INVx1_ASAP7_75t_L g6877 ( 
.A(n_5942),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6018),
.B(n_3664),
.Y(n_6878)
);

INVx2_ASAP7_75t_L g6879 ( 
.A(n_6245),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_5852),
.Y(n_6880)
);

INVx3_ASAP7_75t_L g6881 ( 
.A(n_6308),
.Y(n_6881)
);

BUFx8_ASAP7_75t_L g6882 ( 
.A(n_6052),
.Y(n_6882)
);

NAND2xp5_ASAP7_75t_L g6883 ( 
.A(n_6027),
.B(n_3665),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_6247),
.Y(n_6884)
);

INVx3_ASAP7_75t_L g6885 ( 
.A(n_6316),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6251),
.Y(n_6886)
);

NOR2xp33_ASAP7_75t_L g6887 ( 
.A(n_6230),
.B(n_3669),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6252),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_6255),
.Y(n_6889)
);

NOR2xp33_ASAP7_75t_L g6890 ( 
.A(n_6236),
.B(n_3670),
.Y(n_6890)
);

INVx2_ASAP7_75t_L g6891 ( 
.A(n_6262),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6263),
.Y(n_6892)
);

INVx2_ASAP7_75t_L g6893 ( 
.A(n_6265),
.Y(n_6893)
);

INVx1_ASAP7_75t_SL g6894 ( 
.A(n_6131),
.Y(n_6894)
);

INVx2_ASAP7_75t_L g6895 ( 
.A(n_6269),
.Y(n_6895)
);

BUFx6f_ASAP7_75t_L g6896 ( 
.A(n_6267),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6271),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6272),
.Y(n_6898)
);

NAND2xp5_ASAP7_75t_SL g6899 ( 
.A(n_5819),
.B(n_3672),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_6276),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_6277),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6248),
.B(n_4125),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6075),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6283),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6114),
.Y(n_6905)
);

NOR2xp33_ASAP7_75t_R g6906 ( 
.A(n_5950),
.B(n_4674),
.Y(n_6906)
);

NAND2xp5_ASAP7_75t_SL g6907 ( 
.A(n_5876),
.B(n_3673),
.Y(n_6907)
);

AOI22xp5_ASAP7_75t_L g6908 ( 
.A1(n_6289),
.A2(n_4693),
.B1(n_4710),
.B2(n_4684),
.Y(n_6908)
);

OAI22xp5_ASAP7_75t_SL g6909 ( 
.A1(n_6108),
.A2(n_4738),
.B1(n_4761),
.B2(n_4713),
.Y(n_6909)
);

OA21x2_ASAP7_75t_L g6910 ( 
.A1(n_6043),
.A2(n_3791),
.B(n_3785),
.Y(n_6910)
);

NAND2xp33_ASAP7_75t_L g6911 ( 
.A(n_6027),
.B(n_3677),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_SL g6912 ( 
.A(n_6122),
.B(n_3678),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6008),
.Y(n_6913)
);

OAI21x1_ASAP7_75t_L g6914 ( 
.A1(n_6293),
.A2(n_4535),
.B(n_4512),
.Y(n_6914)
);

NOR2xp33_ASAP7_75t_L g6915 ( 
.A(n_6013),
.B(n_3680),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6273),
.B(n_4187),
.Y(n_6916)
);

BUFx8_ASAP7_75t_L g6917 ( 
.A(n_6073),
.Y(n_6917)
);

NAND2xp5_ASAP7_75t_L g6918 ( 
.A(n_6063),
.B(n_3682),
.Y(n_6918)
);

INVx3_ASAP7_75t_L g6919 ( 
.A(n_6118),
.Y(n_6919)
);

BUFx6f_ASAP7_75t_L g6920 ( 
.A(n_6291),
.Y(n_6920)
);

INVx1_ASAP7_75t_SL g6921 ( 
.A(n_6112),
.Y(n_6921)
);

NAND2xp5_ASAP7_75t_SL g6922 ( 
.A(n_6326),
.B(n_3683),
.Y(n_6922)
);

BUFx6f_ASAP7_75t_L g6923 ( 
.A(n_6092),
.Y(n_6923)
);

INVx1_ASAP7_75t_SL g6924 ( 
.A(n_6145),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6296),
.Y(n_6925)
);

BUFx6f_ASAP7_75t_L g6926 ( 
.A(n_6224),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6298),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_L g6928 ( 
.A(n_6358),
.B(n_3684),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_L g6929 ( 
.A(n_6395),
.B(n_3688),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6039),
.B(n_4187),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_6300),
.Y(n_6931)
);

BUFx6f_ASAP7_75t_L g6932 ( 
.A(n_5879),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_5991),
.Y(n_6933)
);

INVx3_ASAP7_75t_L g6934 ( 
.A(n_6193),
.Y(n_6934)
);

BUFx6f_ASAP7_75t_L g6935 ( 
.A(n_5898),
.Y(n_6935)
);

OA21x2_ASAP7_75t_L g6936 ( 
.A1(n_6097),
.A2(n_3802),
.B(n_3796),
.Y(n_6936)
);

BUFx6f_ASAP7_75t_L g6937 ( 
.A(n_5914),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6292),
.Y(n_6938)
);

AND2x4_ASAP7_75t_L g6939 ( 
.A(n_6302),
.B(n_3807),
.Y(n_6939)
);

INVx2_ASAP7_75t_L g6940 ( 
.A(n_6120),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6123),
.B(n_6284),
.Y(n_6941)
);

BUFx2_ASAP7_75t_L g6942 ( 
.A(n_6306),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6305),
.Y(n_6943)
);

NAND2xp5_ASAP7_75t_L g6944 ( 
.A(n_6301),
.B(n_3689),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6309),
.Y(n_6945)
);

AND2x4_ASAP7_75t_L g6946 ( 
.A(n_6310),
.B(n_6311),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6314),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6318),
.Y(n_6948)
);

NAND2xp5_ASAP7_75t_L g6949 ( 
.A(n_6080),
.B(n_6103),
.Y(n_6949)
);

INVx2_ASAP7_75t_L g6950 ( 
.A(n_6202),
.Y(n_6950)
);

BUFx6f_ASAP7_75t_L g6951 ( 
.A(n_5952),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6288),
.Y(n_6952)
);

INVx2_ASAP7_75t_L g6953 ( 
.A(n_6158),
.Y(n_6953)
);

NAND2xp5_ASAP7_75t_L g6954 ( 
.A(n_6218),
.B(n_3690),
.Y(n_6954)
);

CKINVDCx5p33_ASAP7_75t_R g6955 ( 
.A(n_6222),
.Y(n_6955)
);

NAND2xp5_ASAP7_75t_SL g6956 ( 
.A(n_6333),
.B(n_3694),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6281),
.Y(n_6957)
);

BUFx2_ASAP7_75t_L g6958 ( 
.A(n_6460),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6398),
.Y(n_6959)
);

NAND2xp5_ASAP7_75t_L g6960 ( 
.A(n_6722),
.B(n_3695),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_6397),
.Y(n_6961)
);

NOR2xp33_ASAP7_75t_L g6962 ( 
.A(n_6732),
.B(n_6215),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_6726),
.B(n_3699),
.Y(n_6963)
);

NAND2xp5_ASAP7_75t_L g6964 ( 
.A(n_6728),
.B(n_3700),
.Y(n_6964)
);

NAND2xp5_ASAP7_75t_SL g6965 ( 
.A(n_6488),
.B(n_5977),
.Y(n_6965)
);

INVx3_ASAP7_75t_L g6966 ( 
.A(n_6618),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6399),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6410),
.Y(n_6968)
);

INVx2_ASAP7_75t_L g6969 ( 
.A(n_6402),
.Y(n_6969)
);

NAND2xp5_ASAP7_75t_L g6970 ( 
.A(n_6631),
.B(n_6634),
.Y(n_6970)
);

NAND2xp5_ASAP7_75t_SL g6971 ( 
.A(n_6721),
.B(n_6433),
.Y(n_6971)
);

INVx5_ASAP7_75t_L g6972 ( 
.A(n_6423),
.Y(n_6972)
);

NAND2xp33_ASAP7_75t_L g6973 ( 
.A(n_6635),
.B(n_3704),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_6414),
.Y(n_6974)
);

AND2x2_ASAP7_75t_L g6975 ( 
.A(n_6436),
.B(n_5992),
.Y(n_6975)
);

INVx3_ASAP7_75t_L g6976 ( 
.A(n_6618),
.Y(n_6976)
);

NOR2xp33_ASAP7_75t_L g6977 ( 
.A(n_6532),
.B(n_6084),
.Y(n_6977)
);

INVx2_ASAP7_75t_L g6978 ( 
.A(n_6411),
.Y(n_6978)
);

NAND2xp5_ASAP7_75t_L g6979 ( 
.A(n_6636),
.B(n_3711),
.Y(n_6979)
);

NOR2xp33_ASAP7_75t_L g6980 ( 
.A(n_6453),
.B(n_6111),
.Y(n_6980)
);

INVx2_ASAP7_75t_L g6981 ( 
.A(n_6413),
.Y(n_6981)
);

NAND2xp5_ASAP7_75t_SL g6982 ( 
.A(n_6776),
.B(n_6157),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6522),
.B(n_6115),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_SL g6984 ( 
.A(n_6879),
.B(n_6174),
.Y(n_6984)
);

INVx2_ASAP7_75t_L g6985 ( 
.A(n_6418),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6415),
.Y(n_6986)
);

INVx3_ASAP7_75t_L g6987 ( 
.A(n_6644),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_6434),
.Y(n_6988)
);

BUFx6f_ASAP7_75t_SL g6989 ( 
.A(n_6423),
.Y(n_6989)
);

INVx4_ASAP7_75t_L g6990 ( 
.A(n_6853),
.Y(n_6990)
);

BUFx6f_ASAP7_75t_L g6991 ( 
.A(n_6640),
.Y(n_6991)
);

NOR2xp33_ASAP7_75t_L g6992 ( 
.A(n_6406),
.B(n_6183),
.Y(n_6992)
);

BUFx6f_ASAP7_75t_L g6993 ( 
.A(n_6640),
.Y(n_6993)
);

INVx2_ASAP7_75t_SL g6994 ( 
.A(n_6466),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6435),
.Y(n_6995)
);

OAI22xp5_ASAP7_75t_L g6996 ( 
.A1(n_6913),
.A2(n_4792),
.B1(n_4793),
.B2(n_4783),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_6416),
.Y(n_6997)
);

AOI22xp33_ASAP7_75t_L g6998 ( 
.A1(n_6880),
.A2(n_4816),
.B1(n_4819),
.B2(n_4803),
.Y(n_6998)
);

INVx3_ASAP7_75t_L g6999 ( 
.A(n_6644),
.Y(n_6999)
);

OAI22xp33_ASAP7_75t_L g7000 ( 
.A1(n_6835),
.A2(n_6205),
.B1(n_6364),
.B2(n_5966),
.Y(n_7000)
);

NAND2xp5_ASAP7_75t_L g7001 ( 
.A(n_6638),
.B(n_6642),
.Y(n_7001)
);

NOR2xp33_ASAP7_75t_L g7002 ( 
.A(n_6429),
.B(n_5823),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6417),
.Y(n_7003)
);

AND2x6_ASAP7_75t_L g7004 ( 
.A(n_6396),
.B(n_3809),
.Y(n_7004)
);

OAI22xp33_ASAP7_75t_L g7005 ( 
.A1(n_6876),
.A2(n_6330),
.B1(n_5880),
.B2(n_4840),
.Y(n_7005)
);

INVx3_ASAP7_75t_L g7006 ( 
.A(n_6655),
.Y(n_7006)
);

INVx2_ASAP7_75t_L g7007 ( 
.A(n_6461),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6420),
.Y(n_7008)
);

INVx2_ASAP7_75t_L g7009 ( 
.A(n_6421),
.Y(n_7009)
);

NOR2xp33_ASAP7_75t_L g7010 ( 
.A(n_6752),
.B(n_6235),
.Y(n_7010)
);

INVx2_ASAP7_75t_SL g7011 ( 
.A(n_6605),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6422),
.Y(n_7012)
);

INVx2_ASAP7_75t_L g7013 ( 
.A(n_6427),
.Y(n_7013)
);

INVx2_ASAP7_75t_L g7014 ( 
.A(n_6430),
.Y(n_7014)
);

INVx6_ASAP7_75t_L g7015 ( 
.A(n_6799),
.Y(n_7015)
);

INVxp67_ASAP7_75t_SL g7016 ( 
.A(n_6591),
.Y(n_7016)
);

INVx2_ASAP7_75t_L g7017 ( 
.A(n_6432),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6439),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6443),
.Y(n_7019)
);

BUFx6f_ASAP7_75t_L g7020 ( 
.A(n_6799),
.Y(n_7020)
);

INVx3_ASAP7_75t_L g7021 ( 
.A(n_6655),
.Y(n_7021)
);

NAND3xp33_ASAP7_75t_L g7022 ( 
.A(n_6915),
.B(n_3716),
.C(n_3712),
.Y(n_7022)
);

NAND2xp5_ASAP7_75t_L g7023 ( 
.A(n_6643),
.B(n_3718),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6446),
.Y(n_7024)
);

INVx2_ASAP7_75t_L g7025 ( 
.A(n_6447),
.Y(n_7025)
);

INVx3_ASAP7_75t_L g7026 ( 
.A(n_6675),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6452),
.Y(n_7027)
);

BUFx6f_ASAP7_75t_L g7028 ( 
.A(n_6811),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6454),
.Y(n_7029)
);

OAI22xp5_ASAP7_75t_L g7030 ( 
.A1(n_6877),
.A2(n_4854),
.B1(n_4871),
.B2(n_4833),
.Y(n_7030)
);

INVx2_ASAP7_75t_L g7031 ( 
.A(n_6458),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6463),
.Y(n_7032)
);

AND2x2_ASAP7_75t_L g7033 ( 
.A(n_6551),
.B(n_4288),
.Y(n_7033)
);

BUFx3_ASAP7_75t_L g7034 ( 
.A(n_6811),
.Y(n_7034)
);

NAND2xp5_ASAP7_75t_L g7035 ( 
.A(n_6645),
.B(n_3722),
.Y(n_7035)
);

NOR2xp33_ASAP7_75t_L g7036 ( 
.A(n_6602),
.B(n_6604),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6465),
.Y(n_7037)
);

NAND2xp5_ASAP7_75t_L g7038 ( 
.A(n_6647),
.B(n_6650),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6468),
.Y(n_7039)
);

INVx2_ASAP7_75t_L g7040 ( 
.A(n_6469),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_L g7041 ( 
.A1(n_6809),
.A2(n_4543),
.B1(n_4566),
.B2(n_4541),
.Y(n_7041)
);

INVx2_ASAP7_75t_SL g7042 ( 
.A(n_6626),
.Y(n_7042)
);

NAND2xp5_ASAP7_75t_L g7043 ( 
.A(n_6652),
.B(n_3724),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6470),
.Y(n_7044)
);

INVx2_ASAP7_75t_L g7045 ( 
.A(n_6473),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_6553),
.B(n_4288),
.Y(n_7046)
);

BUFx6f_ASAP7_75t_L g7047 ( 
.A(n_6853),
.Y(n_7047)
);

NOR2xp33_ASAP7_75t_L g7048 ( 
.A(n_6487),
.B(n_3725),
.Y(n_7048)
);

AND3x1_ASAP7_75t_L g7049 ( 
.A(n_6533),
.B(n_6908),
.C(n_6680),
.Y(n_7049)
);

INVx2_ASAP7_75t_SL g7050 ( 
.A(n_6633),
.Y(n_7050)
);

NAND2xp5_ASAP7_75t_SL g7051 ( 
.A(n_6888),
.B(n_3730),
.Y(n_7051)
);

INVx2_ASAP7_75t_L g7052 ( 
.A(n_6477),
.Y(n_7052)
);

INVx3_ASAP7_75t_L g7053 ( 
.A(n_6675),
.Y(n_7053)
);

INVx3_ASAP7_75t_L g7054 ( 
.A(n_6679),
.Y(n_7054)
);

OR2x2_ASAP7_75t_L g7055 ( 
.A(n_6504),
.B(n_3732),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_6479),
.Y(n_7056)
);

AOI22xp5_ASAP7_75t_L g7057 ( 
.A1(n_6654),
.A2(n_3734),
.B1(n_3735),
.B2(n_3733),
.Y(n_7057)
);

NAND2xp5_ASAP7_75t_L g7058 ( 
.A(n_6656),
.B(n_3740),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_6480),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6484),
.Y(n_7060)
);

INVx3_ASAP7_75t_L g7061 ( 
.A(n_6679),
.Y(n_7061)
);

INVx2_ASAP7_75t_L g7062 ( 
.A(n_6491),
.Y(n_7062)
);

INVx2_ASAP7_75t_SL g7063 ( 
.A(n_6407),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_6493),
.Y(n_7064)
);

NAND2xp5_ASAP7_75t_L g7065 ( 
.A(n_6450),
.B(n_6890),
.Y(n_7065)
);

CKINVDCx6p67_ASAP7_75t_R g7066 ( 
.A(n_6609),
.Y(n_7066)
);

AND2x4_ASAP7_75t_L g7067 ( 
.A(n_6405),
.B(n_3818),
.Y(n_7067)
);

INVx2_ASAP7_75t_SL g7068 ( 
.A(n_6472),
.Y(n_7068)
);

INVxp67_ASAP7_75t_L g7069 ( 
.A(n_6431),
.Y(n_7069)
);

AND2x2_ASAP7_75t_L g7070 ( 
.A(n_6717),
.B(n_4333),
.Y(n_7070)
);

NAND3xp33_ASAP7_75t_L g7071 ( 
.A(n_6887),
.B(n_3742),
.C(n_3741),
.Y(n_7071)
);

INVx1_ASAP7_75t_L g7072 ( 
.A(n_6495),
.Y(n_7072)
);

INVx2_ASAP7_75t_SL g7073 ( 
.A(n_6544),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6497),
.Y(n_7074)
);

INVx2_ASAP7_75t_L g7075 ( 
.A(n_6498),
.Y(n_7075)
);

INVx2_ASAP7_75t_L g7076 ( 
.A(n_6499),
.Y(n_7076)
);

NOR2xp33_ASAP7_75t_L g7077 ( 
.A(n_6666),
.B(n_3743),
.Y(n_7077)
);

INVx2_ASAP7_75t_L g7078 ( 
.A(n_6501),
.Y(n_7078)
);

NAND2xp5_ASAP7_75t_L g7079 ( 
.A(n_6653),
.B(n_6729),
.Y(n_7079)
);

INVx2_ASAP7_75t_L g7080 ( 
.A(n_6502),
.Y(n_7080)
);

AND2x2_ASAP7_75t_L g7081 ( 
.A(n_6794),
.B(n_4333),
.Y(n_7081)
);

OR2x6_ASAP7_75t_L g7082 ( 
.A(n_6857),
.B(n_6232),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6508),
.Y(n_7083)
);

INVx2_ASAP7_75t_L g7084 ( 
.A(n_6511),
.Y(n_7084)
);

CKINVDCx5p33_ASAP7_75t_R g7085 ( 
.A(n_6462),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6730),
.B(n_3746),
.Y(n_7086)
);

NOR2xp33_ASAP7_75t_L g7087 ( 
.A(n_6954),
.B(n_3749),
.Y(n_7087)
);

NAND2xp5_ASAP7_75t_L g7088 ( 
.A(n_6731),
.B(n_3750),
.Y(n_7088)
);

INVxp33_ASAP7_75t_SL g7089 ( 
.A(n_6906),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_6514),
.Y(n_7090)
);

INVx1_ASAP7_75t_SL g7091 ( 
.A(n_6586),
.Y(n_7091)
);

INVx2_ASAP7_75t_L g7092 ( 
.A(n_6515),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6516),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_L g7094 ( 
.A(n_6733),
.B(n_3751),
.Y(n_7094)
);

INVx1_ASAP7_75t_SL g7095 ( 
.A(n_6921),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_6467),
.B(n_4458),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_SL g7097 ( 
.A(n_6889),
.B(n_3752),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_6517),
.Y(n_7098)
);

BUFx6f_ASAP7_75t_L g7099 ( 
.A(n_6857),
.Y(n_7099)
);

NAND2xp33_ASAP7_75t_L g7100 ( 
.A(n_6861),
.B(n_3753),
.Y(n_7100)
);

OAI22xp33_ASAP7_75t_L g7101 ( 
.A1(n_6821),
.A2(n_3755),
.B1(n_3759),
.B2(n_3754),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6518),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6520),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_6524),
.Y(n_7104)
);

AND2x2_ASAP7_75t_L g7105 ( 
.A(n_6486),
.B(n_4458),
.Y(n_7105)
);

OAI22xp5_ASAP7_75t_L g7106 ( 
.A1(n_6820),
.A2(n_3761),
.B1(n_3763),
.B2(n_3760),
.Y(n_7106)
);

NAND2xp5_ASAP7_75t_SL g7107 ( 
.A(n_6891),
.B(n_3768),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6525),
.Y(n_7108)
);

INVx2_ASAP7_75t_L g7109 ( 
.A(n_6528),
.Y(n_7109)
);

INVx4_ASAP7_75t_L g7110 ( 
.A(n_6868),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6531),
.Y(n_7111)
);

CKINVDCx20_ASAP7_75t_R g7112 ( 
.A(n_6572),
.Y(n_7112)
);

NAND2xp5_ASAP7_75t_SL g7113 ( 
.A(n_6893),
.B(n_3769),
.Y(n_7113)
);

INVx2_ASAP7_75t_L g7114 ( 
.A(n_6534),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6535),
.Y(n_7115)
);

OAI22xp5_ASAP7_75t_L g7116 ( 
.A1(n_6823),
.A2(n_3771),
.B1(n_3772),
.B2(n_3770),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6401),
.B(n_3774),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6400),
.B(n_3779),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_6536),
.Y(n_7119)
);

INVx3_ASAP7_75t_L g7120 ( 
.A(n_6682),
.Y(n_7120)
);

NAND2xp5_ASAP7_75t_SL g7121 ( 
.A(n_6895),
.B(n_3780),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_SL g7122 ( 
.A(n_6900),
.B(n_6931),
.Y(n_7122)
);

BUFx10_ASAP7_75t_L g7123 ( 
.A(n_6829),
.Y(n_7123)
);

INVx2_ASAP7_75t_L g7124 ( 
.A(n_6542),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_6587),
.B(n_6607),
.Y(n_7125)
);

AO21x2_ASAP7_75t_L g7126 ( 
.A1(n_6664),
.A2(n_3821),
.B(n_3819),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6543),
.Y(n_7127)
);

INVx2_ASAP7_75t_L g7128 ( 
.A(n_6545),
.Y(n_7128)
);

INVx3_ASAP7_75t_L g7129 ( 
.A(n_6682),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_6546),
.Y(n_7130)
);

BUFx6f_ASAP7_75t_L g7131 ( 
.A(n_6868),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6594),
.B(n_3782),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_SL g7133 ( 
.A(n_6884),
.B(n_3783),
.Y(n_7133)
);

INVx2_ASAP7_75t_SL g7134 ( 
.A(n_6566),
.Y(n_7134)
);

INVx2_ASAP7_75t_L g7135 ( 
.A(n_6547),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_6550),
.Y(n_7136)
);

NAND2xp5_ASAP7_75t_L g7137 ( 
.A(n_6557),
.B(n_3786),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6563),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6568),
.Y(n_7139)
);

BUFx10_ASAP7_75t_L g7140 ( 
.A(n_6829),
.Y(n_7140)
);

CKINVDCx5p33_ASAP7_75t_R g7141 ( 
.A(n_6778),
.Y(n_7141)
);

NAND2xp5_ASAP7_75t_L g7142 ( 
.A(n_6570),
.B(n_3788),
.Y(n_7142)
);

BUFx3_ASAP7_75t_L g7143 ( 
.A(n_6871),
.Y(n_7143)
);

BUFx3_ASAP7_75t_L g7144 ( 
.A(n_6871),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6629),
.Y(n_7145)
);

AND3x2_ASAP7_75t_L g7146 ( 
.A(n_6613),
.B(n_3826),
.C(n_3823),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6573),
.Y(n_7147)
);

INVx2_ASAP7_75t_L g7148 ( 
.A(n_6630),
.Y(n_7148)
);

OR2x6_ASAP7_75t_L g7149 ( 
.A(n_6872),
.B(n_3836),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_6575),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6578),
.Y(n_7151)
);

BUFx2_ASAP7_75t_L g7152 ( 
.A(n_6856),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6581),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_L g7154 ( 
.A(n_6677),
.B(n_3789),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6588),
.Y(n_7155)
);

NAND2xp5_ASAP7_75t_L g7156 ( 
.A(n_6707),
.B(n_3792),
.Y(n_7156)
);

INVx1_ASAP7_75t_L g7157 ( 
.A(n_6593),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6596),
.Y(n_7158)
);

INVx3_ASAP7_75t_L g7159 ( 
.A(n_6686),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6597),
.Y(n_7160)
);

BUFx4f_ASAP7_75t_L g7161 ( 
.A(n_6850),
.Y(n_7161)
);

INVx3_ASAP7_75t_L g7162 ( 
.A(n_6686),
.Y(n_7162)
);

CKINVDCx5p33_ASAP7_75t_R g7163 ( 
.A(n_6955),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_6599),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_SL g7165 ( 
.A(n_6886),
.B(n_3797),
.Y(n_7165)
);

INVx4_ASAP7_75t_L g7166 ( 
.A(n_6872),
.Y(n_7166)
);

INVx3_ASAP7_75t_L g7167 ( 
.A(n_6704),
.Y(n_7167)
);

NAND2xp5_ASAP7_75t_SL g7168 ( 
.A(n_6892),
.B(n_3799),
.Y(n_7168)
);

INVxp67_ASAP7_75t_SL g7169 ( 
.A(n_6591),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_6603),
.Y(n_7170)
);

NAND2xp5_ASAP7_75t_SL g7171 ( 
.A(n_6897),
.B(n_3800),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_SL g7172 ( 
.A(n_6898),
.B(n_3808),
.Y(n_7172)
);

BUFx6f_ASAP7_75t_L g7173 ( 
.A(n_6875),
.Y(n_7173)
);

BUFx3_ASAP7_75t_L g7174 ( 
.A(n_6875),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6606),
.Y(n_7175)
);

INVx2_ASAP7_75t_L g7176 ( 
.A(n_6464),
.Y(n_7176)
);

OR2x6_ASAP7_75t_L g7177 ( 
.A(n_6920),
.B(n_3837),
.Y(n_7177)
);

INVx2_ASAP7_75t_L g7178 ( 
.A(n_6471),
.Y(n_7178)
);

INVx2_ASAP7_75t_L g7179 ( 
.A(n_6475),
.Y(n_7179)
);

INVx4_ASAP7_75t_L g7180 ( 
.A(n_6920),
.Y(n_7180)
);

INVx3_ASAP7_75t_L g7181 ( 
.A(n_6704),
.Y(n_7181)
);

NOR2xp33_ASAP7_75t_R g7182 ( 
.A(n_6869),
.B(n_3812),
.Y(n_7182)
);

OR2x2_ASAP7_75t_L g7183 ( 
.A(n_6819),
.B(n_3813),
.Y(n_7183)
);

INVx2_ASAP7_75t_L g7184 ( 
.A(n_6478),
.Y(n_7184)
);

BUFx6f_ASAP7_75t_L g7185 ( 
.A(n_6440),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6482),
.Y(n_7186)
);

AND2x2_ASAP7_75t_L g7187 ( 
.A(n_6779),
.B(n_4502),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_6617),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_6619),
.Y(n_7189)
);

INVx2_ASAP7_75t_L g7190 ( 
.A(n_6483),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_6622),
.Y(n_7191)
);

BUFx4f_ASAP7_75t_L g7192 ( 
.A(n_6850),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_6623),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_6444),
.Y(n_7194)
);

HB1xp67_ASAP7_75t_L g7195 ( 
.A(n_6590),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_6490),
.Y(n_7196)
);

NAND2xp5_ASAP7_75t_L g7197 ( 
.A(n_6724),
.B(n_3817),
.Y(n_7197)
);

NOR2xp33_ASAP7_75t_L g7198 ( 
.A(n_6611),
.B(n_3820),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6494),
.Y(n_7199)
);

INVx2_ASAP7_75t_L g7200 ( 
.A(n_6500),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_6756),
.B(n_3822),
.Y(n_7201)
);

INVx2_ASAP7_75t_L g7202 ( 
.A(n_6509),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_6510),
.Y(n_7203)
);

NAND2xp5_ASAP7_75t_SL g7204 ( 
.A(n_6901),
.B(n_6927),
.Y(n_7204)
);

BUFx4f_ASAP7_75t_L g7205 ( 
.A(n_6896),
.Y(n_7205)
);

INVx2_ASAP7_75t_L g7206 ( 
.A(n_6529),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6530),
.Y(n_7207)
);

NAND3xp33_ASAP7_75t_L g7208 ( 
.A(n_6456),
.B(n_6806),
.C(n_6804),
.Y(n_7208)
);

INVx2_ASAP7_75t_L g7209 ( 
.A(n_6540),
.Y(n_7209)
);

INVx5_ASAP7_75t_L g7210 ( 
.A(n_6896),
.Y(n_7210)
);

INVx2_ASAP7_75t_L g7211 ( 
.A(n_6541),
.Y(n_7211)
);

NOR2xp33_ASAP7_75t_L g7212 ( 
.A(n_6657),
.B(n_3824),
.Y(n_7212)
);

INVx2_ASAP7_75t_L g7213 ( 
.A(n_6554),
.Y(n_7213)
);

AND3x2_ASAP7_75t_L g7214 ( 
.A(n_6761),
.B(n_3852),
.C(n_3841),
.Y(n_7214)
);

CKINVDCx20_ASAP7_75t_R g7215 ( 
.A(n_6715),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_6556),
.Y(n_7216)
);

OAI22xp33_ASAP7_75t_L g7217 ( 
.A1(n_6824),
.A2(n_3831),
.B1(n_3832),
.B2(n_3828),
.Y(n_7217)
);

AOI22xp5_ASAP7_75t_L g7218 ( 
.A1(n_6831),
.A2(n_3838),
.B1(n_3842),
.B2(n_3835),
.Y(n_7218)
);

CKINVDCx5p33_ASAP7_75t_R g7219 ( 
.A(n_6793),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6560),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_6561),
.Y(n_7221)
);

OAI21xp33_ASAP7_75t_SL g7222 ( 
.A1(n_6796),
.A2(n_3854),
.B(n_3853),
.Y(n_7222)
);

NAND2xp5_ASAP7_75t_L g7223 ( 
.A(n_6812),
.B(n_3851),
.Y(n_7223)
);

AOI22xp5_ASAP7_75t_L g7224 ( 
.A1(n_6616),
.A2(n_3858),
.B1(n_3859),
.B2(n_3856),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_6562),
.Y(n_7225)
);

NAND3xp33_ASAP7_75t_L g7226 ( 
.A(n_6938),
.B(n_3861),
.C(n_3860),
.Y(n_7226)
);

NAND2xp5_ASAP7_75t_SL g7227 ( 
.A(n_6813),
.B(n_3862),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6565),
.Y(n_7228)
);

INVx2_ASAP7_75t_L g7229 ( 
.A(n_6582),
.Y(n_7229)
);

AND2x2_ASAP7_75t_L g7230 ( 
.A(n_6789),
.B(n_4502),
.Y(n_7230)
);

NAND2xp5_ASAP7_75t_L g7231 ( 
.A(n_6816),
.B(n_3866),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_6583),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_6601),
.Y(n_7233)
);

INVx2_ASAP7_75t_L g7234 ( 
.A(n_6615),
.Y(n_7234)
);

INVx2_ASAP7_75t_L g7235 ( 
.A(n_6437),
.Y(n_7235)
);

NOR2xp33_ASAP7_75t_L g7236 ( 
.A(n_6827),
.B(n_6903),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_6438),
.Y(n_7237)
);

NOR2xp33_ASAP7_75t_L g7238 ( 
.A(n_6905),
.B(n_3867),
.Y(n_7238)
);

NAND2xp5_ASAP7_75t_L g7239 ( 
.A(n_6825),
.B(n_3872),
.Y(n_7239)
);

INVx2_ASAP7_75t_L g7240 ( 
.A(n_6441),
.Y(n_7240)
);

INVx4_ASAP7_75t_L g7241 ( 
.A(n_6802),
.Y(n_7241)
);

INVx2_ASAP7_75t_SL g7242 ( 
.A(n_6595),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_6442),
.Y(n_7243)
);

INVx2_ASAP7_75t_L g7244 ( 
.A(n_6449),
.Y(n_7244)
);

INVx3_ASAP7_75t_L g7245 ( 
.A(n_6708),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6694),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_6457),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_SL g7248 ( 
.A(n_6828),
.B(n_3876),
.Y(n_7248)
);

INVx5_ASAP7_75t_L g7249 ( 
.A(n_6802),
.Y(n_7249)
);

NOR2xp33_ASAP7_75t_L g7250 ( 
.A(n_6949),
.B(n_3881),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_6695),
.Y(n_7251)
);

OAI22xp33_ASAP7_75t_L g7252 ( 
.A1(n_6846),
.A2(n_3886),
.B1(n_3889),
.B2(n_3884),
.Y(n_7252)
);

INVx6_ASAP7_75t_L g7253 ( 
.A(n_6849),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_SL g7254 ( 
.A(n_6830),
.B(n_3890),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_6696),
.Y(n_7255)
);

NAND2xp5_ASAP7_75t_SL g7256 ( 
.A(n_6838),
.B(n_3894),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_6698),
.Y(n_7257)
);

BUFx6f_ASAP7_75t_L g7258 ( 
.A(n_6440),
.Y(n_7258)
);

INVx3_ASAP7_75t_L g7259 ( 
.A(n_6708),
.Y(n_7259)
);

INVx2_ASAP7_75t_L g7260 ( 
.A(n_6632),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_6699),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_6702),
.Y(n_7262)
);

NAND2xp33_ASAP7_75t_SL g7263 ( 
.A(n_6807),
.B(n_3895),
.Y(n_7263)
);

BUFx6f_ASAP7_75t_SL g7264 ( 
.A(n_6558),
.Y(n_7264)
);

INVx3_ASAP7_75t_L g7265 ( 
.A(n_6713),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_6703),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_6639),
.Y(n_7267)
);

INVx2_ASAP7_75t_L g7268 ( 
.A(n_6651),
.Y(n_7268)
);

NOR2xp33_ASAP7_75t_L g7269 ( 
.A(n_6942),
.B(n_3896),
.Y(n_7269)
);

BUFx3_ASAP7_75t_L g7270 ( 
.A(n_6538),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_6709),
.Y(n_7271)
);

INVx2_ASAP7_75t_L g7272 ( 
.A(n_6663),
.Y(n_7272)
);

INVx2_ASAP7_75t_L g7273 ( 
.A(n_6668),
.Y(n_7273)
);

NOR2xp33_ASAP7_75t_L g7274 ( 
.A(n_6864),
.B(n_3897),
.Y(n_7274)
);

INVx2_ASAP7_75t_L g7275 ( 
.A(n_6685),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_6712),
.Y(n_7276)
);

BUFx10_ASAP7_75t_L g7277 ( 
.A(n_6782),
.Y(n_7277)
);

OAI22xp5_ASAP7_75t_L g7278 ( 
.A1(n_6867),
.A2(n_3900),
.B1(n_3906),
.B2(n_3898),
.Y(n_7278)
);

OAI22xp33_ASAP7_75t_L g7279 ( 
.A1(n_6847),
.A2(n_3912),
.B1(n_3916),
.B2(n_3911),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_6855),
.B(n_4620),
.Y(n_7280)
);

INVx2_ASAP7_75t_L g7281 ( 
.A(n_6688),
.Y(n_7281)
);

CKINVDCx5p33_ASAP7_75t_R g7282 ( 
.A(n_6505),
.Y(n_7282)
);

BUFx2_ASAP7_75t_L g7283 ( 
.A(n_6492),
.Y(n_7283)
);

INVx1_ASAP7_75t_SL g7284 ( 
.A(n_6924),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6716),
.Y(n_7285)
);

OAI22xp33_ASAP7_75t_SL g7286 ( 
.A1(n_6833),
.A2(n_3868),
.B1(n_3870),
.B2(n_3864),
.Y(n_7286)
);

INVx4_ASAP7_75t_L g7287 ( 
.A(n_6926),
.Y(n_7287)
);

INVx2_ASAP7_75t_L g7288 ( 
.A(n_6689),
.Y(n_7288)
);

NAND2xp5_ASAP7_75t_L g7289 ( 
.A(n_6904),
.B(n_3919),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_SL g7290 ( 
.A(n_6925),
.B(n_3920),
.Y(n_7290)
);

OR2x6_ASAP7_75t_L g7291 ( 
.A(n_6919),
.B(n_6934),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_6719),
.Y(n_7292)
);

INVx1_ASAP7_75t_L g7293 ( 
.A(n_6658),
.Y(n_7293)
);

INVx2_ASAP7_75t_L g7294 ( 
.A(n_6697),
.Y(n_7294)
);

INVx2_ASAP7_75t_SL g7295 ( 
.A(n_6818),
.Y(n_7295)
);

INVx2_ASAP7_75t_SL g7296 ( 
.A(n_6834),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_6659),
.Y(n_7297)
);

NAND2xp5_ASAP7_75t_SL g7298 ( 
.A(n_6598),
.B(n_3922),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6661),
.Y(n_7299)
);

INVx2_ASAP7_75t_L g7300 ( 
.A(n_6700),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_SL g7301 ( 
.A(n_6808),
.B(n_6624),
.Y(n_7301)
);

BUFx2_ASAP7_75t_L g7302 ( 
.A(n_6526),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_SL g7303 ( 
.A(n_6624),
.B(n_3924),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6571),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_6620),
.Y(n_7305)
);

INVx2_ASAP7_75t_L g7306 ( 
.A(n_6628),
.Y(n_7306)
);

INVx2_ASAP7_75t_SL g7307 ( 
.A(n_6839),
.Y(n_7307)
);

BUFx6f_ASAP7_75t_L g7308 ( 
.A(n_6455),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_L g7309 ( 
.A(n_6792),
.B(n_3925),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_6637),
.Y(n_7310)
);

INVx5_ASAP7_75t_L g7311 ( 
.A(n_6926),
.Y(n_7311)
);

BUFx6f_ASAP7_75t_L g7312 ( 
.A(n_6455),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6672),
.Y(n_7313)
);

INVx1_ASAP7_75t_L g7314 ( 
.A(n_6690),
.Y(n_7314)
);

INVxp67_ASAP7_75t_L g7315 ( 
.A(n_6576),
.Y(n_7315)
);

OR2x6_ASAP7_75t_L g7316 ( 
.A(n_6932),
.B(n_3875),
.Y(n_7316)
);

NAND2xp33_ASAP7_75t_L g7317 ( 
.A(n_6861),
.B(n_3929),
.Y(n_7317)
);

BUFx6f_ASAP7_75t_L g7318 ( 
.A(n_6459),
.Y(n_7318)
);

OR2x2_ASAP7_75t_L g7319 ( 
.A(n_6537),
.B(n_6564),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_6665),
.Y(n_7320)
);

NAND2xp5_ASAP7_75t_SL g7321 ( 
.A(n_6941),
.B(n_3932),
.Y(n_7321)
);

INVx3_ASAP7_75t_L g7322 ( 
.A(n_6713),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_6815),
.Y(n_7323)
);

INVx2_ASAP7_75t_L g7324 ( 
.A(n_6667),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_SL g7325 ( 
.A(n_6923),
.B(n_3934),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_6669),
.Y(n_7326)
);

AOI22xp33_ASAP7_75t_L g7327 ( 
.A1(n_6670),
.A2(n_4614),
.B1(n_4649),
.B2(n_4605),
.Y(n_7327)
);

CKINVDCx16_ASAP7_75t_R g7328 ( 
.A(n_6641),
.Y(n_7328)
);

NAND2xp5_ASAP7_75t_SL g7329 ( 
.A(n_6923),
.B(n_3935),
.Y(n_7329)
);

BUFx10_ASAP7_75t_L g7330 ( 
.A(n_6946),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_6914),
.Y(n_7331)
);

INVx2_ASAP7_75t_L g7332 ( 
.A(n_6671),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_6795),
.B(n_3937),
.Y(n_7333)
);

INVx1_ASAP7_75t_SL g7334 ( 
.A(n_6693),
.Y(n_7334)
);

INVx2_ASAP7_75t_L g7335 ( 
.A(n_6673),
.Y(n_7335)
);

INVx3_ASAP7_75t_L g7336 ( 
.A(n_6735),
.Y(n_7336)
);

CKINVDCx5p33_ASAP7_75t_R g7337 ( 
.A(n_6932),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_6678),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6684),
.Y(n_7339)
);

OAI22xp5_ASAP7_75t_L g7340 ( 
.A1(n_6870),
.A2(n_3945),
.B1(n_3946),
.B2(n_3940),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6523),
.Y(n_7341)
);

NOR2xp33_ASAP7_75t_L g7342 ( 
.A(n_6734),
.B(n_3949),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6549),
.Y(n_7343)
);

AOI22xp33_ASAP7_75t_L g7344 ( 
.A1(n_6687),
.A2(n_4810),
.B1(n_4825),
.B2(n_4750),
.Y(n_7344)
);

INVx2_ASAP7_75t_L g7345 ( 
.A(n_6691),
.Y(n_7345)
);

NOR2xp33_ASAP7_75t_L g7346 ( 
.A(n_6943),
.B(n_6945),
.Y(n_7346)
);

INVx2_ASAP7_75t_L g7347 ( 
.A(n_6692),
.Y(n_7347)
);

NOR2xp33_ASAP7_75t_L g7348 ( 
.A(n_6947),
.B(n_3950),
.Y(n_7348)
);

INVx2_ASAP7_75t_L g7349 ( 
.A(n_6425),
.Y(n_7349)
);

INVx2_ASAP7_75t_L g7350 ( 
.A(n_6627),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_SL g7351 ( 
.A(n_6928),
.B(n_3954),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6790),
.Y(n_7352)
);

INVx3_ASAP7_75t_L g7353 ( 
.A(n_6735),
.Y(n_7353)
);

NAND2xp5_ASAP7_75t_L g7354 ( 
.A(n_6936),
.B(n_3955),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_6780),
.Y(n_7355)
);

BUFx6f_ASAP7_75t_L g7356 ( 
.A(n_6459),
.Y(n_7356)
);

OR2x2_ASAP7_75t_L g7357 ( 
.A(n_6567),
.B(n_6584),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_6559),
.Y(n_7358)
);

INVx3_ASAP7_75t_L g7359 ( 
.A(n_6742),
.Y(n_7359)
);

INVx2_ASAP7_75t_L g7360 ( 
.A(n_6527),
.Y(n_7360)
);

INVx2_ASAP7_75t_L g7361 ( 
.A(n_6474),
.Y(n_7361)
);

NAND2xp5_ASAP7_75t_L g7362 ( 
.A(n_6863),
.B(n_3956),
.Y(n_7362)
);

INVx2_ASAP7_75t_SL g7363 ( 
.A(n_6939),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6785),
.Y(n_7364)
);

BUFx10_ASAP7_75t_L g7365 ( 
.A(n_6957),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_6701),
.Y(n_7366)
);

BUFx6f_ASAP7_75t_L g7367 ( 
.A(n_6503),
.Y(n_7367)
);

INVx2_ASAP7_75t_L g7368 ( 
.A(n_6711),
.Y(n_7368)
);

INVx2_ASAP7_75t_L g7369 ( 
.A(n_6714),
.Y(n_7369)
);

NAND2xp5_ASAP7_75t_SL g7370 ( 
.A(n_6929),
.B(n_3958),
.Y(n_7370)
);

NAND2xp5_ASAP7_75t_L g7371 ( 
.A(n_6621),
.B(n_3967),
.Y(n_7371)
);

CKINVDCx5p33_ASAP7_75t_R g7372 ( 
.A(n_6935),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6718),
.Y(n_7373)
);

INVx2_ASAP7_75t_L g7374 ( 
.A(n_6725),
.Y(n_7374)
);

NOR2xp33_ASAP7_75t_L g7375 ( 
.A(n_6933),
.B(n_3969),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6786),
.Y(n_7376)
);

BUFx2_ASAP7_75t_L g7377 ( 
.A(n_6845),
.Y(n_7377)
);

OAI22xp33_ASAP7_75t_SL g7378 ( 
.A1(n_6409),
.A2(n_6918),
.B1(n_6842),
.B2(n_6840),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_6803),
.B(n_3970),
.Y(n_7379)
);

BUFx6f_ASAP7_75t_L g7380 ( 
.A(n_6503),
.Y(n_7380)
);

AND2x2_ASAP7_75t_L g7381 ( 
.A(n_6745),
.B(n_4620),
.Y(n_7381)
);

INVxp67_ASAP7_75t_SL g7382 ( 
.A(n_6592),
.Y(n_7382)
);

NAND2xp5_ASAP7_75t_SL g7383 ( 
.A(n_6944),
.B(n_3971),
.Y(n_7383)
);

NAND2xp5_ASAP7_75t_SL g7384 ( 
.A(n_6940),
.B(n_3972),
.Y(n_7384)
);

INVx3_ASAP7_75t_L g7385 ( 
.A(n_6742),
.Y(n_7385)
);

INVx3_ASAP7_75t_L g7386 ( 
.A(n_6744),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_6791),
.Y(n_7387)
);

AOI22xp33_ASAP7_75t_L g7388 ( 
.A1(n_6614),
.A2(n_6861),
.B1(n_6910),
.B2(n_6445),
.Y(n_7388)
);

INVx2_ASAP7_75t_L g7389 ( 
.A(n_6738),
.Y(n_7389)
);

INVx2_ASAP7_75t_L g7390 ( 
.A(n_6740),
.Y(n_7390)
);

INVx2_ASAP7_75t_L g7391 ( 
.A(n_6743),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_6754),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_6403),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_6577),
.B(n_3973),
.Y(n_7394)
);

INVx2_ASAP7_75t_SL g7395 ( 
.A(n_6513),
.Y(n_7395)
);

AND2x2_ASAP7_75t_L g7396 ( 
.A(n_6768),
.B(n_4661),
.Y(n_7396)
);

NAND2xp5_ASAP7_75t_L g7397 ( 
.A(n_6580),
.B(n_3974),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6404),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_6408),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6412),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_SL g7401 ( 
.A(n_6822),
.B(n_3977),
.Y(n_7401)
);

NOR2xp33_ASAP7_75t_L g7402 ( 
.A(n_6948),
.B(n_3979),
.Y(n_7402)
);

CKINVDCx5p33_ASAP7_75t_R g7403 ( 
.A(n_6935),
.Y(n_7403)
);

INVx2_ASAP7_75t_L g7404 ( 
.A(n_6755),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_6762),
.Y(n_7405)
);

NAND2xp33_ASAP7_75t_SL g7406 ( 
.A(n_6860),
.B(n_3981),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_SL g7407 ( 
.A(n_6814),
.B(n_3982),
.Y(n_7407)
);

OAI22xp33_ASAP7_75t_L g7408 ( 
.A1(n_6419),
.A2(n_3987),
.B1(n_3988),
.B2(n_3983),
.Y(n_7408)
);

INVx3_ASAP7_75t_L g7409 ( 
.A(n_6744),
.Y(n_7409)
);

AOI22xp5_ASAP7_75t_L g7410 ( 
.A1(n_6648),
.A2(n_3994),
.B1(n_3998),
.B2(n_3989),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6476),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_6481),
.Y(n_7412)
);

INVx1_ASAP7_75t_L g7413 ( 
.A(n_6485),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_6506),
.Y(n_7414)
);

NAND2xp5_ASAP7_75t_L g7415 ( 
.A(n_6548),
.B(n_4001),
.Y(n_7415)
);

BUFx2_ASAP7_75t_L g7416 ( 
.A(n_6787),
.Y(n_7416)
);

NAND2xp5_ASAP7_75t_SL g7417 ( 
.A(n_6953),
.B(n_6773),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6552),
.Y(n_7418)
);

INVxp67_ASAP7_75t_SL g7419 ( 
.A(n_6592),
.Y(n_7419)
);

AOI22xp33_ASAP7_75t_L g7420 ( 
.A1(n_6810),
.A2(n_3892),
.B1(n_3899),
.B2(n_3877),
.Y(n_7420)
);

INVx3_ASAP7_75t_L g7421 ( 
.A(n_6747),
.Y(n_7421)
);

INVx2_ASAP7_75t_SL g7422 ( 
.A(n_6513),
.Y(n_7422)
);

INVx3_ASAP7_75t_L g7423 ( 
.A(n_6747),
.Y(n_7423)
);

INVx2_ASAP7_75t_L g7424 ( 
.A(n_6763),
.Y(n_7424)
);

OR2x2_ASAP7_75t_L g7425 ( 
.A(n_6600),
.B(n_4005),
.Y(n_7425)
);

INVx2_ASAP7_75t_L g7426 ( 
.A(n_6769),
.Y(n_7426)
);

INVx2_ASAP7_75t_SL g7427 ( 
.A(n_6519),
.Y(n_7427)
);

INVx1_ASAP7_75t_L g7428 ( 
.A(n_6736),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_6760),
.Y(n_7429)
);

AOI22xp33_ASAP7_75t_L g7430 ( 
.A1(n_6810),
.A2(n_3909),
.B1(n_3917),
.B2(n_3901),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_6737),
.Y(n_7431)
);

INVx2_ASAP7_75t_L g7432 ( 
.A(n_6512),
.Y(n_7432)
);

INVx4_ASAP7_75t_L g7433 ( 
.A(n_6937),
.Y(n_7433)
);

NAND2xp5_ASAP7_75t_L g7434 ( 
.A(n_6781),
.B(n_4006),
.Y(n_7434)
);

BUFx2_ASAP7_75t_L g7435 ( 
.A(n_6608),
.Y(n_7435)
);

NOR2xp33_ASAP7_75t_L g7436 ( 
.A(n_6956),
.B(n_4008),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_6746),
.Y(n_7437)
);

NOR2xp33_ASAP7_75t_R g7438 ( 
.A(n_6676),
.B(n_4015),
.Y(n_7438)
);

NOR2xp33_ASAP7_75t_L g7439 ( 
.A(n_6496),
.B(n_4018),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6750),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_6753),
.Y(n_7441)
);

INVxp33_ASAP7_75t_SL g7442 ( 
.A(n_6424),
.Y(n_7442)
);

BUFx6f_ASAP7_75t_L g7443 ( 
.A(n_6519),
.Y(n_7443)
);

CKINVDCx11_ASAP7_75t_R g7444 ( 
.A(n_6894),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_SL g7445 ( 
.A(n_6902),
.B(n_4019),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6758),
.Y(n_7446)
);

NAND2xp5_ASAP7_75t_L g7447 ( 
.A(n_6930),
.B(n_4020),
.Y(n_7447)
);

INVx2_ASAP7_75t_SL g7448 ( 
.A(n_6539),
.Y(n_7448)
);

NAND3xp33_ASAP7_75t_L g7449 ( 
.A(n_6706),
.B(n_6451),
.C(n_6574),
.Y(n_7449)
);

INVx2_ASAP7_75t_L g7450 ( 
.A(n_6759),
.Y(n_7450)
);

NAND2xp5_ASAP7_75t_L g7451 ( 
.A(n_6800),
.B(n_4021),
.Y(n_7451)
);

INVx2_ASAP7_75t_SL g7452 ( 
.A(n_6539),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_L g7453 ( 
.A(n_6771),
.B(n_4022),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_6426),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_SL g7455 ( 
.A(n_6916),
.B(n_4023),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_6610),
.Y(n_7456)
);

INVx2_ASAP7_75t_L g7457 ( 
.A(n_6428),
.Y(n_7457)
);

INVx2_ASAP7_75t_SL g7458 ( 
.A(n_6569),
.Y(n_7458)
);

NAND3xp33_ASAP7_75t_L g7459 ( 
.A(n_6662),
.B(n_4029),
.C(n_4026),
.Y(n_7459)
);

NAND2xp5_ASAP7_75t_SL g7460 ( 
.A(n_6801),
.B(n_4031),
.Y(n_7460)
);

INVx2_ASAP7_75t_L g7461 ( 
.A(n_6448),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_6727),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6798),
.Y(n_7463)
);

INVx3_ASAP7_75t_L g7464 ( 
.A(n_6751),
.Y(n_7464)
);

INVx2_ASAP7_75t_L g7465 ( 
.A(n_6507),
.Y(n_7465)
);

INVx3_ASAP7_75t_L g7466 ( 
.A(n_6751),
.Y(n_7466)
);

CKINVDCx5p33_ASAP7_75t_R g7467 ( 
.A(n_6937),
.Y(n_7467)
);

CKINVDCx6p67_ASAP7_75t_R g7468 ( 
.A(n_6489),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_6797),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_6764),
.Y(n_7470)
);

INVxp67_ASAP7_75t_R g7471 ( 
.A(n_6909),
.Y(n_7471)
);

BUFx10_ASAP7_75t_L g7472 ( 
.A(n_6951),
.Y(n_7472)
);

BUFx6f_ASAP7_75t_L g7473 ( 
.A(n_6569),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6770),
.Y(n_7474)
);

BUFx6f_ASAP7_75t_L g7475 ( 
.A(n_6579),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_6774),
.Y(n_7476)
);

BUFx6f_ASAP7_75t_L g7477 ( 
.A(n_6579),
.Y(n_7477)
);

INVxp33_ASAP7_75t_L g7478 ( 
.A(n_6683),
.Y(n_7478)
);

INVx4_ASAP7_75t_SL g7479 ( 
.A(n_6810),
.Y(n_7479)
);

NOR2xp33_ASAP7_75t_L g7480 ( 
.A(n_6674),
.B(n_4036),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_6521),
.Y(n_7481)
);

INVx2_ASAP7_75t_L g7482 ( 
.A(n_6757),
.Y(n_7482)
);

OR2x6_ASAP7_75t_L g7483 ( 
.A(n_6951),
.B(n_3926),
.Y(n_7483)
);

INVx2_ASAP7_75t_L g7484 ( 
.A(n_6757),
.Y(n_7484)
);

INVx2_ASAP7_75t_L g7485 ( 
.A(n_6767),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_SL g7486 ( 
.A(n_6858),
.B(n_4037),
.Y(n_7486)
);

INVx5_ASAP7_75t_L g7487 ( 
.A(n_6826),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_6767),
.Y(n_7488)
);

INVx2_ASAP7_75t_L g7489 ( 
.A(n_6649),
.Y(n_7489)
);

INVx3_ASAP7_75t_L g7490 ( 
.A(n_6585),
.Y(n_7490)
);

NAND2xp5_ASAP7_75t_SL g7491 ( 
.A(n_6865),
.B(n_4039),
.Y(n_7491)
);

OR2x6_ASAP7_75t_L g7492 ( 
.A(n_6950),
.B(n_3931),
.Y(n_7492)
);

OAI22xp5_ASAP7_75t_L g7493 ( 
.A1(n_6866),
.A2(n_4041),
.B1(n_4042),
.B2(n_4040),
.Y(n_7493)
);

INVx1_ASAP7_75t_SL g7494 ( 
.A(n_6612),
.Y(n_7494)
);

NAND2xp5_ASAP7_75t_SL g7495 ( 
.A(n_6873),
.B(n_4043),
.Y(n_7495)
);

AND2x2_ASAP7_75t_L g7496 ( 
.A(n_6705),
.B(n_4661),
.Y(n_7496)
);

INVx2_ASAP7_75t_L g7497 ( 
.A(n_6555),
.Y(n_7497)
);

NAND3xp33_ASAP7_75t_L g7498 ( 
.A(n_6720),
.B(n_6723),
.C(n_6646),
.Y(n_7498)
);

INVx2_ASAP7_75t_L g7499 ( 
.A(n_6765),
.Y(n_7499)
);

AOI22xp33_ASAP7_75t_L g7500 ( 
.A1(n_6625),
.A2(n_3944),
.B1(n_3952),
.B2(n_3936),
.Y(n_7500)
);

INVx2_ASAP7_75t_L g7501 ( 
.A(n_6766),
.Y(n_7501)
);

OAI22xp33_ASAP7_75t_L g7502 ( 
.A1(n_6748),
.A2(n_4049),
.B1(n_4050),
.B2(n_4047),
.Y(n_7502)
);

INVx3_ASAP7_75t_L g7503 ( 
.A(n_6585),
.Y(n_7503)
);

INVx2_ASAP7_75t_L g7504 ( 
.A(n_6777),
.Y(n_7504)
);

INVx1_ASAP7_75t_L g7505 ( 
.A(n_6783),
.Y(n_7505)
);

NAND2xp33_ASAP7_75t_L g7506 ( 
.A(n_6817),
.B(n_4051),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_6784),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_6788),
.Y(n_7508)
);

INVx2_ASAP7_75t_L g7509 ( 
.A(n_6741),
.Y(n_7509)
);

INVx1_ASAP7_75t_L g7510 ( 
.A(n_6772),
.Y(n_7510)
);

NOR2xp33_ASAP7_75t_L g7511 ( 
.A(n_6832),
.B(n_4054),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_6959),
.Y(n_7512)
);

XNOR2xp5_ASAP7_75t_L g7513 ( 
.A(n_7215),
.B(n_6710),
.Y(n_7513)
);

AND2x6_ASAP7_75t_L g7514 ( 
.A(n_7393),
.B(n_6952),
.Y(n_7514)
);

CKINVDCx5p33_ASAP7_75t_R g7515 ( 
.A(n_7085),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_6967),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_6968),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_6974),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_6986),
.Y(n_7519)
);

AND2x2_ASAP7_75t_L g7520 ( 
.A(n_7125),
.B(n_6837),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_6997),
.Y(n_7521)
);

NOR2xp33_ASAP7_75t_SL g7522 ( 
.A(n_7141),
.B(n_6882),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7003),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7008),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7012),
.Y(n_7525)
);

OAI21xp5_ASAP7_75t_L g7526 ( 
.A1(n_7065),
.A2(n_6878),
.B(n_6836),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7018),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7019),
.Y(n_7528)
);

CKINVDCx20_ASAP7_75t_R g7529 ( 
.A(n_7112),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_7024),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7029),
.Y(n_7531)
);

XOR2xp5_ASAP7_75t_L g7532 ( 
.A(n_7282),
.B(n_6681),
.Y(n_7532)
);

INVx2_ASAP7_75t_L g7533 ( 
.A(n_7009),
.Y(n_7533)
);

INVx1_ASAP7_75t_L g7534 ( 
.A(n_7039),
.Y(n_7534)
);

INVxp67_ASAP7_75t_SL g7535 ( 
.A(n_7047),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_7070),
.B(n_6843),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7044),
.Y(n_7537)
);

INVxp33_ASAP7_75t_L g7538 ( 
.A(n_6980),
.Y(n_7538)
);

AND2x4_ASAP7_75t_L g7539 ( 
.A(n_7249),
.B(n_6881),
.Y(n_7539)
);

INVx2_ASAP7_75t_L g7540 ( 
.A(n_7013),
.Y(n_7540)
);

INVx2_ASAP7_75t_L g7541 ( 
.A(n_7014),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7056),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7059),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7060),
.Y(n_7544)
);

CKINVDCx16_ASAP7_75t_R g7545 ( 
.A(n_7328),
.Y(n_7545)
);

NAND2xp5_ASAP7_75t_L g7546 ( 
.A(n_7194),
.B(n_6775),
.Y(n_7546)
);

NOR2xp33_ASAP7_75t_SL g7547 ( 
.A(n_7163),
.B(n_6917),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7187),
.B(n_6844),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7064),
.Y(n_7549)
);

NOR2xp33_ASAP7_75t_L g7550 ( 
.A(n_6971),
.B(n_6739),
.Y(n_7550)
);

INVx2_ASAP7_75t_L g7551 ( 
.A(n_7017),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7072),
.Y(n_7552)
);

INVx1_ASAP7_75t_L g7553 ( 
.A(n_7074),
.Y(n_7553)
);

NOR2xp67_ASAP7_75t_L g7554 ( 
.A(n_7249),
.B(n_7311),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_7083),
.Y(n_7555)
);

INVx2_ASAP7_75t_L g7556 ( 
.A(n_7025),
.Y(n_7556)
);

BUFx5_ASAP7_75t_L g7557 ( 
.A(n_7323),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7093),
.Y(n_7558)
);

OR2x2_ASAP7_75t_L g7559 ( 
.A(n_7095),
.B(n_7284),
.Y(n_7559)
);

AOI21xp5_ASAP7_75t_L g7560 ( 
.A1(n_7079),
.A2(n_6660),
.B(n_6899),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7102),
.Y(n_7561)
);

AND2x4_ASAP7_75t_L g7562 ( 
.A(n_7311),
.B(n_6885),
.Y(n_7562)
);

INVx2_ASAP7_75t_L g7563 ( 
.A(n_7027),
.Y(n_7563)
);

NOR2x1_ASAP7_75t_L g7564 ( 
.A(n_6990),
.B(n_6851),
.Y(n_7564)
);

AND2x4_ASAP7_75t_L g7565 ( 
.A(n_6972),
.B(n_6749),
.Y(n_7565)
);

NOR2xp33_ASAP7_75t_SL g7566 ( 
.A(n_7337),
.B(n_6883),
.Y(n_7566)
);

INVx2_ASAP7_75t_L g7567 ( 
.A(n_7031),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7103),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_7104),
.Y(n_7569)
);

BUFx3_ASAP7_75t_L g7570 ( 
.A(n_7047),
.Y(n_7570)
);

AND2x2_ASAP7_75t_L g7571 ( 
.A(n_7230),
.B(n_6859),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7108),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7111),
.Y(n_7573)
);

NOR2xp67_ASAP7_75t_L g7574 ( 
.A(n_7487),
.B(n_6862),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7115),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7127),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7136),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_7138),
.Y(n_7578)
);

NAND2xp33_ASAP7_75t_R g7579 ( 
.A(n_7182),
.B(n_6874),
.Y(n_7579)
);

INVx2_ASAP7_75t_L g7580 ( 
.A(n_7032),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7037),
.Y(n_7581)
);

BUFx2_ASAP7_75t_L g7582 ( 
.A(n_6958),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7040),
.Y(n_7583)
);

CKINVDCx20_ASAP7_75t_R g7584 ( 
.A(n_7444),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7045),
.Y(n_7585)
);

OR2x2_ASAP7_75t_L g7586 ( 
.A(n_7319),
.B(n_6907),
.Y(n_7586)
);

AND2x2_ASAP7_75t_L g7587 ( 
.A(n_7280),
.B(n_6912),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_7052),
.Y(n_7588)
);

BUFx6f_ASAP7_75t_L g7589 ( 
.A(n_7099),
.Y(n_7589)
);

AND2x6_ASAP7_75t_L g7590 ( 
.A(n_7398),
.B(n_6848),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7062),
.Y(n_7591)
);

AND2x4_ASAP7_75t_L g7592 ( 
.A(n_6972),
.B(n_6589),
.Y(n_7592)
);

OR2x2_ASAP7_75t_SL g7593 ( 
.A(n_7449),
.B(n_7022),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_7075),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_7076),
.Y(n_7595)
);

INVxp67_ASAP7_75t_SL g7596 ( 
.A(n_7099),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_7078),
.Y(n_7597)
);

INVxp33_ASAP7_75t_L g7598 ( 
.A(n_6975),
.Y(n_7598)
);

NOR2xp67_ASAP7_75t_L g7599 ( 
.A(n_7487),
.B(n_6922),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_7080),
.Y(n_7600)
);

AND2x4_ASAP7_75t_L g7601 ( 
.A(n_7241),
.B(n_7287),
.Y(n_7601)
);

NOR2xp33_ASAP7_75t_L g7602 ( 
.A(n_7399),
.B(n_6805),
.Y(n_7602)
);

INVx2_ASAP7_75t_L g7603 ( 
.A(n_7084),
.Y(n_7603)
);

INVxp67_ASAP7_75t_L g7604 ( 
.A(n_7152),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_7090),
.Y(n_7605)
);

CKINVDCx5p33_ASAP7_75t_R g7606 ( 
.A(n_7372),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7092),
.Y(n_7607)
);

NAND2xp33_ASAP7_75t_R g7608 ( 
.A(n_7442),
.B(n_6852),
.Y(n_7608)
);

NOR2xp33_ASAP7_75t_L g7609 ( 
.A(n_7400),
.B(n_6589),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_7098),
.Y(n_7610)
);

INVxp33_ASAP7_75t_L g7611 ( 
.A(n_7357),
.Y(n_7611)
);

NOR2xp33_ASAP7_75t_L g7612 ( 
.A(n_7411),
.B(n_6911),
.Y(n_7612)
);

AND2x2_ASAP7_75t_L g7613 ( 
.A(n_7346),
.B(n_6841),
.Y(n_7613)
);

NOR2xp33_ASAP7_75t_L g7614 ( 
.A(n_7412),
.B(n_6854),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7109),
.Y(n_7615)
);

NOR2xp33_ASAP7_75t_L g7616 ( 
.A(n_7413),
.B(n_4055),
.Y(n_7616)
);

XNOR2xp5_ASAP7_75t_L g7617 ( 
.A(n_7049),
.B(n_4057),
.Y(n_7617)
);

AND2x2_ASAP7_75t_L g7618 ( 
.A(n_6983),
.B(n_4678),
.Y(n_7618)
);

INVx1_ASAP7_75t_SL g7619 ( 
.A(n_7091),
.Y(n_7619)
);

NOR2xp33_ASAP7_75t_L g7620 ( 
.A(n_7414),
.B(n_4061),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7114),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7119),
.Y(n_7622)
);

OR2x2_ASAP7_75t_L g7623 ( 
.A(n_6994),
.B(n_4068),
.Y(n_7623)
);

XOR2xp5_ASAP7_75t_L g7624 ( 
.A(n_7089),
.B(n_4069),
.Y(n_7624)
);

INVxp67_ASAP7_75t_L g7625 ( 
.A(n_7377),
.Y(n_7625)
);

AND2x2_ASAP7_75t_L g7626 ( 
.A(n_7081),
.B(n_4678),
.Y(n_7626)
);

NOR2xp67_ASAP7_75t_L g7627 ( 
.A(n_7433),
.B(n_4071),
.Y(n_7627)
);

NOR2xp33_ASAP7_75t_L g7628 ( 
.A(n_7418),
.B(n_4076),
.Y(n_7628)
);

OR2x6_ASAP7_75t_L g7629 ( 
.A(n_7015),
.B(n_6991),
.Y(n_7629)
);

INVx2_ASAP7_75t_L g7630 ( 
.A(n_7124),
.Y(n_7630)
);

BUFx6f_ASAP7_75t_L g7631 ( 
.A(n_7131),
.Y(n_7631)
);

CKINVDCx5p33_ASAP7_75t_R g7632 ( 
.A(n_7403),
.Y(n_7632)
);

XOR2xp5_ASAP7_75t_L g7633 ( 
.A(n_7219),
.B(n_4079),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7128),
.Y(n_7634)
);

XOR2xp5_ASAP7_75t_L g7635 ( 
.A(n_7467),
.B(n_4080),
.Y(n_7635)
);

CKINVDCx20_ASAP7_75t_R g7636 ( 
.A(n_7066),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7130),
.Y(n_7637)
);

CKINVDCx20_ASAP7_75t_R g7638 ( 
.A(n_7468),
.Y(n_7638)
);

INVx1_ASAP7_75t_L g7639 ( 
.A(n_7135),
.Y(n_7639)
);

AND2x4_ASAP7_75t_L g7640 ( 
.A(n_7110),
.B(n_3960),
.Y(n_7640)
);

AND2x2_ASAP7_75t_L g7641 ( 
.A(n_7033),
.B(n_4690),
.Y(n_7641)
);

AND2x2_ASAP7_75t_L g7642 ( 
.A(n_7046),
.B(n_7381),
.Y(n_7642)
);

INVx1_ASAP7_75t_L g7643 ( 
.A(n_7139),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_7320),
.Y(n_7644)
);

INVx1_ASAP7_75t_L g7645 ( 
.A(n_7246),
.Y(n_7645)
);

AND2x2_ASAP7_75t_L g7646 ( 
.A(n_7396),
.B(n_4690),
.Y(n_7646)
);

INVxp33_ASAP7_75t_SL g7647 ( 
.A(n_6962),
.Y(n_7647)
);

BUFx6f_ASAP7_75t_L g7648 ( 
.A(n_7131),
.Y(n_7648)
);

NAND2x1p5_ASAP7_75t_L g7649 ( 
.A(n_7166),
.B(n_3961),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7251),
.Y(n_7650)
);

NOR2xp33_ASAP7_75t_L g7651 ( 
.A(n_7236),
.B(n_4083),
.Y(n_7651)
);

INVx1_ASAP7_75t_L g7652 ( 
.A(n_7255),
.Y(n_7652)
);

INVxp67_ASAP7_75t_L g7653 ( 
.A(n_7416),
.Y(n_7653)
);

BUFx5_ASAP7_75t_L g7654 ( 
.A(n_7331),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7257),
.Y(n_7655)
);

CKINVDCx20_ASAP7_75t_R g7656 ( 
.A(n_7270),
.Y(n_7656)
);

NOR2xp33_ASAP7_75t_L g7657 ( 
.A(n_6996),
.B(n_7030),
.Y(n_7657)
);

BUFx2_ASAP7_75t_L g7658 ( 
.A(n_7283),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_7261),
.Y(n_7659)
);

OR2x2_ASAP7_75t_L g7660 ( 
.A(n_7302),
.B(n_4085),
.Y(n_7660)
);

XOR2x2_ASAP7_75t_L g7661 ( 
.A(n_7010),
.B(n_6998),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_SL g7662 ( 
.A(n_6970),
.B(n_4088),
.Y(n_7662)
);

CKINVDCx5p33_ASAP7_75t_R g7663 ( 
.A(n_7264),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7262),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7266),
.Y(n_7665)
);

INVx2_ASAP7_75t_L g7666 ( 
.A(n_7324),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_7271),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7276),
.Y(n_7668)
);

INVx2_ASAP7_75t_L g7669 ( 
.A(n_7326),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_7285),
.Y(n_7670)
);

OAI21xp5_ASAP7_75t_L g7671 ( 
.A1(n_7001),
.A2(n_3984),
.B(n_3962),
.Y(n_7671)
);

INVxp33_ASAP7_75t_L g7672 ( 
.A(n_7173),
.Y(n_7672)
);

INVx2_ASAP7_75t_L g7673 ( 
.A(n_7332),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_7292),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7335),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7188),
.Y(n_7676)
);

HB1xp67_ASAP7_75t_L g7677 ( 
.A(n_7011),
.Y(n_7677)
);

CKINVDCx20_ASAP7_75t_R g7678 ( 
.A(n_7205),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_7189),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7191),
.Y(n_7680)
);

NAND2x1p5_ASAP7_75t_L g7681 ( 
.A(n_7180),
.B(n_3991),
.Y(n_7681)
);

INVx2_ASAP7_75t_L g7682 ( 
.A(n_7338),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_7193),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_7038),
.B(n_4089),
.Y(n_7684)
);

AND2x2_ASAP7_75t_L g7685 ( 
.A(n_7048),
.B(n_7238),
.Y(n_7685)
);

NAND2xp5_ASAP7_75t_L g7686 ( 
.A(n_7087),
.B(n_4090),
.Y(n_7686)
);

INVx2_ASAP7_75t_L g7687 ( 
.A(n_7339),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7147),
.Y(n_7688)
);

XNOR2xp5_ASAP7_75t_L g7689 ( 
.A(n_7082),
.B(n_4092),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_7150),
.Y(n_7690)
);

INVx1_ASAP7_75t_L g7691 ( 
.A(n_7151),
.Y(n_7691)
);

XOR2x2_ASAP7_75t_L g7692 ( 
.A(n_7500),
.B(n_5),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_7153),
.Y(n_7693)
);

AND2x2_ASAP7_75t_L g7694 ( 
.A(n_7274),
.B(n_4826),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7345),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7155),
.Y(n_7696)
);

INVx4_ASAP7_75t_L g7697 ( 
.A(n_7173),
.Y(n_7697)
);

BUFx8_ASAP7_75t_L g7698 ( 
.A(n_6989),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7157),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7158),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_7160),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7347),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7164),
.Y(n_7703)
);

INVx4_ASAP7_75t_SL g7704 ( 
.A(n_7253),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7170),
.Y(n_7705)
);

INVx1_ASAP7_75t_L g7706 ( 
.A(n_7175),
.Y(n_7706)
);

CKINVDCx5p33_ASAP7_75t_R g7707 ( 
.A(n_7210),
.Y(n_7707)
);

INVx2_ASAP7_75t_SL g7708 ( 
.A(n_7472),
.Y(n_7708)
);

NOR2xp33_ASAP7_75t_L g7709 ( 
.A(n_7510),
.B(n_4095),
.Y(n_7709)
);

INVx1_ASAP7_75t_L g7710 ( 
.A(n_7304),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7428),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7196),
.Y(n_7712)
);

NAND2xp5_ASAP7_75t_L g7713 ( 
.A(n_7118),
.B(n_4100),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_7199),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_7207),
.Y(n_7715)
);

INVx1_ASAP7_75t_L g7716 ( 
.A(n_7216),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7221),
.Y(n_7717)
);

INVx3_ASAP7_75t_L g7718 ( 
.A(n_6991),
.Y(n_7718)
);

AND2x2_ASAP7_75t_L g7719 ( 
.A(n_7375),
.B(n_4826),
.Y(n_7719)
);

CKINVDCx5p33_ASAP7_75t_R g7720 ( 
.A(n_7210),
.Y(n_7720)
);

INVx1_ASAP7_75t_SL g7721 ( 
.A(n_7334),
.Y(n_7721)
);

BUFx6f_ASAP7_75t_SL g7722 ( 
.A(n_7123),
.Y(n_7722)
);

OR2x2_ASAP7_75t_L g7723 ( 
.A(n_7055),
.B(n_7362),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7225),
.Y(n_7724)
);

INVxp33_ASAP7_75t_L g7725 ( 
.A(n_7195),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_6961),
.Y(n_7726)
);

NOR2xp33_ASAP7_75t_L g7727 ( 
.A(n_7250),
.B(n_4103),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7228),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_7232),
.Y(n_7729)
);

NAND2xp33_ASAP7_75t_SL g7730 ( 
.A(n_7478),
.B(n_4112),
.Y(n_7730)
);

INVxp33_ASAP7_75t_L g7731 ( 
.A(n_7269),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7233),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7237),
.Y(n_7733)
);

NOR2xp33_ASAP7_75t_L g7734 ( 
.A(n_7036),
.B(n_4114),
.Y(n_7734)
);

INVx1_ASAP7_75t_L g7735 ( 
.A(n_6969),
.Y(n_7735)
);

CKINVDCx20_ASAP7_75t_R g7736 ( 
.A(n_7034),
.Y(n_7736)
);

AND2x2_ASAP7_75t_L g7737 ( 
.A(n_7315),
.B(n_4850),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_6978),
.Y(n_7738)
);

OR2x2_ASAP7_75t_L g7739 ( 
.A(n_7447),
.B(n_4117),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6981),
.Y(n_7740)
);

XOR2xp5_ASAP7_75t_L g7741 ( 
.A(n_7498),
.B(n_4119),
.Y(n_7741)
);

INVx1_ASAP7_75t_L g7742 ( 
.A(n_6985),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_6988),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_6995),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7007),
.Y(n_7745)
);

BUFx6f_ASAP7_75t_L g7746 ( 
.A(n_6993),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7145),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7148),
.Y(n_7748)
);

CKINVDCx20_ASAP7_75t_R g7749 ( 
.A(n_7143),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7463),
.Y(n_7750)
);

INVx1_ASAP7_75t_L g7751 ( 
.A(n_7176),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7178),
.Y(n_7752)
);

NAND2xp5_ASAP7_75t_L g7753 ( 
.A(n_7197),
.B(n_4120),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_7179),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7184),
.Y(n_7755)
);

XOR2xp5_ASAP7_75t_L g7756 ( 
.A(n_7459),
.B(n_4121),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7186),
.Y(n_7757)
);

AND2x2_ASAP7_75t_L g7758 ( 
.A(n_7069),
.B(n_4850),
.Y(n_7758)
);

NOR2xp67_ASAP7_75t_L g7759 ( 
.A(n_7042),
.B(n_4129),
.Y(n_7759)
);

AND2x2_ASAP7_75t_L g7760 ( 
.A(n_7348),
.B(n_4134),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7190),
.Y(n_7761)
);

INVx1_ASAP7_75t_L g7762 ( 
.A(n_7200),
.Y(n_7762)
);

CKINVDCx5p33_ASAP7_75t_R g7763 ( 
.A(n_7082),
.Y(n_7763)
);

NAND2xp33_ASAP7_75t_SL g7764 ( 
.A(n_7185),
.B(n_4135),
.Y(n_7764)
);

INVx1_ASAP7_75t_L g7765 ( 
.A(n_7202),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7203),
.Y(n_7766)
);

INVx1_ASAP7_75t_L g7767 ( 
.A(n_7206),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7209),
.Y(n_7768)
);

XOR2x2_ASAP7_75t_L g7769 ( 
.A(n_7436),
.B(n_5),
.Y(n_7769)
);

INVx1_ASAP7_75t_L g7770 ( 
.A(n_7211),
.Y(n_7770)
);

INVx2_ASAP7_75t_SL g7771 ( 
.A(n_7144),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7213),
.Y(n_7772)
);

INVx3_ASAP7_75t_L g7773 ( 
.A(n_6993),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_7220),
.Y(n_7774)
);

AND2x4_ASAP7_75t_L g7775 ( 
.A(n_7174),
.B(n_3996),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_7229),
.Y(n_7776)
);

BUFx2_ASAP7_75t_L g7777 ( 
.A(n_7435),
.Y(n_7777)
);

XOR2xp5_ASAP7_75t_L g7778 ( 
.A(n_7378),
.B(n_7071),
.Y(n_7778)
);

AND2x6_ASAP7_75t_L g7779 ( 
.A(n_7469),
.B(n_7293),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7234),
.Y(n_7780)
);

INVx1_ASAP7_75t_L g7781 ( 
.A(n_7235),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7240),
.Y(n_7782)
);

AND2x4_ASAP7_75t_L g7783 ( 
.A(n_7016),
.B(n_4000),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7243),
.Y(n_7784)
);

NOR2xp33_ASAP7_75t_L g7785 ( 
.A(n_7132),
.B(n_4139),
.Y(n_7785)
);

INVx1_ASAP7_75t_L g7786 ( 
.A(n_7244),
.Y(n_7786)
);

AOI21xp5_ASAP7_75t_L g7787 ( 
.A1(n_7358),
.A2(n_4004),
.B(n_4003),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7355),
.Y(n_7788)
);

AND2x2_ASAP7_75t_L g7789 ( 
.A(n_7402),
.B(n_4143),
.Y(n_7789)
);

CKINVDCx20_ASAP7_75t_R g7790 ( 
.A(n_7020),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_7364),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7376),
.Y(n_7792)
);

CKINVDCx5p33_ASAP7_75t_R g7793 ( 
.A(n_7020),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7387),
.Y(n_7794)
);

NAND2xp5_ASAP7_75t_L g7795 ( 
.A(n_7117),
.B(n_7154),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7470),
.Y(n_7796)
);

NOR2xp33_ASAP7_75t_SL g7797 ( 
.A(n_6992),
.B(n_4145),
.Y(n_7797)
);

NOR2xp33_ASAP7_75t_L g7798 ( 
.A(n_6977),
.B(n_4148),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7474),
.Y(n_7799)
);

OAI21xp5_ASAP7_75t_L g7800 ( 
.A1(n_7371),
.A2(n_4025),
.B(n_4016),
.Y(n_7800)
);

INVxp33_ASAP7_75t_L g7801 ( 
.A(n_7028),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_7297),
.Y(n_7802)
);

AND2x4_ASAP7_75t_L g7803 ( 
.A(n_7169),
.B(n_4030),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7299),
.Y(n_7804)
);

INVx2_ASAP7_75t_L g7805 ( 
.A(n_7247),
.Y(n_7805)
);

NOR2xp33_ASAP7_75t_L g7806 ( 
.A(n_7201),
.B(n_4149),
.Y(n_7806)
);

INVx1_ASAP7_75t_L g7807 ( 
.A(n_7352),
.Y(n_7807)
);

INVxp33_ASAP7_75t_L g7808 ( 
.A(n_7028),
.Y(n_7808)
);

XOR2x2_ASAP7_75t_L g7809 ( 
.A(n_6984),
.B(n_6),
.Y(n_7809)
);

CKINVDCx20_ASAP7_75t_R g7810 ( 
.A(n_7140),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_7504),
.Y(n_7811)
);

XNOR2xp5_ASAP7_75t_L g7812 ( 
.A(n_7000),
.B(n_4150),
.Y(n_7812)
);

CKINVDCx5p33_ASAP7_75t_R g7813 ( 
.A(n_7291),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_7507),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7260),
.Y(n_7815)
);

AND2x2_ASAP7_75t_L g7816 ( 
.A(n_7050),
.B(n_4152),
.Y(n_7816)
);

INVx1_ASAP7_75t_L g7817 ( 
.A(n_7267),
.Y(n_7817)
);

AND2x2_ASAP7_75t_L g7818 ( 
.A(n_7096),
.B(n_4154),
.Y(n_7818)
);

AND2x2_ASAP7_75t_L g7819 ( 
.A(n_7105),
.B(n_4155),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7268),
.Y(n_7820)
);

AND2x2_ASAP7_75t_L g7821 ( 
.A(n_7077),
.B(n_4156),
.Y(n_7821)
);

NAND2x1p5_ASAP7_75t_L g7822 ( 
.A(n_6966),
.B(n_4033),
.Y(n_7822)
);

NOR2xp33_ASAP7_75t_L g7823 ( 
.A(n_7156),
.B(n_7415),
.Y(n_7823)
);

NOR2xp33_ASAP7_75t_L g7824 ( 
.A(n_6960),
.B(n_4158),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_7272),
.Y(n_7825)
);

INVx1_ASAP7_75t_L g7826 ( 
.A(n_7273),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7275),
.Y(n_7827)
);

XNOR2xp5_ASAP7_75t_L g7828 ( 
.A(n_6965),
.B(n_4159),
.Y(n_7828)
);

INVx1_ASAP7_75t_L g7829 ( 
.A(n_7281),
.Y(n_7829)
);

NAND2xp5_ASAP7_75t_SL g7830 ( 
.A(n_6963),
.B(n_4163),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7288),
.Y(n_7831)
);

INVx1_ASAP7_75t_L g7832 ( 
.A(n_7294),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7300),
.Y(n_7833)
);

BUFx6f_ASAP7_75t_L g7834 ( 
.A(n_7185),
.Y(n_7834)
);

INVxp33_ASAP7_75t_L g7835 ( 
.A(n_7511),
.Y(n_7835)
);

CKINVDCx20_ASAP7_75t_R g7836 ( 
.A(n_7161),
.Y(n_7836)
);

NOR2xp33_ASAP7_75t_L g7837 ( 
.A(n_6964),
.B(n_4166),
.Y(n_7837)
);

AND2x2_ASAP7_75t_L g7838 ( 
.A(n_7198),
.B(n_4170),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7476),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7505),
.Y(n_7840)
);

INVx8_ASAP7_75t_L g7841 ( 
.A(n_7291),
.Y(n_7841)
);

INVx2_ASAP7_75t_L g7842 ( 
.A(n_7306),
.Y(n_7842)
);

XOR2xp5_ASAP7_75t_L g7843 ( 
.A(n_6982),
.B(n_4175),
.Y(n_7843)
);

INVx2_ASAP7_75t_L g7844 ( 
.A(n_7366),
.Y(n_7844)
);

AND2x4_ASAP7_75t_L g7845 ( 
.A(n_7295),
.B(n_4038),
.Y(n_7845)
);

INVx1_ASAP7_75t_L g7846 ( 
.A(n_7508),
.Y(n_7846)
);

NOR2xp67_ASAP7_75t_L g7847 ( 
.A(n_7208),
.B(n_4180),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7305),
.Y(n_7848)
);

INVx1_ASAP7_75t_L g7849 ( 
.A(n_7310),
.Y(n_7849)
);

NOR2xp33_ASAP7_75t_L g7850 ( 
.A(n_6979),
.B(n_4182),
.Y(n_7850)
);

INVx1_ASAP7_75t_L g7851 ( 
.A(n_7313),
.Y(n_7851)
);

BUFx6f_ASAP7_75t_L g7852 ( 
.A(n_7258),
.Y(n_7852)
);

CKINVDCx16_ASAP7_75t_R g7853 ( 
.A(n_7330),
.Y(n_7853)
);

AND2x2_ASAP7_75t_L g7854 ( 
.A(n_7212),
.B(n_4183),
.Y(n_7854)
);

INVx1_ASAP7_75t_L g7855 ( 
.A(n_7314),
.Y(n_7855)
);

CKINVDCx20_ASAP7_75t_R g7856 ( 
.A(n_7192),
.Y(n_7856)
);

INVx1_ASAP7_75t_L g7857 ( 
.A(n_7368),
.Y(n_7857)
);

BUFx6f_ASAP7_75t_L g7858 ( 
.A(n_7258),
.Y(n_7858)
);

NOR2xp33_ASAP7_75t_L g7859 ( 
.A(n_7023),
.B(n_4188),
.Y(n_7859)
);

NAND2xp5_ASAP7_75t_L g7860 ( 
.A(n_7035),
.B(n_4194),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7369),
.Y(n_7861)
);

INVx2_ASAP7_75t_SL g7862 ( 
.A(n_7308),
.Y(n_7862)
);

BUFx6f_ASAP7_75t_L g7863 ( 
.A(n_7308),
.Y(n_7863)
);

INVx1_ASAP7_75t_L g7864 ( 
.A(n_7373),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7374),
.Y(n_7865)
);

INVx1_ASAP7_75t_L g7866 ( 
.A(n_7389),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7390),
.Y(n_7867)
);

AND2x2_ASAP7_75t_L g7868 ( 
.A(n_7496),
.B(n_4203),
.Y(n_7868)
);

INVx2_ASAP7_75t_L g7869 ( 
.A(n_7391),
.Y(n_7869)
);

OR2x6_ASAP7_75t_L g7870 ( 
.A(n_7316),
.B(n_4048),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7392),
.Y(n_7871)
);

INVxp67_ASAP7_75t_SL g7872 ( 
.A(n_7312),
.Y(n_7872)
);

NAND2xp5_ASAP7_75t_L g7873 ( 
.A(n_7043),
.B(n_4204),
.Y(n_7873)
);

INVx2_ASAP7_75t_L g7874 ( 
.A(n_7404),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7405),
.Y(n_7875)
);

NOR2xp33_ASAP7_75t_L g7876 ( 
.A(n_7058),
.B(n_4206),
.Y(n_7876)
);

AND2x2_ASAP7_75t_L g7877 ( 
.A(n_7363),
.B(n_7439),
.Y(n_7877)
);

CKINVDCx20_ASAP7_75t_R g7878 ( 
.A(n_7263),
.Y(n_7878)
);

INVx1_ASAP7_75t_L g7879 ( 
.A(n_7424),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_7426),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7429),
.Y(n_7881)
);

AO21x1_ASAP7_75t_L g7882 ( 
.A1(n_7342),
.A2(n_4059),
.B(n_4053),
.Y(n_7882)
);

NOR2xp33_ASAP7_75t_SL g7883 ( 
.A(n_7002),
.B(n_4209),
.Y(n_7883)
);

INVx1_ASAP7_75t_L g7884 ( 
.A(n_7431),
.Y(n_7884)
);

INVx1_ASAP7_75t_L g7885 ( 
.A(n_7437),
.Y(n_7885)
);

AND2x2_ASAP7_75t_L g7886 ( 
.A(n_7316),
.B(n_4212),
.Y(n_7886)
);

INVx2_ASAP7_75t_SL g7887 ( 
.A(n_7312),
.Y(n_7887)
);

NOR2xp67_ASAP7_75t_L g7888 ( 
.A(n_7226),
.B(n_4213),
.Y(n_7888)
);

INVx1_ASAP7_75t_L g7889 ( 
.A(n_7440),
.Y(n_7889)
);

AND2x2_ASAP7_75t_L g7890 ( 
.A(n_7483),
.B(n_7086),
.Y(n_7890)
);

BUFx8_ASAP7_75t_L g7891 ( 
.A(n_7318),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_7441),
.Y(n_7892)
);

XOR2xp5_ASAP7_75t_L g7893 ( 
.A(n_7388),
.B(n_4215),
.Y(n_7893)
);

INVx1_ASAP7_75t_L g7894 ( 
.A(n_7446),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7394),
.B(n_4217),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_7450),
.Y(n_7896)
);

INVx1_ASAP7_75t_L g7897 ( 
.A(n_7122),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_7204),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_7341),
.Y(n_7899)
);

INVx1_ASAP7_75t_L g7900 ( 
.A(n_7343),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7223),
.Y(n_7901)
);

NAND2xp5_ASAP7_75t_L g7902 ( 
.A(n_7397),
.B(n_4218),
.Y(n_7902)
);

XOR2x2_ASAP7_75t_L g7903 ( 
.A(n_7480),
.B(n_6),
.Y(n_7903)
);

NAND2x1p5_ASAP7_75t_L g7904 ( 
.A(n_6976),
.B(n_4062),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7231),
.Y(n_7905)
);

OAI21xp5_ASAP7_75t_L g7906 ( 
.A1(n_7349),
.A2(n_4070),
.B(n_4066),
.Y(n_7906)
);

AOI21xp5_ASAP7_75t_L g7907 ( 
.A1(n_7350),
.A2(n_4074),
.B(n_4073),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7239),
.Y(n_7908)
);

NOR2xp33_ASAP7_75t_L g7909 ( 
.A(n_7453),
.B(n_4219),
.Y(n_7909)
);

BUFx2_ASAP7_75t_L g7910 ( 
.A(n_7318),
.Y(n_7910)
);

AND2x2_ASAP7_75t_L g7911 ( 
.A(n_7483),
.B(n_7088),
.Y(n_7911)
);

NAND2xp5_ASAP7_75t_L g7912 ( 
.A(n_7094),
.B(n_4221),
.Y(n_7912)
);

INVx1_ASAP7_75t_L g7913 ( 
.A(n_7289),
.Y(n_7913)
);

XOR2xp5_ASAP7_75t_L g7914 ( 
.A(n_7325),
.B(n_4222),
.Y(n_7914)
);

BUFx2_ASAP7_75t_L g7915 ( 
.A(n_7356),
.Y(n_7915)
);

AND2x2_ASAP7_75t_L g7916 ( 
.A(n_7365),
.B(n_4223),
.Y(n_7916)
);

INVxp33_ASAP7_75t_L g7917 ( 
.A(n_7356),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7137),
.Y(n_7918)
);

INVx1_ASAP7_75t_L g7919 ( 
.A(n_7142),
.Y(n_7919)
);

CKINVDCx5p33_ASAP7_75t_R g7920 ( 
.A(n_7438),
.Y(n_7920)
);

INVx1_ASAP7_75t_L g7921 ( 
.A(n_7126),
.Y(n_7921)
);

NOR2xp33_ASAP7_75t_SL g7922 ( 
.A(n_7494),
.B(n_4224),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7222),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7354),
.Y(n_7924)
);

INVx1_ASAP7_75t_L g7925 ( 
.A(n_7451),
.Y(n_7925)
);

INVx2_ASAP7_75t_L g7926 ( 
.A(n_7361),
.Y(n_7926)
);

INVx2_ASAP7_75t_L g7927 ( 
.A(n_7360),
.Y(n_7927)
);

XOR2xp5_ASAP7_75t_L g7928 ( 
.A(n_7329),
.B(n_4225),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_7301),
.Y(n_7929)
);

OR2x6_ASAP7_75t_L g7930 ( 
.A(n_7149),
.B(n_4077),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7454),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7457),
.Y(n_7932)
);

NOR2xp33_ASAP7_75t_L g7933 ( 
.A(n_7502),
.B(n_4228),
.Y(n_7933)
);

INVx2_ASAP7_75t_L g7934 ( 
.A(n_7432),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_7461),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_7465),
.Y(n_7936)
);

INVx1_ASAP7_75t_L g7937 ( 
.A(n_7481),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7497),
.Y(n_7938)
);

INVx1_ASAP7_75t_L g7939 ( 
.A(n_7509),
.Y(n_7939)
);

INVx1_ASAP7_75t_L g7940 ( 
.A(n_7309),
.Y(n_7940)
);

AND2x2_ASAP7_75t_L g7941 ( 
.A(n_7073),
.B(n_4229),
.Y(n_7941)
);

OR2x6_ASAP7_75t_L g7942 ( 
.A(n_7149),
.B(n_4081),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7333),
.Y(n_7943)
);

NOR2xp33_ASAP7_75t_L g7944 ( 
.A(n_7401),
.B(n_4231),
.Y(n_7944)
);

NAND2x1p5_ASAP7_75t_L g7945 ( 
.A(n_6987),
.B(n_4082),
.Y(n_7945)
);

AOI21x1_ASAP7_75t_L g7946 ( 
.A1(n_7489),
.A2(n_7321),
.B(n_7351),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7499),
.Y(n_7947)
);

XNOR2x2_ASAP7_75t_L g7948 ( 
.A(n_7218),
.B(n_4086),
.Y(n_7948)
);

BUFx6f_ASAP7_75t_L g7949 ( 
.A(n_7367),
.Y(n_7949)
);

INVx1_ASAP7_75t_L g7950 ( 
.A(n_7501),
.Y(n_7950)
);

AND2x2_ASAP7_75t_L g7951 ( 
.A(n_7134),
.B(n_4233),
.Y(n_7951)
);

NOR2xp33_ASAP7_75t_L g7952 ( 
.A(n_7445),
.B(n_4239),
.Y(n_7952)
);

XOR2x2_ASAP7_75t_L g7953 ( 
.A(n_7298),
.B(n_6),
.Y(n_7953)
);

INVx1_ASAP7_75t_L g7954 ( 
.A(n_7379),
.Y(n_7954)
);

INVx1_ASAP7_75t_L g7955 ( 
.A(n_7456),
.Y(n_7955)
);

NAND2xp5_ASAP7_75t_L g7956 ( 
.A(n_6973),
.B(n_4240),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_7462),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7482),
.Y(n_7958)
);

INVx1_ASAP7_75t_L g7959 ( 
.A(n_7484),
.Y(n_7959)
);

NAND2xp5_ASAP7_75t_L g7960 ( 
.A(n_7408),
.B(n_4242),
.Y(n_7960)
);

AND2x4_ASAP7_75t_L g7961 ( 
.A(n_7296),
.B(n_4091),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_7485),
.Y(n_7962)
);

CKINVDCx20_ASAP7_75t_R g7963 ( 
.A(n_7406),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7488),
.Y(n_7964)
);

NAND2xp5_ASAP7_75t_L g7965 ( 
.A(n_7327),
.B(n_4244),
.Y(n_7965)
);

NOR2xp33_ASAP7_75t_L g7966 ( 
.A(n_7455),
.B(n_4245),
.Y(n_7966)
);

AND2x2_ASAP7_75t_L g7967 ( 
.A(n_7242),
.B(n_4247),
.Y(n_7967)
);

INVx2_ASAP7_75t_L g7968 ( 
.A(n_6999),
.Y(n_7968)
);

INVx1_ASAP7_75t_L g7969 ( 
.A(n_7004),
.Y(n_7969)
);

XOR2xp5_ASAP7_75t_L g7970 ( 
.A(n_7370),
.B(n_7224),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_7004),
.Y(n_7971)
);

NAND2xp5_ASAP7_75t_L g7972 ( 
.A(n_7344),
.B(n_7004),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_7434),
.Y(n_7973)
);

BUFx6f_ASAP7_75t_L g7974 ( 
.A(n_7367),
.Y(n_7974)
);

XNOR2x2_ASAP7_75t_L g7975 ( 
.A(n_7410),
.B(n_4094),
.Y(n_7975)
);

NOR2xp33_ASAP7_75t_L g7976 ( 
.A(n_7101),
.B(n_4248),
.Y(n_7976)
);

AND2x2_ASAP7_75t_SL g7977 ( 
.A(n_7100),
.B(n_4097),
.Y(n_7977)
);

INVx1_ASAP7_75t_L g7978 ( 
.A(n_7417),
.Y(n_7978)
);

HB1xp67_ASAP7_75t_L g7979 ( 
.A(n_7380),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7384),
.Y(n_7980)
);

AND2x2_ASAP7_75t_L g7981 ( 
.A(n_7183),
.B(n_4249),
.Y(n_7981)
);

AND2x4_ASAP7_75t_L g7982 ( 
.A(n_7307),
.B(n_4107),
.Y(n_7982)
);

XOR2xp5_ASAP7_75t_L g7983 ( 
.A(n_7383),
.B(n_4253),
.Y(n_7983)
);

INVx2_ASAP7_75t_L g7984 ( 
.A(n_7006),
.Y(n_7984)
);

CKINVDCx20_ASAP7_75t_R g7985 ( 
.A(n_7277),
.Y(n_7985)
);

NOR2xp33_ASAP7_75t_L g7986 ( 
.A(n_7217),
.B(n_7425),
.Y(n_7986)
);

OAI21xp5_ASAP7_75t_L g7987 ( 
.A1(n_7133),
.A2(n_4118),
.B(n_4116),
.Y(n_7987)
);

INVx1_ASAP7_75t_L g7988 ( 
.A(n_7227),
.Y(n_7988)
);

AND2x2_ASAP7_75t_L g7989 ( 
.A(n_7063),
.B(n_7068),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7248),
.Y(n_7990)
);

INVx1_ASAP7_75t_L g7991 ( 
.A(n_7254),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7256),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_7290),
.Y(n_7993)
);

AND2x4_ASAP7_75t_L g7994 ( 
.A(n_7382),
.B(n_4122),
.Y(n_7994)
);

AND2x2_ASAP7_75t_L g7995 ( 
.A(n_7471),
.B(n_4263),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_7051),
.Y(n_7996)
);

AND2x2_ASAP7_75t_L g7997 ( 
.A(n_7067),
.B(n_4264),
.Y(n_7997)
);

BUFx3_ASAP7_75t_L g7998 ( 
.A(n_7380),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_7097),
.Y(n_7999)
);

AND2x2_ASAP7_75t_L g8000 ( 
.A(n_7177),
.B(n_4265),
.Y(n_8000)
);

HB1xp67_ASAP7_75t_L g8001 ( 
.A(n_7443),
.Y(n_8001)
);

XNOR2xp5_ASAP7_75t_L g8002 ( 
.A(n_7005),
.B(n_7407),
.Y(n_8002)
);

INVx1_ASAP7_75t_L g8003 ( 
.A(n_7107),
.Y(n_8003)
);

XOR2xp5_ASAP7_75t_L g8004 ( 
.A(n_7303),
.B(n_7486),
.Y(n_8004)
);

CKINVDCx20_ASAP7_75t_R g8005 ( 
.A(n_7479),
.Y(n_8005)
);

NOR2xp33_ASAP7_75t_L g8006 ( 
.A(n_7252),
.B(n_4270),
.Y(n_8006)
);

OAI21xp5_ASAP7_75t_L g8007 ( 
.A1(n_7165),
.A2(n_4128),
.B(n_4126),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_7113),
.Y(n_8008)
);

BUFx3_ASAP7_75t_L g8009 ( 
.A(n_7443),
.Y(n_8009)
);

INVx1_ASAP7_75t_L g8010 ( 
.A(n_7121),
.Y(n_8010)
);

INVx1_ASAP7_75t_L g8011 ( 
.A(n_7419),
.Y(n_8011)
);

AND2x2_ASAP7_75t_L g8012 ( 
.A(n_7177),
.B(n_4271),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_7021),
.Y(n_8013)
);

INVx2_ASAP7_75t_SL g8014 ( 
.A(n_7473),
.Y(n_8014)
);

OR2x6_ASAP7_75t_L g8015 ( 
.A(n_7473),
.B(n_4142),
.Y(n_8015)
);

NAND2xp5_ASAP7_75t_L g8016 ( 
.A(n_7041),
.B(n_4273),
.Y(n_8016)
);

INVxp33_ASAP7_75t_L g8017 ( 
.A(n_7475),
.Y(n_8017)
);

CKINVDCx20_ASAP7_75t_R g8018 ( 
.A(n_7475),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7026),
.Y(n_8019)
);

INVx1_ASAP7_75t_L g8020 ( 
.A(n_7053),
.Y(n_8020)
);

INVx1_ASAP7_75t_L g8021 ( 
.A(n_7512),
.Y(n_8021)
);

NAND2xp5_ASAP7_75t_L g8022 ( 
.A(n_7685),
.B(n_7286),
.Y(n_8022)
);

INVx2_ASAP7_75t_L g8023 ( 
.A(n_7516),
.Y(n_8023)
);

NAND2xp5_ASAP7_75t_SL g8024 ( 
.A(n_7731),
.B(n_7477),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7517),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7518),
.Y(n_8026)
);

AOI22xp5_ASAP7_75t_SL g8027 ( 
.A1(n_7812),
.A2(n_7116),
.B1(n_7106),
.B2(n_7278),
.Y(n_8027)
);

INVx2_ASAP7_75t_SL g8028 ( 
.A(n_7891),
.Y(n_8028)
);

NAND2xp5_ASAP7_75t_L g8029 ( 
.A(n_7823),
.B(n_7168),
.Y(n_8029)
);

INVx2_ASAP7_75t_L g8030 ( 
.A(n_7519),
.Y(n_8030)
);

NAND2xp5_ASAP7_75t_SL g8031 ( 
.A(n_7538),
.B(n_7835),
.Y(n_8031)
);

NOR2xp33_ASAP7_75t_L g8032 ( 
.A(n_7647),
.B(n_7171),
.Y(n_8032)
);

NAND2xp5_ASAP7_75t_SL g8033 ( 
.A(n_7723),
.B(n_7477),
.Y(n_8033)
);

BUFx3_ASAP7_75t_L g8034 ( 
.A(n_7790),
.Y(n_8034)
);

AOI221xp5_ASAP7_75t_L g8035 ( 
.A1(n_7657),
.A2(n_7651),
.B1(n_8006),
.B2(n_7976),
.C(n_7734),
.Y(n_8035)
);

NOR2xp33_ASAP7_75t_L g8036 ( 
.A(n_7727),
.B(n_7172),
.Y(n_8036)
);

AND2x2_ASAP7_75t_L g8037 ( 
.A(n_7694),
.B(n_7057),
.Y(n_8037)
);

NOR2xp33_ASAP7_75t_L g8038 ( 
.A(n_7925),
.B(n_7279),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_SL g8039 ( 
.A(n_7598),
.B(n_7054),
.Y(n_8039)
);

INVx2_ASAP7_75t_L g8040 ( 
.A(n_7521),
.Y(n_8040)
);

BUFx2_ASAP7_75t_L g8041 ( 
.A(n_8018),
.Y(n_8041)
);

NAND2xp5_ASAP7_75t_L g8042 ( 
.A(n_7795),
.B(n_7495),
.Y(n_8042)
);

NAND2xp5_ASAP7_75t_SL g8043 ( 
.A(n_7877),
.B(n_7061),
.Y(n_8043)
);

AOI22xp5_ASAP7_75t_L g8044 ( 
.A1(n_7661),
.A2(n_7506),
.B1(n_7317),
.B2(n_7460),
.Y(n_8044)
);

NAND2x1p5_ASAP7_75t_L g8045 ( 
.A(n_7554),
.B(n_7120),
.Y(n_8045)
);

INVx1_ASAP7_75t_L g8046 ( 
.A(n_7523),
.Y(n_8046)
);

INVx2_ASAP7_75t_L g8047 ( 
.A(n_7524),
.Y(n_8047)
);

O2A1O1Ixp33_ASAP7_75t_L g8048 ( 
.A1(n_7800),
.A2(n_7493),
.B(n_7491),
.C(n_7340),
.Y(n_8048)
);

INVx2_ASAP7_75t_L g8049 ( 
.A(n_7525),
.Y(n_8049)
);

INVx2_ASAP7_75t_L g8050 ( 
.A(n_7527),
.Y(n_8050)
);

INVx8_ASAP7_75t_L g8051 ( 
.A(n_7629),
.Y(n_8051)
);

INVx2_ASAP7_75t_L g8052 ( 
.A(n_7528),
.Y(n_8052)
);

INVxp67_ASAP7_75t_SL g8053 ( 
.A(n_7677),
.Y(n_8053)
);

INVx1_ASAP7_75t_L g8054 ( 
.A(n_7530),
.Y(n_8054)
);

HB1xp67_ASAP7_75t_L g8055 ( 
.A(n_7658),
.Y(n_8055)
);

OR2x6_ASAP7_75t_L g8056 ( 
.A(n_7841),
.B(n_7395),
.Y(n_8056)
);

CKINVDCx20_ASAP7_75t_R g8057 ( 
.A(n_7529),
.Y(n_8057)
);

NAND2xp5_ASAP7_75t_L g8058 ( 
.A(n_7918),
.B(n_7420),
.Y(n_8058)
);

NAND2xp5_ASAP7_75t_L g8059 ( 
.A(n_7919),
.B(n_7430),
.Y(n_8059)
);

NAND2xp5_ASAP7_75t_L g8060 ( 
.A(n_7940),
.B(n_7129),
.Y(n_8060)
);

NAND2xp5_ASAP7_75t_L g8061 ( 
.A(n_7943),
.B(n_7159),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_SL g8062 ( 
.A(n_7642),
.B(n_7162),
.Y(n_8062)
);

NAND2xp5_ASAP7_75t_L g8063 ( 
.A(n_7954),
.B(n_7167),
.Y(n_8063)
);

AND2x2_ASAP7_75t_L g8064 ( 
.A(n_7719),
.B(n_7492),
.Y(n_8064)
);

INVx2_ASAP7_75t_L g8065 ( 
.A(n_7531),
.Y(n_8065)
);

AOI22xp5_ASAP7_75t_L g8066 ( 
.A1(n_7986),
.A2(n_7492),
.B1(n_7181),
.B2(n_7259),
.Y(n_8066)
);

NOR2xp33_ASAP7_75t_L g8067 ( 
.A(n_7611),
.B(n_7245),
.Y(n_8067)
);

INVx2_ASAP7_75t_L g8068 ( 
.A(n_7534),
.Y(n_8068)
);

NOR2xp33_ASAP7_75t_L g8069 ( 
.A(n_7798),
.B(n_7265),
.Y(n_8069)
);

INVx1_ASAP7_75t_L g8070 ( 
.A(n_7537),
.Y(n_8070)
);

AOI22xp33_ASAP7_75t_L g8071 ( 
.A1(n_7933),
.A2(n_7336),
.B1(n_7353),
.B2(n_7322),
.Y(n_8071)
);

NOR2xp33_ASAP7_75t_L g8072 ( 
.A(n_7686),
.B(n_7359),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_L g8073 ( 
.A(n_7546),
.B(n_7385),
.Y(n_8073)
);

HB1xp67_ASAP7_75t_L g8074 ( 
.A(n_7582),
.Y(n_8074)
);

NOR2xp33_ASAP7_75t_L g8075 ( 
.A(n_7973),
.B(n_7386),
.Y(n_8075)
);

AND2x2_ASAP7_75t_L g8076 ( 
.A(n_7520),
.B(n_7409),
.Y(n_8076)
);

INVx2_ASAP7_75t_L g8077 ( 
.A(n_7542),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7543),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7544),
.Y(n_8079)
);

AND2x2_ASAP7_75t_L g8080 ( 
.A(n_7548),
.B(n_7421),
.Y(n_8080)
);

OAI22xp33_ASAP7_75t_L g8081 ( 
.A1(n_7797),
.A2(n_7423),
.B1(n_7466),
.B2(n_7464),
.Y(n_8081)
);

NAND2xp5_ASAP7_75t_L g8082 ( 
.A(n_7785),
.B(n_7490),
.Y(n_8082)
);

NOR2xp33_ASAP7_75t_L g8083 ( 
.A(n_7806),
.B(n_7503),
.Y(n_8083)
);

AOI22xp5_ASAP7_75t_L g8084 ( 
.A1(n_7890),
.A2(n_7427),
.B1(n_7448),
.B2(n_7422),
.Y(n_8084)
);

NAND2xp5_ASAP7_75t_L g8085 ( 
.A(n_7909),
.B(n_7452),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_7549),
.Y(n_8086)
);

NAND2xp5_ASAP7_75t_L g8087 ( 
.A(n_7901),
.B(n_7458),
.Y(n_8087)
);

AOI22xp33_ASAP7_75t_L g8088 ( 
.A1(n_7617),
.A2(n_7214),
.B1(n_7146),
.B2(n_4151),
.Y(n_8088)
);

HB1xp67_ASAP7_75t_L g8089 ( 
.A(n_7777),
.Y(n_8089)
);

NAND2xp5_ASAP7_75t_SL g8090 ( 
.A(n_7612),
.B(n_4277),
.Y(n_8090)
);

INVx2_ASAP7_75t_SL g8091 ( 
.A(n_7629),
.Y(n_8091)
);

NOR2xp33_ASAP7_75t_SL g8092 ( 
.A(n_7515),
.B(n_7606),
.Y(n_8092)
);

INVx2_ASAP7_75t_L g8093 ( 
.A(n_7552),
.Y(n_8093)
);

NAND2xp5_ASAP7_75t_L g8094 ( 
.A(n_7905),
.B(n_4144),
.Y(n_8094)
);

AOI21xp5_ASAP7_75t_L g8095 ( 
.A1(n_7526),
.A2(n_4164),
.B(n_4162),
.Y(n_8095)
);

AOI22xp33_ASAP7_75t_L g8096 ( 
.A1(n_7893),
.A2(n_4176),
.B1(n_4179),
.B2(n_4169),
.Y(n_8096)
);

INVx2_ASAP7_75t_SL g8097 ( 
.A(n_7793),
.Y(n_8097)
);

NAND2xp5_ASAP7_75t_L g8098 ( 
.A(n_7908),
.B(n_4184),
.Y(n_8098)
);

NAND3xp33_ASAP7_75t_L g8099 ( 
.A(n_7824),
.B(n_4283),
.C(n_4281),
.Y(n_8099)
);

NOR2xp33_ASAP7_75t_L g8100 ( 
.A(n_7559),
.B(n_4284),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_L g8101 ( 
.A(n_7913),
.B(n_4185),
.Y(n_8101)
);

NAND2xp5_ASAP7_75t_L g8102 ( 
.A(n_7837),
.B(n_4186),
.Y(n_8102)
);

NAND2xp5_ASAP7_75t_SL g8103 ( 
.A(n_7602),
.B(n_4286),
.Y(n_8103)
);

O2A1O1Ixp33_ASAP7_75t_L g8104 ( 
.A1(n_7960),
.A2(n_4191),
.B(n_4192),
.C(n_4189),
.Y(n_8104)
);

INVx1_ASAP7_75t_L g8105 ( 
.A(n_7553),
.Y(n_8105)
);

INVx2_ASAP7_75t_SL g8106 ( 
.A(n_7592),
.Y(n_8106)
);

INVx1_ASAP7_75t_L g8107 ( 
.A(n_7555),
.Y(n_8107)
);

INVxp67_ASAP7_75t_L g8108 ( 
.A(n_7721),
.Y(n_8108)
);

NOR2xp33_ASAP7_75t_L g8109 ( 
.A(n_7850),
.B(n_4287),
.Y(n_8109)
);

NAND2x1p5_ASAP7_75t_L g8110 ( 
.A(n_7697),
.B(n_4193),
.Y(n_8110)
);

NAND2xp5_ASAP7_75t_L g8111 ( 
.A(n_7859),
.B(n_4195),
.Y(n_8111)
);

NAND2xp5_ASAP7_75t_L g8112 ( 
.A(n_7876),
.B(n_4197),
.Y(n_8112)
);

NOR2xp33_ASAP7_75t_L g8113 ( 
.A(n_7653),
.B(n_4291),
.Y(n_8113)
);

INVx2_ASAP7_75t_L g8114 ( 
.A(n_7558),
.Y(n_8114)
);

NAND2xp5_ASAP7_75t_L g8115 ( 
.A(n_7684),
.B(n_4200),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7561),
.Y(n_8116)
);

NAND2xp5_ASAP7_75t_L g8117 ( 
.A(n_7571),
.B(n_4205),
.Y(n_8117)
);

NAND2xp5_ASAP7_75t_SL g8118 ( 
.A(n_7536),
.B(n_4293),
.Y(n_8118)
);

INVx2_ASAP7_75t_L g8119 ( 
.A(n_7568),
.Y(n_8119)
);

INVx2_ASAP7_75t_L g8120 ( 
.A(n_7569),
.Y(n_8120)
);

NOR2xp33_ASAP7_75t_L g8121 ( 
.A(n_7619),
.B(n_4295),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_7572),
.Y(n_8122)
);

NAND2xp5_ASAP7_75t_L g8123 ( 
.A(n_7616),
.B(n_4207),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_SL g8124 ( 
.A(n_7609),
.B(n_4296),
.Y(n_8124)
);

NAND2xp5_ASAP7_75t_L g8125 ( 
.A(n_7620),
.B(n_4216),
.Y(n_8125)
);

NAND2xp5_ASAP7_75t_L g8126 ( 
.A(n_7628),
.B(n_4227),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_7789),
.B(n_4232),
.Y(n_8127)
);

NAND3xp33_ASAP7_75t_L g8128 ( 
.A(n_7671),
.B(n_4298),
.C(n_4297),
.Y(n_8128)
);

BUFx6f_ASAP7_75t_L g8129 ( 
.A(n_7589),
.Y(n_8129)
);

NAND2xp5_ASAP7_75t_SL g8130 ( 
.A(n_7550),
.B(n_4299),
.Y(n_8130)
);

INVx2_ASAP7_75t_L g8131 ( 
.A(n_7573),
.Y(n_8131)
);

NAND2xp5_ASAP7_75t_L g8132 ( 
.A(n_7760),
.B(n_4236),
.Y(n_8132)
);

NAND2xp5_ASAP7_75t_L g8133 ( 
.A(n_7821),
.B(n_4243),
.Y(n_8133)
);

NAND2xp5_ASAP7_75t_L g8134 ( 
.A(n_7838),
.B(n_4266),
.Y(n_8134)
);

CKINVDCx5p33_ASAP7_75t_R g8135 ( 
.A(n_7632),
.Y(n_8135)
);

AND2x2_ASAP7_75t_L g8136 ( 
.A(n_7868),
.B(n_4300),
.Y(n_8136)
);

NOR2xp33_ASAP7_75t_L g8137 ( 
.A(n_7604),
.B(n_4301),
.Y(n_8137)
);

NOR2xp67_ASAP7_75t_L g8138 ( 
.A(n_7625),
.B(n_7),
.Y(n_8138)
);

BUFx3_ASAP7_75t_L g8139 ( 
.A(n_7656),
.Y(n_8139)
);

NOR2xp33_ASAP7_75t_L g8140 ( 
.A(n_7725),
.B(n_4302),
.Y(n_8140)
);

NAND2xp5_ASAP7_75t_SL g8141 ( 
.A(n_7911),
.B(n_4303),
.Y(n_8141)
);

AOI221xp5_ASAP7_75t_L g8142 ( 
.A1(n_7741),
.A2(n_4279),
.B1(n_4285),
.B2(n_4276),
.C(n_4267),
.Y(n_8142)
);

NAND2xp5_ASAP7_75t_L g8143 ( 
.A(n_7854),
.B(n_4292),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_7575),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7576),
.Y(n_8145)
);

NAND2xp5_ASAP7_75t_L g8146 ( 
.A(n_7613),
.B(n_4311),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_7577),
.Y(n_8147)
);

NAND2xp5_ASAP7_75t_SL g8148 ( 
.A(n_7922),
.B(n_4306),
.Y(n_8148)
);

INVx2_ASAP7_75t_L g8149 ( 
.A(n_7578),
.Y(n_8149)
);

NAND2xp5_ASAP7_75t_L g8150 ( 
.A(n_7709),
.B(n_7713),
.Y(n_8150)
);

NAND2xp5_ASAP7_75t_L g8151 ( 
.A(n_7614),
.B(n_4313),
.Y(n_8151)
);

AOI22xp5_ASAP7_75t_L g8152 ( 
.A1(n_7970),
.A2(n_4309),
.B1(n_4310),
.B2(n_4308),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7645),
.Y(n_8153)
);

INVx1_ASAP7_75t_SL g8154 ( 
.A(n_7736),
.Y(n_8154)
);

NOR2xp33_ASAP7_75t_SL g8155 ( 
.A(n_7836),
.B(n_7856),
.Y(n_8155)
);

NAND2xp5_ASAP7_75t_L g8156 ( 
.A(n_7753),
.B(n_4318),
.Y(n_8156)
);

OR2x2_ASAP7_75t_L g8157 ( 
.A(n_7660),
.B(n_4312),
.Y(n_8157)
);

HB1xp67_ASAP7_75t_L g8158 ( 
.A(n_7746),
.Y(n_8158)
);

NOR2xp33_ASAP7_75t_SL g8159 ( 
.A(n_7678),
.B(n_4315),
.Y(n_8159)
);

AND2x2_ASAP7_75t_L g8160 ( 
.A(n_7818),
.B(n_4317),
.Y(n_8160)
);

OAI22xp5_ASAP7_75t_SL g8161 ( 
.A1(n_8002),
.A2(n_4320),
.B1(n_4321),
.B2(n_4319),
.Y(n_8161)
);

NOR2xp33_ASAP7_75t_L g8162 ( 
.A(n_7895),
.B(n_4322),
.Y(n_8162)
);

INVx1_ASAP7_75t_L g8163 ( 
.A(n_7650),
.Y(n_8163)
);

AOI22xp5_ASAP7_75t_L g8164 ( 
.A1(n_7778),
.A2(n_7579),
.B1(n_7587),
.B2(n_7995),
.Y(n_8164)
);

NAND2xp5_ASAP7_75t_L g8165 ( 
.A(n_7860),
.B(n_4328),
.Y(n_8165)
);

NOR2xp33_ASAP7_75t_L g8166 ( 
.A(n_7902),
.B(n_4323),
.Y(n_8166)
);

AND2x6_ASAP7_75t_SL g8167 ( 
.A(n_8015),
.B(n_4337),
.Y(n_8167)
);

NAND2xp5_ASAP7_75t_L g8168 ( 
.A(n_7873),
.B(n_7912),
.Y(n_8168)
);

NOR2xp33_ASAP7_75t_L g8169 ( 
.A(n_7586),
.B(n_4324),
.Y(n_8169)
);

INVx4_ASAP7_75t_L g8170 ( 
.A(n_7746),
.Y(n_8170)
);

NAND2xp33_ASAP7_75t_L g8171 ( 
.A(n_7779),
.B(n_4325),
.Y(n_8171)
);

INVx1_ASAP7_75t_SL g8172 ( 
.A(n_7749),
.Y(n_8172)
);

NAND2xp5_ASAP7_75t_L g8173 ( 
.A(n_7924),
.B(n_4344),
.Y(n_8173)
);

NAND2xp5_ASAP7_75t_L g8174 ( 
.A(n_7898),
.B(n_4351),
.Y(n_8174)
);

NAND2xp5_ASAP7_75t_L g8175 ( 
.A(n_7652),
.B(n_4354),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_L g8176 ( 
.A(n_7655),
.B(n_4355),
.Y(n_8176)
);

NAND2xp5_ASAP7_75t_L g8177 ( 
.A(n_7659),
.B(n_7664),
.Y(n_8177)
);

OAI22xp5_ASAP7_75t_L g8178 ( 
.A1(n_7593),
.A2(n_7667),
.B1(n_7668),
.B2(n_7665),
.Y(n_8178)
);

OAI21xp5_ASAP7_75t_L g8179 ( 
.A1(n_7906),
.A2(n_4364),
.B(n_4356),
.Y(n_8179)
);

INVx4_ASAP7_75t_L g8180 ( 
.A(n_7589),
.Y(n_8180)
);

INVx3_ASAP7_75t_L g8181 ( 
.A(n_7601),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7670),
.Y(n_8182)
);

OR2x2_ASAP7_75t_L g8183 ( 
.A(n_7739),
.B(n_7623),
.Y(n_8183)
);

INVx2_ASAP7_75t_L g8184 ( 
.A(n_7674),
.Y(n_8184)
);

BUFx6f_ASAP7_75t_L g8185 ( 
.A(n_7631),
.Y(n_8185)
);

OAI22xp5_ASAP7_75t_L g8186 ( 
.A1(n_7676),
.A2(n_4332),
.B1(n_4334),
.B2(n_4327),
.Y(n_8186)
);

NAND2xp5_ASAP7_75t_L g8187 ( 
.A(n_7560),
.B(n_7710),
.Y(n_8187)
);

OAI221xp5_ASAP7_75t_L g8188 ( 
.A1(n_7952),
.A2(n_4394),
.B1(n_4401),
.B2(n_4375),
.C(n_4374),
.Y(n_8188)
);

NAND2xp5_ASAP7_75t_L g8189 ( 
.A(n_7711),
.B(n_4405),
.Y(n_8189)
);

A2O1A1Ixp33_ASAP7_75t_L g8190 ( 
.A1(n_7847),
.A2(n_4421),
.B(n_4429),
.C(n_4415),
.Y(n_8190)
);

NAND2xp5_ASAP7_75t_L g8191 ( 
.A(n_7788),
.B(n_4432),
.Y(n_8191)
);

OAI21xp33_ASAP7_75t_L g8192 ( 
.A1(n_7903),
.A2(n_4336),
.B(n_4335),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7679),
.Y(n_8193)
);

AOI22xp5_ASAP7_75t_L g8194 ( 
.A1(n_7730),
.A2(n_4340),
.B1(n_4343),
.B2(n_4339),
.Y(n_8194)
);

NAND2xp5_ASAP7_75t_SL g8195 ( 
.A(n_7545),
.B(n_4347),
.Y(n_8195)
);

INVx2_ASAP7_75t_L g8196 ( 
.A(n_7802),
.Y(n_8196)
);

INVx2_ASAP7_75t_L g8197 ( 
.A(n_7804),
.Y(n_8197)
);

INVxp67_ASAP7_75t_SL g8198 ( 
.A(n_7557),
.Y(n_8198)
);

NAND2xp5_ASAP7_75t_L g8199 ( 
.A(n_7791),
.B(n_4436),
.Y(n_8199)
);

NAND2xp5_ASAP7_75t_L g8200 ( 
.A(n_7792),
.B(n_4437),
.Y(n_8200)
);

INVx2_ASAP7_75t_L g8201 ( 
.A(n_7680),
.Y(n_8201)
);

NAND2xp5_ASAP7_75t_SL g8202 ( 
.A(n_7566),
.B(n_7977),
.Y(n_8202)
);

AND2x2_ASAP7_75t_L g8203 ( 
.A(n_7819),
.B(n_4349),
.Y(n_8203)
);

AND2x2_ASAP7_75t_L g8204 ( 
.A(n_7981),
.B(n_4357),
.Y(n_8204)
);

INVx2_ASAP7_75t_SL g8205 ( 
.A(n_7841),
.Y(n_8205)
);

BUFx3_ASAP7_75t_L g8206 ( 
.A(n_7570),
.Y(n_8206)
);

NAND2xp5_ASAP7_75t_L g8207 ( 
.A(n_7794),
.B(n_4438),
.Y(n_8207)
);

NOR2xp33_ASAP7_75t_L g8208 ( 
.A(n_7662),
.B(n_4361),
.Y(n_8208)
);

AND2x2_ASAP7_75t_L g8209 ( 
.A(n_7618),
.B(n_7626),
.Y(n_8209)
);

NAND2xp5_ASAP7_75t_L g8210 ( 
.A(n_7796),
.B(n_4444),
.Y(n_8210)
);

INVx2_ASAP7_75t_SL g8211 ( 
.A(n_7631),
.Y(n_8211)
);

NAND2xp5_ASAP7_75t_L g8212 ( 
.A(n_7799),
.B(n_7581),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_7583),
.B(n_4450),
.Y(n_8213)
);

NAND2xp5_ASAP7_75t_L g8214 ( 
.A(n_7585),
.B(n_4460),
.Y(n_8214)
);

AND2x2_ASAP7_75t_L g8215 ( 
.A(n_7641),
.B(n_4362),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7683),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_SL g8217 ( 
.A(n_7883),
.B(n_4363),
.Y(n_8217)
);

NAND2xp5_ASAP7_75t_L g8218 ( 
.A(n_7588),
.B(n_4481),
.Y(n_8218)
);

BUFx5_ASAP7_75t_L g8219 ( 
.A(n_7779),
.Y(n_8219)
);

NOR2xp33_ASAP7_75t_L g8220 ( 
.A(n_7633),
.B(n_4365),
.Y(n_8220)
);

OR2x6_ASAP7_75t_L g8221 ( 
.A(n_7708),
.B(n_4489),
.Y(n_8221)
);

NAND2xp33_ASAP7_75t_L g8222 ( 
.A(n_7779),
.B(n_4368),
.Y(n_8222)
);

AND2x2_ASAP7_75t_L g8223 ( 
.A(n_7646),
.B(n_4369),
.Y(n_8223)
);

INVx2_ASAP7_75t_SL g8224 ( 
.A(n_7648),
.Y(n_8224)
);

INVx2_ASAP7_75t_L g8225 ( 
.A(n_7688),
.Y(n_8225)
);

INVx2_ASAP7_75t_SL g8226 ( 
.A(n_7648),
.Y(n_8226)
);

AND2x6_ASAP7_75t_SL g8227 ( 
.A(n_8015),
.B(n_4494),
.Y(n_8227)
);

NOR2xp33_ASAP7_75t_L g8228 ( 
.A(n_7980),
.B(n_4370),
.Y(n_8228)
);

INVx2_ASAP7_75t_SL g8229 ( 
.A(n_7834),
.Y(n_8229)
);

NOR2xp33_ASAP7_75t_L g8230 ( 
.A(n_7830),
.B(n_4372),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_7591),
.B(n_4497),
.Y(n_8231)
);

NOR2xp67_ASAP7_75t_L g8232 ( 
.A(n_7920),
.B(n_8),
.Y(n_8232)
);

NAND3xp33_ASAP7_75t_L g8233 ( 
.A(n_7966),
.B(n_7944),
.C(n_7956),
.Y(n_8233)
);

INVxp33_ASAP7_75t_L g8234 ( 
.A(n_7532),
.Y(n_8234)
);

INVx3_ASAP7_75t_L g8235 ( 
.A(n_7539),
.Y(n_8235)
);

INVx2_ASAP7_75t_SL g8236 ( 
.A(n_7834),
.Y(n_8236)
);

NAND2xp5_ASAP7_75t_L g8237 ( 
.A(n_7594),
.B(n_4499),
.Y(n_8237)
);

INVx8_ASAP7_75t_L g8238 ( 
.A(n_7722),
.Y(n_8238)
);

AOI22xp5_ASAP7_75t_L g8239 ( 
.A1(n_7624),
.A2(n_4379),
.B1(n_4381),
.B2(n_4376),
.Y(n_8239)
);

INVx2_ASAP7_75t_L g8240 ( 
.A(n_7690),
.Y(n_8240)
);

AND2x4_ASAP7_75t_L g8241 ( 
.A(n_7562),
.B(n_4506),
.Y(n_8241)
);

INVx1_ASAP7_75t_L g8242 ( 
.A(n_7691),
.Y(n_8242)
);

AOI22xp33_ASAP7_75t_L g8243 ( 
.A1(n_7948),
.A2(n_4513),
.B1(n_4516),
.B2(n_4510),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7693),
.Y(n_8244)
);

NOR3xp33_ASAP7_75t_L g8245 ( 
.A(n_7916),
.B(n_4527),
.C(n_4521),
.Y(n_8245)
);

NAND2xp5_ASAP7_75t_SL g8246 ( 
.A(n_8011),
.B(n_4382),
.Y(n_8246)
);

NOR2xp33_ASAP7_75t_L g8247 ( 
.A(n_7996),
.B(n_4388),
.Y(n_8247)
);

BUFx5_ASAP7_75t_L g8248 ( 
.A(n_7590),
.Y(n_8248)
);

AND2x2_ASAP7_75t_L g8249 ( 
.A(n_7816),
.B(n_4389),
.Y(n_8249)
);

NOR2xp33_ASAP7_75t_L g8250 ( 
.A(n_7999),
.B(n_4391),
.Y(n_8250)
);

INVx2_ASAP7_75t_L g8251 ( 
.A(n_7696),
.Y(n_8251)
);

NAND2xp5_ASAP7_75t_L g8252 ( 
.A(n_7595),
.B(n_4530),
.Y(n_8252)
);

O2A1O1Ixp5_ASAP7_75t_L g8253 ( 
.A1(n_7882),
.A2(n_4534),
.B(n_4546),
.C(n_4532),
.Y(n_8253)
);

INVx1_ASAP7_75t_L g8254 ( 
.A(n_7699),
.Y(n_8254)
);

NOR2xp67_ASAP7_75t_L g8255 ( 
.A(n_7929),
.B(n_8),
.Y(n_8255)
);

NAND2xp5_ASAP7_75t_SL g8256 ( 
.A(n_7599),
.B(n_4392),
.Y(n_8256)
);

INVx2_ASAP7_75t_L g8257 ( 
.A(n_7700),
.Y(n_8257)
);

NOR2xp33_ASAP7_75t_L g8258 ( 
.A(n_8003),
.B(n_4397),
.Y(n_8258)
);

INVx1_ASAP7_75t_L g8259 ( 
.A(n_7701),
.Y(n_8259)
);

NOR3xp33_ASAP7_75t_L g8260 ( 
.A(n_7987),
.B(n_8007),
.C(n_7886),
.Y(n_8260)
);

NAND2xp5_ASAP7_75t_SL g8261 ( 
.A(n_7533),
.B(n_4398),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_7703),
.Y(n_8262)
);

NAND2xp5_ASAP7_75t_SL g8263 ( 
.A(n_7540),
.B(n_4403),
.Y(n_8263)
);

NAND2xp5_ASAP7_75t_SL g8264 ( 
.A(n_7541),
.B(n_4408),
.Y(n_8264)
);

NAND2xp5_ASAP7_75t_L g8265 ( 
.A(n_7597),
.B(n_4552),
.Y(n_8265)
);

INVx2_ASAP7_75t_SL g8266 ( 
.A(n_7852),
.Y(n_8266)
);

NAND2xp5_ASAP7_75t_L g8267 ( 
.A(n_7600),
.B(n_7607),
.Y(n_8267)
);

AND2x2_ASAP7_75t_L g8268 ( 
.A(n_7783),
.B(n_4409),
.Y(n_8268)
);

INVx1_ASAP7_75t_L g8269 ( 
.A(n_7705),
.Y(n_8269)
);

INVx2_ASAP7_75t_L g8270 ( 
.A(n_7706),
.Y(n_8270)
);

NAND2xp33_ASAP7_75t_L g8271 ( 
.A(n_7590),
.B(n_4410),
.Y(n_8271)
);

A2O1A1Ixp33_ASAP7_75t_L g8272 ( 
.A1(n_7923),
.A2(n_4565),
.B(n_4570),
.C(n_4561),
.Y(n_8272)
);

INVx2_ASAP7_75t_SL g8273 ( 
.A(n_7852),
.Y(n_8273)
);

AOI22xp33_ASAP7_75t_L g8274 ( 
.A1(n_7975),
.A2(n_4573),
.B1(n_4579),
.B2(n_4571),
.Y(n_8274)
);

NAND2xp5_ASAP7_75t_L g8275 ( 
.A(n_7610),
.B(n_4581),
.Y(n_8275)
);

NOR2xp33_ASAP7_75t_L g8276 ( 
.A(n_8008),
.B(n_4411),
.Y(n_8276)
);

OAI22xp5_ASAP7_75t_SL g8277 ( 
.A1(n_7513),
.A2(n_4419),
.B1(n_4420),
.B2(n_4414),
.Y(n_8277)
);

OAI22xp33_ASAP7_75t_L g8278 ( 
.A1(n_7522),
.A2(n_4426),
.B1(n_4427),
.B2(n_4424),
.Y(n_8278)
);

NAND2xp5_ASAP7_75t_L g8279 ( 
.A(n_7615),
.B(n_4583),
.Y(n_8279)
);

NAND2xp5_ASAP7_75t_L g8280 ( 
.A(n_7621),
.B(n_7622),
.Y(n_8280)
);

INVx5_ASAP7_75t_L g8281 ( 
.A(n_7858),
.Y(n_8281)
);

INVx1_ASAP7_75t_L g8282 ( 
.A(n_7644),
.Y(n_8282)
);

NAND2xp5_ASAP7_75t_L g8283 ( 
.A(n_7634),
.B(n_4594),
.Y(n_8283)
);

NOR2xp33_ASAP7_75t_L g8284 ( 
.A(n_8010),
.B(n_4428),
.Y(n_8284)
);

INVx3_ASAP7_75t_L g8285 ( 
.A(n_7565),
.Y(n_8285)
);

NOR2xp33_ASAP7_75t_L g8286 ( 
.A(n_7988),
.B(n_4430),
.Y(n_8286)
);

INVx2_ASAP7_75t_SL g8287 ( 
.A(n_7858),
.Y(n_8287)
);

AND2x2_ASAP7_75t_L g8288 ( 
.A(n_7803),
.B(n_4431),
.Y(n_8288)
);

AND2x2_ASAP7_75t_L g8289 ( 
.A(n_7994),
.B(n_4435),
.Y(n_8289)
);

OAI22xp33_ASAP7_75t_L g8290 ( 
.A1(n_7547),
.A2(n_7870),
.B1(n_7608),
.B2(n_7930),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_7666),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7926),
.Y(n_8292)
);

AOI21xp5_ASAP7_75t_L g8293 ( 
.A1(n_7907),
.A2(n_4609),
.B(n_4599),
.Y(n_8293)
);

INVx2_ASAP7_75t_L g8294 ( 
.A(n_7669),
.Y(n_8294)
);

INVx1_ASAP7_75t_L g8295 ( 
.A(n_7673),
.Y(n_8295)
);

NAND2xp5_ASAP7_75t_SL g8296 ( 
.A(n_7551),
.B(n_4441),
.Y(n_8296)
);

NAND2xp5_ASAP7_75t_L g8297 ( 
.A(n_7637),
.B(n_4622),
.Y(n_8297)
);

NAND2xp5_ASAP7_75t_L g8298 ( 
.A(n_7639),
.B(n_4627),
.Y(n_8298)
);

NAND2xp5_ASAP7_75t_SL g8299 ( 
.A(n_7556),
.B(n_4443),
.Y(n_8299)
);

INVx2_ASAP7_75t_L g8300 ( 
.A(n_7675),
.Y(n_8300)
);

INVx1_ASAP7_75t_L g8301 ( 
.A(n_7682),
.Y(n_8301)
);

NOR2xp33_ASAP7_75t_L g8302 ( 
.A(n_7990),
.B(n_4445),
.Y(n_8302)
);

NAND2xp5_ASAP7_75t_L g8303 ( 
.A(n_7643),
.B(n_4629),
.Y(n_8303)
);

INVx2_ASAP7_75t_L g8304 ( 
.A(n_7687),
.Y(n_8304)
);

INVx2_ASAP7_75t_SL g8305 ( 
.A(n_7863),
.Y(n_8305)
);

XNOR2xp5_ASAP7_75t_L g8306 ( 
.A(n_7584),
.B(n_4452),
.Y(n_8306)
);

NAND2xp5_ASAP7_75t_L g8307 ( 
.A(n_7563),
.B(n_4634),
.Y(n_8307)
);

O2A1O1Ixp5_ASAP7_75t_L g8308 ( 
.A1(n_7787),
.A2(n_4641),
.B(n_4644),
.C(n_4636),
.Y(n_8308)
);

NAND2xp5_ASAP7_75t_L g8309 ( 
.A(n_7567),
.B(n_4646),
.Y(n_8309)
);

CKINVDCx5p33_ASAP7_75t_R g8310 ( 
.A(n_7698),
.Y(n_8310)
);

BUFx3_ASAP7_75t_L g8311 ( 
.A(n_7998),
.Y(n_8311)
);

INVx2_ASAP7_75t_L g8312 ( 
.A(n_7695),
.Y(n_8312)
);

NAND2xp5_ASAP7_75t_L g8313 ( 
.A(n_7580),
.B(n_4657),
.Y(n_8313)
);

OAI21xp5_ASAP7_75t_L g8314 ( 
.A1(n_7972),
.A2(n_4662),
.B(n_4658),
.Y(n_8314)
);

INVx2_ASAP7_75t_L g8315 ( 
.A(n_7702),
.Y(n_8315)
);

INVx3_ASAP7_75t_L g8316 ( 
.A(n_7863),
.Y(n_8316)
);

AND2x2_ASAP7_75t_L g8317 ( 
.A(n_7941),
.B(n_4454),
.Y(n_8317)
);

AOI22xp5_ASAP7_75t_L g8318 ( 
.A1(n_7983),
.A2(n_4456),
.B1(n_4459),
.B2(n_4455),
.Y(n_8318)
);

NOR2xp33_ASAP7_75t_L g8319 ( 
.A(n_7991),
.B(n_4461),
.Y(n_8319)
);

NOR2xp33_ASAP7_75t_L g8320 ( 
.A(n_7992),
.B(n_4466),
.Y(n_8320)
);

NOR2xp33_ASAP7_75t_SL g8321 ( 
.A(n_7707),
.B(n_4467),
.Y(n_8321)
);

INVx2_ASAP7_75t_SL g8322 ( 
.A(n_7949),
.Y(n_8322)
);

NAND2xp5_ASAP7_75t_SL g8323 ( 
.A(n_7603),
.B(n_4469),
.Y(n_8323)
);

HB1xp67_ASAP7_75t_L g8324 ( 
.A(n_8009),
.Y(n_8324)
);

NAND2xp5_ASAP7_75t_L g8325 ( 
.A(n_7605),
.B(n_4671),
.Y(n_8325)
);

NAND2xp5_ASAP7_75t_L g8326 ( 
.A(n_7630),
.B(n_4672),
.Y(n_8326)
);

AOI21xp5_ASAP7_75t_L g8327 ( 
.A1(n_7927),
.A2(n_4686),
.B(n_4676),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_L g8328 ( 
.A(n_7750),
.B(n_7807),
.Y(n_8328)
);

INVx3_ASAP7_75t_L g8329 ( 
.A(n_7949),
.Y(n_8329)
);

INVx3_ASAP7_75t_L g8330 ( 
.A(n_7974),
.Y(n_8330)
);

BUFx3_ASAP7_75t_L g8331 ( 
.A(n_7974),
.Y(n_8331)
);

NAND2xp5_ASAP7_75t_L g8332 ( 
.A(n_7839),
.B(n_4691),
.Y(n_8332)
);

OAI22xp5_ASAP7_75t_SL g8333 ( 
.A1(n_7689),
.A2(n_7928),
.B1(n_7914),
.B2(n_7769),
.Y(n_8333)
);

INVx2_ASAP7_75t_L g8334 ( 
.A(n_7712),
.Y(n_8334)
);

NOR2xp33_ASAP7_75t_L g8335 ( 
.A(n_7993),
.B(n_7801),
.Y(n_8335)
);

NOR2xp33_ASAP7_75t_L g8336 ( 
.A(n_7808),
.B(n_4470),
.Y(n_8336)
);

AOI22xp5_ASAP7_75t_L g8337 ( 
.A1(n_8004),
.A2(n_4475),
.B1(n_4477),
.B2(n_4473),
.Y(n_8337)
);

NAND2xp5_ASAP7_75t_SL g8338 ( 
.A(n_7828),
.B(n_4478),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_7884),
.Y(n_8339)
);

INVx2_ASAP7_75t_SL g8340 ( 
.A(n_7718),
.Y(n_8340)
);

INVx1_ASAP7_75t_L g8341 ( 
.A(n_7885),
.Y(n_8341)
);

NAND2xp5_ASAP7_75t_L g8342 ( 
.A(n_7840),
.B(n_4701),
.Y(n_8342)
);

NAND2xp5_ASAP7_75t_L g8343 ( 
.A(n_7846),
.B(n_4702),
.Y(n_8343)
);

NAND2xp5_ASAP7_75t_L g8344 ( 
.A(n_7714),
.B(n_4707),
.Y(n_8344)
);

AND2x6_ASAP7_75t_L g8345 ( 
.A(n_7969),
.B(n_4708),
.Y(n_8345)
);

NAND2xp5_ASAP7_75t_L g8346 ( 
.A(n_7715),
.B(n_4721),
.Y(n_8346)
);

INVx1_ASAP7_75t_L g8347 ( 
.A(n_7889),
.Y(n_8347)
);

INVx2_ASAP7_75t_L g8348 ( 
.A(n_7716),
.Y(n_8348)
);

NOR2xp33_ASAP7_75t_L g8349 ( 
.A(n_7978),
.B(n_4479),
.Y(n_8349)
);

NOR2xp33_ASAP7_75t_L g8350 ( 
.A(n_7756),
.B(n_4480),
.Y(n_8350)
);

NOR2xp67_ASAP7_75t_SL g8351 ( 
.A(n_7720),
.B(n_4482),
.Y(n_8351)
);

NOR2xp33_ASAP7_75t_L g8352 ( 
.A(n_7672),
.B(n_4487),
.Y(n_8352)
);

INVx1_ASAP7_75t_L g8353 ( 
.A(n_7892),
.Y(n_8353)
);

NAND2xp5_ASAP7_75t_L g8354 ( 
.A(n_7717),
.B(n_4735),
.Y(n_8354)
);

AND2x2_ASAP7_75t_L g8355 ( 
.A(n_7951),
.B(n_4490),
.Y(n_8355)
);

NAND2xp5_ASAP7_75t_L g8356 ( 
.A(n_7724),
.B(n_4740),
.Y(n_8356)
);

NAND2xp5_ASAP7_75t_L g8357 ( 
.A(n_7728),
.B(n_4746),
.Y(n_8357)
);

AOI21xp5_ASAP7_75t_L g8358 ( 
.A1(n_7934),
.A2(n_4752),
.B(n_4751),
.Y(n_8358)
);

NOR2xp33_ASAP7_75t_L g8359 ( 
.A(n_7917),
.B(n_4493),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7894),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_7729),
.Y(n_8361)
);

NAND2xp5_ASAP7_75t_L g8362 ( 
.A(n_7732),
.B(n_4766),
.Y(n_8362)
);

OR2x6_ASAP7_75t_L g8363 ( 
.A(n_7910),
.B(n_4780),
.Y(n_8363)
);

AND2x2_ASAP7_75t_L g8364 ( 
.A(n_7967),
.B(n_4495),
.Y(n_8364)
);

NAND2xp5_ASAP7_75t_L g8365 ( 
.A(n_7733),
.B(n_4781),
.Y(n_8365)
);

NAND2xp5_ASAP7_75t_L g8366 ( 
.A(n_7897),
.B(n_4787),
.Y(n_8366)
);

NAND2xp5_ASAP7_75t_L g8367 ( 
.A(n_7514),
.B(n_4801),
.Y(n_8367)
);

INVxp67_ASAP7_75t_L g8368 ( 
.A(n_7979),
.Y(n_8368)
);

OAI22xp5_ASAP7_75t_L g8369 ( 
.A1(n_7896),
.A2(n_4503),
.B1(n_4505),
.B2(n_4500),
.Y(n_8369)
);

NOR2xp33_ASAP7_75t_L g8370 ( 
.A(n_8017),
.B(n_7635),
.Y(n_8370)
);

NAND2xp5_ASAP7_75t_L g8371 ( 
.A(n_7514),
.B(n_4805),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_7735),
.Y(n_8372)
);

OR2x2_ASAP7_75t_L g8373 ( 
.A(n_7955),
.B(n_4508),
.Y(n_8373)
);

NAND2xp5_ASAP7_75t_L g8374 ( 
.A(n_7514),
.B(n_4817),
.Y(n_8374)
);

AND2x2_ASAP7_75t_L g8375 ( 
.A(n_7758),
.B(n_4511),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7738),
.Y(n_8376)
);

NAND2xp5_ASAP7_75t_SL g8377 ( 
.A(n_7989),
.B(n_4514),
.Y(n_8377)
);

NAND2xp5_ASAP7_75t_L g8378 ( 
.A(n_7811),
.B(n_4832),
.Y(n_8378)
);

AOI22xp5_ASAP7_75t_L g8379 ( 
.A1(n_7878),
.A2(n_4517),
.B1(n_4518),
.B2(n_4515),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7740),
.Y(n_8380)
);

NAND2xp5_ASAP7_75t_L g8381 ( 
.A(n_7814),
.B(n_4846),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_7742),
.Y(n_8382)
);

NOR2xp33_ASAP7_75t_L g8383 ( 
.A(n_7842),
.B(n_4520),
.Y(n_8383)
);

HB1xp67_ASAP7_75t_L g8384 ( 
.A(n_7915),
.Y(n_8384)
);

INVx3_ASAP7_75t_L g8385 ( 
.A(n_7773),
.Y(n_8385)
);

INVx2_ASAP7_75t_SL g8386 ( 
.A(n_8001),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7743),
.Y(n_8387)
);

NOR3xp33_ASAP7_75t_L g8388 ( 
.A(n_8000),
.B(n_4855),
.C(n_4848),
.Y(n_8388)
);

AND2x2_ASAP7_75t_L g8389 ( 
.A(n_7737),
.B(n_4524),
.Y(n_8389)
);

INVx2_ASAP7_75t_L g8390 ( 
.A(n_7726),
.Y(n_8390)
);

INVx2_ASAP7_75t_SL g8391 ( 
.A(n_7771),
.Y(n_8391)
);

CKINVDCx11_ASAP7_75t_R g8392 ( 
.A(n_7704),
.Y(n_8392)
);

NOR2xp33_ASAP7_75t_L g8393 ( 
.A(n_7958),
.B(n_4526),
.Y(n_8393)
);

NOR2xp33_ASAP7_75t_L g8394 ( 
.A(n_7959),
.B(n_4528),
.Y(n_8394)
);

NAND2xp5_ASAP7_75t_L g8395 ( 
.A(n_7744),
.B(n_4856),
.Y(n_8395)
);

NAND2xp5_ASAP7_75t_L g8396 ( 
.A(n_7745),
.B(n_4859),
.Y(n_8396)
);

NOR2xp33_ASAP7_75t_L g8397 ( 
.A(n_7962),
.B(n_7964),
.Y(n_8397)
);

INVx8_ASAP7_75t_L g8398 ( 
.A(n_7810),
.Y(n_8398)
);

INVx2_ASAP7_75t_L g8399 ( 
.A(n_7747),
.Y(n_8399)
);

INVx2_ASAP7_75t_L g8400 ( 
.A(n_7748),
.Y(n_8400)
);

INVx3_ASAP7_75t_L g8401 ( 
.A(n_7853),
.Y(n_8401)
);

AND2x4_ASAP7_75t_SL g8402 ( 
.A(n_7638),
.B(n_4860),
.Y(n_8402)
);

NAND2xp5_ASAP7_75t_SL g8403 ( 
.A(n_7957),
.B(n_4529),
.Y(n_8403)
);

AND2x6_ASAP7_75t_L g8404 ( 
.A(n_7971),
.B(n_4861),
.Y(n_8404)
);

INVx3_ASAP7_75t_L g8405 ( 
.A(n_7813),
.Y(n_8405)
);

AND2x4_ASAP7_75t_L g8406 ( 
.A(n_7535),
.B(n_4863),
.Y(n_8406)
);

NAND2xp5_ASAP7_75t_L g8407 ( 
.A(n_7751),
.B(n_7752),
.Y(n_8407)
);

OR2x6_ASAP7_75t_L g8408 ( 
.A(n_7862),
.B(n_871),
.Y(n_8408)
);

INVx2_ASAP7_75t_L g8409 ( 
.A(n_7754),
.Y(n_8409)
);

NOR2xp33_ASAP7_75t_L g8410 ( 
.A(n_7931),
.B(n_4531),
.Y(n_8410)
);

NAND2xp5_ASAP7_75t_L g8411 ( 
.A(n_7755),
.B(n_4533),
.Y(n_8411)
);

NOR2xp33_ASAP7_75t_L g8412 ( 
.A(n_7932),
.B(n_4536),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_7757),
.Y(n_8413)
);

AND2x6_ASAP7_75t_SL g8414 ( 
.A(n_7930),
.B(n_4537),
.Y(n_8414)
);

NAND2x1_ASAP7_75t_L g8415 ( 
.A(n_7590),
.B(n_871),
.Y(n_8415)
);

INVx2_ASAP7_75t_L g8416 ( 
.A(n_7761),
.Y(n_8416)
);

NAND2xp33_ASAP7_75t_L g8417 ( 
.A(n_7557),
.B(n_7654),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_7762),
.Y(n_8418)
);

NAND2xp5_ASAP7_75t_L g8419 ( 
.A(n_7765),
.B(n_4539),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_7766),
.Y(n_8420)
);

OR2x6_ASAP7_75t_L g8421 ( 
.A(n_7887),
.B(n_872),
.Y(n_8421)
);

NAND2xp5_ASAP7_75t_SL g8422 ( 
.A(n_7759),
.B(n_4540),
.Y(n_8422)
);

INVx2_ASAP7_75t_L g8423 ( 
.A(n_7767),
.Y(n_8423)
);

AND2x2_ASAP7_75t_L g8424 ( 
.A(n_7845),
.B(n_7961),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_7768),
.Y(n_8425)
);

NOR2xp33_ASAP7_75t_L g8426 ( 
.A(n_7935),
.B(n_4542),
.Y(n_8426)
);

NAND2xp5_ASAP7_75t_L g8427 ( 
.A(n_7770),
.B(n_4544),
.Y(n_8427)
);

INVxp67_ASAP7_75t_L g8428 ( 
.A(n_7775),
.Y(n_8428)
);

NAND2xp5_ASAP7_75t_L g8429 ( 
.A(n_7772),
.B(n_4545),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_7774),
.Y(n_8430)
);

AOI21xp5_ASAP7_75t_L g8431 ( 
.A1(n_7921),
.A2(n_4548),
.B(n_4547),
.Y(n_8431)
);

NAND2xp5_ASAP7_75t_L g8432 ( 
.A(n_7776),
.B(n_4550),
.Y(n_8432)
);

NAND2xp5_ASAP7_75t_SL g8433 ( 
.A(n_8012),
.B(n_4553),
.Y(n_8433)
);

INVx2_ASAP7_75t_L g8434 ( 
.A(n_7780),
.Y(n_8434)
);

BUFx3_ASAP7_75t_L g8435 ( 
.A(n_8014),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7781),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_L g8437 ( 
.A(n_7782),
.B(n_4554),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7784),
.Y(n_8438)
);

AND2x2_ASAP7_75t_L g8439 ( 
.A(n_7982),
.B(n_4555),
.Y(n_8439)
);

OR2x2_ASAP7_75t_L g8440 ( 
.A(n_8016),
.B(n_4557),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_7786),
.B(n_4560),
.Y(n_8441)
);

NAND2xp5_ASAP7_75t_L g8442 ( 
.A(n_7805),
.B(n_4568),
.Y(n_8442)
);

NAND2xp5_ASAP7_75t_L g8443 ( 
.A(n_7815),
.B(n_4572),
.Y(n_8443)
);

CKINVDCx5p33_ASAP7_75t_R g8444 ( 
.A(n_7663),
.Y(n_8444)
);

AOI22xp5_ASAP7_75t_L g8445 ( 
.A1(n_7963),
.A2(n_4575),
.B1(n_4577),
.B2(n_4574),
.Y(n_8445)
);

OAI221xp5_ASAP7_75t_L g8446 ( 
.A1(n_7843),
.A2(n_4585),
.B1(n_4586),
.B2(n_4580),
.C(n_4578),
.Y(n_8446)
);

NAND2xp5_ASAP7_75t_L g8447 ( 
.A(n_7817),
.B(n_4592),
.Y(n_8447)
);

BUFx2_ASAP7_75t_L g8448 ( 
.A(n_7596),
.Y(n_8448)
);

INVxp67_ASAP7_75t_L g8449 ( 
.A(n_7997),
.Y(n_8449)
);

INVx1_ASAP7_75t_L g8450 ( 
.A(n_7881),
.Y(n_8450)
);

INVx2_ASAP7_75t_L g8451 ( 
.A(n_7844),
.Y(n_8451)
);

NAND2xp5_ASAP7_75t_L g8452 ( 
.A(n_7820),
.B(n_4600),
.Y(n_8452)
);

NAND2xp5_ASAP7_75t_SL g8453 ( 
.A(n_7822),
.B(n_4602),
.Y(n_8453)
);

NAND2xp5_ASAP7_75t_SL g8454 ( 
.A(n_7904),
.B(n_7945),
.Y(n_8454)
);

NAND2xp5_ASAP7_75t_SL g8455 ( 
.A(n_7640),
.B(n_7574),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_7825),
.B(n_4606),
.Y(n_8456)
);

AOI22xp33_ASAP7_75t_L g8457 ( 
.A1(n_7692),
.A2(n_4610),
.B1(n_4611),
.B2(n_4607),
.Y(n_8457)
);

NAND2xp33_ASAP7_75t_L g8458 ( 
.A(n_7557),
.B(n_4612),
.Y(n_8458)
);

NOR2xp33_ASAP7_75t_L g8459 ( 
.A(n_7936),
.B(n_4617),
.Y(n_8459)
);

INVx2_ASAP7_75t_SL g8460 ( 
.A(n_7968),
.Y(n_8460)
);

INVx3_ASAP7_75t_L g8461 ( 
.A(n_7984),
.Y(n_8461)
);

NAND2xp5_ASAP7_75t_SL g8462 ( 
.A(n_7869),
.B(n_4618),
.Y(n_8462)
);

OR2x2_ASAP7_75t_L g8463 ( 
.A(n_7826),
.B(n_4623),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_7827),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_L g8465 ( 
.A(n_7829),
.B(n_4624),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_7831),
.Y(n_8466)
);

AOI22xp5_ASAP7_75t_L g8467 ( 
.A1(n_7888),
.A2(n_4630),
.B1(n_4631),
.B2(n_4626),
.Y(n_8467)
);

INVx1_ASAP7_75t_L g8468 ( 
.A(n_7832),
.Y(n_8468)
);

INVx2_ASAP7_75t_L g8469 ( 
.A(n_7874),
.Y(n_8469)
);

NAND2xp5_ASAP7_75t_L g8470 ( 
.A(n_7833),
.B(n_7857),
.Y(n_8470)
);

INVx3_ASAP7_75t_L g8471 ( 
.A(n_8013),
.Y(n_8471)
);

NAND2xp5_ASAP7_75t_L g8472 ( 
.A(n_7861),
.B(n_4632),
.Y(n_8472)
);

AND2x2_ASAP7_75t_L g8473 ( 
.A(n_7953),
.B(n_7870),
.Y(n_8473)
);

AOI22xp5_ASAP7_75t_L g8474 ( 
.A1(n_7627),
.A2(n_4643),
.B1(n_4648),
.B2(n_4635),
.Y(n_8474)
);

INVxp33_ASAP7_75t_L g8475 ( 
.A(n_7564),
.Y(n_8475)
);

INVxp33_ASAP7_75t_SL g8476 ( 
.A(n_7763),
.Y(n_8476)
);

NAND2xp5_ASAP7_75t_SL g8477 ( 
.A(n_7937),
.B(n_4650),
.Y(n_8477)
);

NOR2xp33_ASAP7_75t_L g8478 ( 
.A(n_7938),
.B(n_4652),
.Y(n_8478)
);

NOR2xp67_ASAP7_75t_L g8479 ( 
.A(n_7939),
.B(n_8),
.Y(n_8479)
);

INVx2_ASAP7_75t_L g8480 ( 
.A(n_7557),
.Y(n_8480)
);

AO22x1_ASAP7_75t_L g8481 ( 
.A1(n_7872),
.A2(n_4660),
.B1(n_4664),
.B2(n_4655),
.Y(n_8481)
);

BUFx5_ASAP7_75t_L g8482 ( 
.A(n_7864),
.Y(n_8482)
);

INVxp67_ASAP7_75t_L g8483 ( 
.A(n_7764),
.Y(n_8483)
);

NAND2xp5_ASAP7_75t_L g8484 ( 
.A(n_7865),
.B(n_4665),
.Y(n_8484)
);

NAND2xp5_ASAP7_75t_L g8485 ( 
.A(n_7866),
.B(n_4666),
.Y(n_8485)
);

O2A1O1Ixp5_ASAP7_75t_L g8486 ( 
.A1(n_7946),
.A2(n_874),
.B(n_875),
.C(n_872),
.Y(n_8486)
);

INVx2_ASAP7_75t_SL g8487 ( 
.A(n_8019),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_7867),
.Y(n_8488)
);

AOI21xp5_ASAP7_75t_L g8489 ( 
.A1(n_7965),
.A2(n_4669),
.B(n_4667),
.Y(n_8489)
);

NAND2xp5_ASAP7_75t_SL g8490 ( 
.A(n_7947),
.B(n_4670),
.Y(n_8490)
);

INVx1_ASAP7_75t_L g8491 ( 
.A(n_7871),
.Y(n_8491)
);

NAND2xp5_ASAP7_75t_L g8492 ( 
.A(n_7875),
.B(n_7879),
.Y(n_8492)
);

NAND3xp33_ASAP7_75t_L g8493 ( 
.A(n_7942),
.B(n_4677),
.C(n_4675),
.Y(n_8493)
);

AND2x2_ASAP7_75t_L g8494 ( 
.A(n_7880),
.B(n_4680),
.Y(n_8494)
);

AND2x2_ASAP7_75t_L g8495 ( 
.A(n_7950),
.B(n_4681),
.Y(n_8495)
);

INVx1_ASAP7_75t_L g8496 ( 
.A(n_7848),
.Y(n_8496)
);

AOI22xp5_ASAP7_75t_L g8497 ( 
.A1(n_7985),
.A2(n_4687),
.B1(n_4688),
.B2(n_4685),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_7849),
.Y(n_8498)
);

OAI22xp33_ASAP7_75t_L g8499 ( 
.A1(n_7942),
.A2(n_4694),
.B1(n_4699),
.B2(n_4689),
.Y(n_8499)
);

NAND2xp5_ASAP7_75t_L g8500 ( 
.A(n_7851),
.B(n_4703),
.Y(n_8500)
);

INVx3_ASAP7_75t_L g8501 ( 
.A(n_8020),
.Y(n_8501)
);

AND2x2_ASAP7_75t_L g8502 ( 
.A(n_7649),
.B(n_7681),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_SL g8503 ( 
.A(n_7855),
.B(n_7899),
.Y(n_8503)
);

NAND2xp5_ASAP7_75t_L g8504 ( 
.A(n_7900),
.B(n_4704),
.Y(n_8504)
);

HB1xp67_ASAP7_75t_L g8505 ( 
.A(n_7704),
.Y(n_8505)
);

OAI22xp5_ASAP7_75t_L g8506 ( 
.A1(n_8005),
.A2(n_4706),
.B1(n_4709),
.B2(n_4705),
.Y(n_8506)
);

NOR2xp33_ASAP7_75t_L g8507 ( 
.A(n_7636),
.B(n_4717),
.Y(n_8507)
);

NAND2xp5_ASAP7_75t_L g8508 ( 
.A(n_7654),
.B(n_4719),
.Y(n_8508)
);

NOR2xp33_ASAP7_75t_L g8509 ( 
.A(n_7654),
.B(n_4722),
.Y(n_8509)
);

NAND2xp5_ASAP7_75t_L g8510 ( 
.A(n_7654),
.B(n_4723),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_7809),
.Y(n_8511)
);

NAND2xp5_ASAP7_75t_L g8512 ( 
.A(n_7685),
.B(n_4724),
.Y(n_8512)
);

INVx2_ASAP7_75t_L g8513 ( 
.A(n_7512),
.Y(n_8513)
);

NAND2xp5_ASAP7_75t_L g8514 ( 
.A(n_7685),
.B(n_4726),
.Y(n_8514)
);

INVx2_ASAP7_75t_L g8515 ( 
.A(n_7512),
.Y(n_8515)
);

OR2x2_ASAP7_75t_L g8516 ( 
.A(n_7559),
.B(n_4728),
.Y(n_8516)
);

INVxp67_ASAP7_75t_L g8517 ( 
.A(n_7559),
.Y(n_8517)
);

INVx2_ASAP7_75t_L g8518 ( 
.A(n_7512),
.Y(n_8518)
);

NAND2xp5_ASAP7_75t_SL g8519 ( 
.A(n_7685),
.B(n_4729),
.Y(n_8519)
);

NAND2xp5_ASAP7_75t_L g8520 ( 
.A(n_7685),
.B(n_4731),
.Y(n_8520)
);

AND2x6_ASAP7_75t_SL g8521 ( 
.A(n_7629),
.B(n_4741),
.Y(n_8521)
);

AOI22xp5_ASAP7_75t_L g8522 ( 
.A1(n_7685),
.A2(n_4743),
.B1(n_4744),
.B2(n_4742),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_7512),
.Y(n_8523)
);

NAND2xp5_ASAP7_75t_L g8524 ( 
.A(n_7685),
.B(n_4745),
.Y(n_8524)
);

NAND2xp5_ASAP7_75t_SL g8525 ( 
.A(n_7685),
.B(n_4747),
.Y(n_8525)
);

NAND2xp33_ASAP7_75t_L g8526 ( 
.A(n_7779),
.B(n_4748),
.Y(n_8526)
);

AOI22xp33_ASAP7_75t_L g8527 ( 
.A1(n_7657),
.A2(n_4754),
.B1(n_4755),
.B2(n_4753),
.Y(n_8527)
);

OAI22x1_ASAP7_75t_L g8528 ( 
.A1(n_7657),
.A2(n_4757),
.B1(n_4758),
.B2(n_4756),
.Y(n_8528)
);

NAND2xp5_ASAP7_75t_SL g8529 ( 
.A(n_7685),
.B(n_4759),
.Y(n_8529)
);

INVx1_ASAP7_75t_L g8530 ( 
.A(n_7512),
.Y(n_8530)
);

INVx2_ASAP7_75t_SL g8531 ( 
.A(n_8051),
.Y(n_8531)
);

AND2x2_ASAP7_75t_L g8532 ( 
.A(n_8209),
.B(n_4762),
.Y(n_8532)
);

AOI22xp5_ASAP7_75t_SL g8533 ( 
.A1(n_8036),
.A2(n_4764),
.B1(n_4769),
.B2(n_4763),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_L g8534 ( 
.A(n_8035),
.B(n_4770),
.Y(n_8534)
);

AND2x4_ASAP7_75t_L g8535 ( 
.A(n_8206),
.B(n_4777),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_SL g8536 ( 
.A(n_8150),
.B(n_4778),
.Y(n_8536)
);

OR2x2_ASAP7_75t_L g8537 ( 
.A(n_8517),
.B(n_4788),
.Y(n_8537)
);

NOR2xp33_ASAP7_75t_L g8538 ( 
.A(n_8031),
.B(n_4790),
.Y(n_8538)
);

NAND2xp5_ASAP7_75t_L g8539 ( 
.A(n_8168),
.B(n_8109),
.Y(n_8539)
);

NAND2xp5_ASAP7_75t_SL g8540 ( 
.A(n_8233),
.B(n_4800),
.Y(n_8540)
);

OAI21xp33_ASAP7_75t_L g8541 ( 
.A1(n_8123),
.A2(n_4804),
.B(n_4802),
.Y(n_8541)
);

NAND2xp5_ASAP7_75t_L g8542 ( 
.A(n_8038),
.B(n_4809),
.Y(n_8542)
);

NOR2xp33_ASAP7_75t_L g8543 ( 
.A(n_8069),
.B(n_4811),
.Y(n_8543)
);

INVx4_ASAP7_75t_L g8544 ( 
.A(n_8281),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_8177),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_SL g8546 ( 
.A(n_8083),
.B(n_4812),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_8029),
.B(n_4814),
.Y(n_8547)
);

INVx2_ASAP7_75t_L g8548 ( 
.A(n_8023),
.Y(n_8548)
);

INVx2_ASAP7_75t_L g8549 ( 
.A(n_8026),
.Y(n_8549)
);

INVx3_ASAP7_75t_L g8550 ( 
.A(n_8311),
.Y(n_8550)
);

INVxp67_ASAP7_75t_SL g8551 ( 
.A(n_8053),
.Y(n_8551)
);

NAND2xp5_ASAP7_75t_SL g8552 ( 
.A(n_8085),
.B(n_4815),
.Y(n_8552)
);

AOI21xp5_ASAP7_75t_L g8553 ( 
.A1(n_8417),
.A2(n_8187),
.B(n_8458),
.Y(n_8553)
);

INVx2_ASAP7_75t_L g8554 ( 
.A(n_8030),
.Y(n_8554)
);

AOI22xp33_ASAP7_75t_L g8555 ( 
.A1(n_8260),
.A2(n_4828),
.B1(n_4830),
.B2(n_4820),
.Y(n_8555)
);

INVx1_ASAP7_75t_L g8556 ( 
.A(n_8328),
.Y(n_8556)
);

BUFx3_ASAP7_75t_L g8557 ( 
.A(n_8051),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_8040),
.Y(n_8558)
);

INVx2_ASAP7_75t_L g8559 ( 
.A(n_8047),
.Y(n_8559)
);

CKINVDCx5p33_ASAP7_75t_R g8560 ( 
.A(n_8392),
.Y(n_8560)
);

NAND2xp5_ASAP7_75t_L g8561 ( 
.A(n_8169),
.B(n_4835),
.Y(n_8561)
);

NAND2xp5_ASAP7_75t_SL g8562 ( 
.A(n_8082),
.B(n_4837),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_8049),
.Y(n_8563)
);

NAND2xp5_ASAP7_75t_SL g8564 ( 
.A(n_8164),
.B(n_4838),
.Y(n_8564)
);

INVx1_ASAP7_75t_SL g8565 ( 
.A(n_8074),
.Y(n_8565)
);

NOR2xp33_ASAP7_75t_R g8566 ( 
.A(n_8057),
.B(n_4841),
.Y(n_8566)
);

INVx3_ASAP7_75t_L g8567 ( 
.A(n_8181),
.Y(n_8567)
);

INVx1_ASAP7_75t_L g8568 ( 
.A(n_8050),
.Y(n_8568)
);

AND2x4_ASAP7_75t_L g8569 ( 
.A(n_8106),
.B(n_4842),
.Y(n_8569)
);

AND2x4_ASAP7_75t_L g8570 ( 
.A(n_8034),
.B(n_4844),
.Y(n_8570)
);

INVx2_ASAP7_75t_SL g8571 ( 
.A(n_8281),
.Y(n_8571)
);

AOI22xp33_ASAP7_75t_SL g8572 ( 
.A1(n_8333),
.A2(n_4847),
.B1(n_4852),
.B2(n_4845),
.Y(n_8572)
);

AND2x4_ASAP7_75t_L g8573 ( 
.A(n_8285),
.B(n_4853),
.Y(n_8573)
);

OAI22xp5_ASAP7_75t_L g8574 ( 
.A1(n_8044),
.A2(n_4864),
.B1(n_4866),
.B2(n_4858),
.Y(n_8574)
);

BUFx6f_ASAP7_75t_L g8575 ( 
.A(n_8129),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_L g8576 ( 
.A(n_8037),
.B(n_4867),
.Y(n_8576)
);

CKINVDCx5p33_ASAP7_75t_R g8577 ( 
.A(n_8135),
.Y(n_8577)
);

BUFx2_ASAP7_75t_L g8578 ( 
.A(n_8055),
.Y(n_8578)
);

NOR2xp33_ASAP7_75t_L g8579 ( 
.A(n_8350),
.B(n_4868),
.Y(n_8579)
);

NOR2xp33_ASAP7_75t_L g8580 ( 
.A(n_8108),
.B(n_4869),
.Y(n_8580)
);

OR2x2_ASAP7_75t_L g8581 ( 
.A(n_8022),
.B(n_4870),
.Y(n_8581)
);

OAI21xp5_ASAP7_75t_L g8582 ( 
.A1(n_8102),
.A2(n_4872),
.B(n_9),
.Y(n_8582)
);

NAND2xp5_ASAP7_75t_L g8583 ( 
.A(n_8073),
.B(n_9),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_8052),
.Y(n_8584)
);

OAI21xp5_ASAP7_75t_L g8585 ( 
.A1(n_8111),
.A2(n_9),
.B(n_10),
.Y(n_8585)
);

NAND2xp5_ASAP7_75t_L g8586 ( 
.A(n_8042),
.B(n_10),
.Y(n_8586)
);

OAI21xp5_ASAP7_75t_L g8587 ( 
.A1(n_8112),
.A2(n_10),
.B(n_11),
.Y(n_8587)
);

INVx2_ASAP7_75t_L g8588 ( 
.A(n_8065),
.Y(n_8588)
);

INVx1_ASAP7_75t_L g8589 ( 
.A(n_8068),
.Y(n_8589)
);

NOR2xp33_ASAP7_75t_L g8590 ( 
.A(n_8220),
.B(n_874),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_8077),
.Y(n_8591)
);

OAI21xp5_ASAP7_75t_L g8592 ( 
.A1(n_8128),
.A2(n_11),
.B(n_12),
.Y(n_8592)
);

AOI22xp5_ASAP7_75t_L g8593 ( 
.A1(n_8032),
.A2(n_8096),
.B1(n_8202),
.B2(n_8064),
.Y(n_8593)
);

AOI22xp33_ASAP7_75t_L g8594 ( 
.A1(n_8161),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_8594)
);

NAND2xp5_ASAP7_75t_L g8595 ( 
.A(n_8072),
.B(n_12),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_8093),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_8114),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_8116),
.Y(n_8598)
);

NAND2xp5_ASAP7_75t_L g8599 ( 
.A(n_8162),
.B(n_13),
.Y(n_8599)
);

CKINVDCx5p33_ASAP7_75t_R g8600 ( 
.A(n_8444),
.Y(n_8600)
);

NAND2xp5_ASAP7_75t_L g8601 ( 
.A(n_8166),
.B(n_13),
.Y(n_8601)
);

NAND2xp5_ASAP7_75t_L g8602 ( 
.A(n_8076),
.B(n_14),
.Y(n_8602)
);

NAND2xp5_ASAP7_75t_SL g8603 ( 
.A(n_8290),
.B(n_875),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8119),
.Y(n_8604)
);

AOI21xp5_ASAP7_75t_L g8605 ( 
.A1(n_8198),
.A2(n_877),
.B(n_876),
.Y(n_8605)
);

NAND2xp5_ASAP7_75t_L g8606 ( 
.A(n_8125),
.B(n_14),
.Y(n_8606)
);

AOI22xp33_ASAP7_75t_L g8607 ( 
.A1(n_8388),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_8607)
);

AOI22xp5_ASAP7_75t_L g8608 ( 
.A1(n_8230),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_8608)
);

INVx2_ASAP7_75t_SL g8609 ( 
.A(n_8281),
.Y(n_8609)
);

INVx1_ASAP7_75t_L g8610 ( 
.A(n_8120),
.Y(n_8610)
);

NOR2xp33_ASAP7_75t_R g8611 ( 
.A(n_8155),
.B(n_878),
.Y(n_8611)
);

NAND2xp5_ASAP7_75t_SL g8612 ( 
.A(n_8066),
.B(n_8183),
.Y(n_8612)
);

BUFx12f_ASAP7_75t_SL g8613 ( 
.A(n_8056),
.Y(n_8613)
);

INVx2_ASAP7_75t_L g8614 ( 
.A(n_8131),
.Y(n_8614)
);

NOR2xp33_ASAP7_75t_R g8615 ( 
.A(n_8092),
.B(n_878),
.Y(n_8615)
);

BUFx3_ASAP7_75t_L g8616 ( 
.A(n_8331),
.Y(n_8616)
);

NAND2xp5_ASAP7_75t_L g8617 ( 
.A(n_8126),
.B(n_17),
.Y(n_8617)
);

NAND2xp5_ASAP7_75t_L g8618 ( 
.A(n_8080),
.B(n_17),
.Y(n_8618)
);

NOR2xp33_ASAP7_75t_L g8619 ( 
.A(n_8154),
.B(n_879),
.Y(n_8619)
);

NAND2xp5_ASAP7_75t_L g8620 ( 
.A(n_8058),
.B(n_18),
.Y(n_8620)
);

NOR2x1p5_ASAP7_75t_L g8621 ( 
.A(n_8235),
.B(n_8401),
.Y(n_8621)
);

AND2x4_ASAP7_75t_L g8622 ( 
.A(n_8205),
.B(n_881),
.Y(n_8622)
);

INVx1_ASAP7_75t_L g8623 ( 
.A(n_8149),
.Y(n_8623)
);

NOR3xp33_ASAP7_75t_SL g8624 ( 
.A(n_8446),
.B(n_18),
.C(n_19),
.Y(n_8624)
);

NAND2xp5_ASAP7_75t_L g8625 ( 
.A(n_8059),
.B(n_8424),
.Y(n_8625)
);

INVx2_ASAP7_75t_L g8626 ( 
.A(n_8153),
.Y(n_8626)
);

AOI22xp5_ASAP7_75t_L g8627 ( 
.A1(n_8208),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_8627)
);

NOR2x1_ASAP7_75t_R g8628 ( 
.A(n_8310),
.B(n_881),
.Y(n_8628)
);

NAND2xp5_ASAP7_75t_L g8629 ( 
.A(n_8100),
.B(n_8512),
.Y(n_8629)
);

AO21x1_ASAP7_75t_L g8630 ( 
.A1(n_8314),
.A2(n_8178),
.B(n_8095),
.Y(n_8630)
);

INVx1_ASAP7_75t_L g8631 ( 
.A(n_8184),
.Y(n_8631)
);

INVx1_ASAP7_75t_L g8632 ( 
.A(n_8196),
.Y(n_8632)
);

BUFx3_ASAP7_75t_L g8633 ( 
.A(n_8129),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_8197),
.Y(n_8634)
);

NAND2x1p5_ASAP7_75t_L g8635 ( 
.A(n_8139),
.B(n_883),
.Y(n_8635)
);

A2O1A1Ixp33_ASAP7_75t_L g8636 ( 
.A1(n_8048),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_8636)
);

INVx2_ASAP7_75t_L g8637 ( 
.A(n_8201),
.Y(n_8637)
);

NAND2xp5_ASAP7_75t_L g8638 ( 
.A(n_8514),
.B(n_8520),
.Y(n_8638)
);

NAND2xp5_ASAP7_75t_L g8639 ( 
.A(n_8524),
.B(n_8075),
.Y(n_8639)
);

INVx1_ASAP7_75t_L g8640 ( 
.A(n_8225),
.Y(n_8640)
);

INVx2_ASAP7_75t_L g8641 ( 
.A(n_8240),
.Y(n_8641)
);

NAND2xp5_ASAP7_75t_L g8642 ( 
.A(n_8335),
.B(n_21),
.Y(n_8642)
);

NOR2x1_ASAP7_75t_R g8643 ( 
.A(n_8028),
.B(n_883),
.Y(n_8643)
);

NAND2xp5_ASAP7_75t_L g8644 ( 
.A(n_8146),
.B(n_21),
.Y(n_8644)
);

INVx2_ASAP7_75t_L g8645 ( 
.A(n_8251),
.Y(n_8645)
);

OR2x6_ASAP7_75t_L g8646 ( 
.A(n_8238),
.B(n_884),
.Y(n_8646)
);

BUFx6f_ASAP7_75t_L g8647 ( 
.A(n_8185),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8257),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_8270),
.Y(n_8649)
);

INVx2_ASAP7_75t_L g8650 ( 
.A(n_8513),
.Y(n_8650)
);

OR2x6_ASAP7_75t_SL g8651 ( 
.A(n_8493),
.B(n_22),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_L g8652 ( 
.A(n_8087),
.B(n_22),
.Y(n_8652)
);

INVx1_ASAP7_75t_L g8653 ( 
.A(n_8515),
.Y(n_8653)
);

AOI21xp5_ASAP7_75t_L g8654 ( 
.A1(n_8509),
.A2(n_885),
.B(n_884),
.Y(n_8654)
);

NOR2xp33_ASAP7_75t_L g8655 ( 
.A(n_8172),
.B(n_885),
.Y(n_8655)
);

BUFx3_ASAP7_75t_L g8656 ( 
.A(n_8185),
.Y(n_8656)
);

BUFx12f_ASAP7_75t_L g8657 ( 
.A(n_8041),
.Y(n_8657)
);

INVx2_ASAP7_75t_L g8658 ( 
.A(n_8518),
.Y(n_8658)
);

NAND2xp5_ASAP7_75t_SL g8659 ( 
.A(n_8027),
.B(n_886),
.Y(n_8659)
);

AOI21xp5_ASAP7_75t_L g8660 ( 
.A1(n_8179),
.A2(n_887),
.B(n_886),
.Y(n_8660)
);

NAND2xp5_ASAP7_75t_L g8661 ( 
.A(n_8151),
.B(n_22),
.Y(n_8661)
);

NAND2x1p5_ASAP7_75t_L g8662 ( 
.A(n_8097),
.B(n_887),
.Y(n_8662)
);

INVx5_ASAP7_75t_L g8663 ( 
.A(n_8238),
.Y(n_8663)
);

NOR2xp33_ASAP7_75t_L g8664 ( 
.A(n_8449),
.B(n_888),
.Y(n_8664)
);

HB1xp67_ASAP7_75t_L g8665 ( 
.A(n_8089),
.Y(n_8665)
);

INVxp67_ASAP7_75t_L g8666 ( 
.A(n_8384),
.Y(n_8666)
);

AND2x2_ASAP7_75t_L g8667 ( 
.A(n_8204),
.B(n_23),
.Y(n_8667)
);

AND2x2_ASAP7_75t_SL g8668 ( 
.A(n_8473),
.B(n_888),
.Y(n_8668)
);

NAND2xp5_ASAP7_75t_L g8669 ( 
.A(n_8115),
.B(n_8117),
.Y(n_8669)
);

NAND2xp5_ASAP7_75t_SL g8670 ( 
.A(n_8081),
.B(n_889),
.Y(n_8670)
);

AOI22xp5_ASAP7_75t_L g8671 ( 
.A1(n_8338),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_8671)
);

BUFx6f_ASAP7_75t_L g8672 ( 
.A(n_8170),
.Y(n_8672)
);

AOI22xp5_ASAP7_75t_L g8673 ( 
.A1(n_8483),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_8673)
);

AOI22x1_ASAP7_75t_L g8674 ( 
.A1(n_8528),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_8674)
);

NAND2xp5_ASAP7_75t_L g8675 ( 
.A(n_8156),
.B(n_26),
.Y(n_8675)
);

INVx2_ASAP7_75t_L g8676 ( 
.A(n_8334),
.Y(n_8676)
);

HB1xp67_ASAP7_75t_L g8677 ( 
.A(n_8324),
.Y(n_8677)
);

AOI22xp5_ASAP7_75t_L g8678 ( 
.A1(n_8099),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_8678)
);

INVx1_ASAP7_75t_L g8679 ( 
.A(n_8021),
.Y(n_8679)
);

INVx1_ASAP7_75t_L g8680 ( 
.A(n_8025),
.Y(n_8680)
);

NAND2xp33_ASAP7_75t_SL g8681 ( 
.A(n_8475),
.B(n_889),
.Y(n_8681)
);

INVx2_ASAP7_75t_SL g8682 ( 
.A(n_8316),
.Y(n_8682)
);

INVx3_ASAP7_75t_L g8683 ( 
.A(n_8180),
.Y(n_8683)
);

NOR2xp33_ASAP7_75t_L g8684 ( 
.A(n_8234),
.B(n_890),
.Y(n_8684)
);

AOI22xp5_ASAP7_75t_L g8685 ( 
.A1(n_8519),
.A2(n_8529),
.B1(n_8525),
.B2(n_8217),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_8046),
.Y(n_8686)
);

NOR2xp33_ASAP7_75t_L g8687 ( 
.A(n_8192),
.B(n_890),
.Y(n_8687)
);

INVx1_ASAP7_75t_L g8688 ( 
.A(n_8054),
.Y(n_8688)
);

AOI22xp33_ASAP7_75t_L g8689 ( 
.A1(n_8245),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8070),
.Y(n_8690)
);

NOR2xp33_ASAP7_75t_L g8691 ( 
.A(n_8370),
.B(n_891),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_8348),
.Y(n_8692)
);

INVx4_ASAP7_75t_L g8693 ( 
.A(n_8056),
.Y(n_8693)
);

BUFx6f_ASAP7_75t_L g8694 ( 
.A(n_8435),
.Y(n_8694)
);

NAND2xp5_ASAP7_75t_SL g8695 ( 
.A(n_8033),
.B(n_892),
.Y(n_8695)
);

HB1xp67_ASAP7_75t_L g8696 ( 
.A(n_8158),
.Y(n_8696)
);

CKINVDCx5p33_ASAP7_75t_R g8697 ( 
.A(n_8476),
.Y(n_8697)
);

OR2x6_ASAP7_75t_L g8698 ( 
.A(n_8398),
.B(n_892),
.Y(n_8698)
);

INVx1_ASAP7_75t_L g8699 ( 
.A(n_8078),
.Y(n_8699)
);

INVx4_ASAP7_75t_SL g8700 ( 
.A(n_8345),
.Y(n_8700)
);

INVx2_ASAP7_75t_L g8701 ( 
.A(n_8294),
.Y(n_8701)
);

OAI22xp5_ASAP7_75t_SL g8702 ( 
.A1(n_8511),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_8702)
);

INVx5_ASAP7_75t_L g8703 ( 
.A(n_8398),
.Y(n_8703)
);

INVx2_ASAP7_75t_L g8704 ( 
.A(n_8300),
.Y(n_8704)
);

NAND2xp5_ASAP7_75t_SL g8705 ( 
.A(n_8502),
.B(n_8060),
.Y(n_8705)
);

INVx3_ASAP7_75t_L g8706 ( 
.A(n_8329),
.Y(n_8706)
);

NAND2x1_ASAP7_75t_L g8707 ( 
.A(n_8480),
.B(n_893),
.Y(n_8707)
);

NAND2xp5_ASAP7_75t_SL g8708 ( 
.A(n_8061),
.B(n_893),
.Y(n_8708)
);

INVx2_ASAP7_75t_SL g8709 ( 
.A(n_8330),
.Y(n_8709)
);

NAND2xp5_ASAP7_75t_L g8710 ( 
.A(n_8165),
.B(n_29),
.Y(n_8710)
);

NAND2xp5_ASAP7_75t_SL g8711 ( 
.A(n_8063),
.B(n_894),
.Y(n_8711)
);

BUFx2_ASAP7_75t_L g8712 ( 
.A(n_8448),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_8079),
.Y(n_8713)
);

INVx2_ASAP7_75t_SL g8714 ( 
.A(n_8505),
.Y(n_8714)
);

OR2x2_ASAP7_75t_L g8715 ( 
.A(n_8173),
.B(n_8516),
.Y(n_8715)
);

NAND2xp5_ASAP7_75t_L g8716 ( 
.A(n_8249),
.B(n_30),
.Y(n_8716)
);

INVx3_ASAP7_75t_L g8717 ( 
.A(n_8385),
.Y(n_8717)
);

NAND2x1_ASAP7_75t_L g8718 ( 
.A(n_8361),
.B(n_895),
.Y(n_8718)
);

OAI22xp33_ASAP7_75t_L g8719 ( 
.A1(n_8152),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_8719)
);

O2A1O1Ixp33_ASAP7_75t_L g8720 ( 
.A1(n_8103),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_8720)
);

NAND2xp5_ASAP7_75t_SL g8721 ( 
.A(n_8067),
.B(n_8228),
.Y(n_8721)
);

OR2x6_ASAP7_75t_L g8722 ( 
.A(n_8091),
.B(n_895),
.Y(n_8722)
);

AND3x1_ASAP7_75t_SL g8723 ( 
.A(n_8188),
.B(n_31),
.C(n_32),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8086),
.Y(n_8724)
);

AND2x2_ASAP7_75t_L g8725 ( 
.A(n_8160),
.B(n_33),
.Y(n_8725)
);

INVx2_ASAP7_75t_L g8726 ( 
.A(n_8304),
.Y(n_8726)
);

INVx1_ASAP7_75t_L g8727 ( 
.A(n_8105),
.Y(n_8727)
);

NOR3xp33_ASAP7_75t_L g8728 ( 
.A(n_8104),
.B(n_33),
.C(n_34),
.Y(n_8728)
);

AOI22xp5_ASAP7_75t_L g8729 ( 
.A1(n_8507),
.A2(n_8141),
.B1(n_8250),
.B2(n_8247),
.Y(n_8729)
);

AND2x4_ASAP7_75t_L g8730 ( 
.A(n_8386),
.B(n_896),
.Y(n_8730)
);

INVx4_ASAP7_75t_L g8731 ( 
.A(n_8045),
.Y(n_8731)
);

NAND2xp5_ASAP7_75t_L g8732 ( 
.A(n_8094),
.B(n_35),
.Y(n_8732)
);

INVx4_ASAP7_75t_L g8733 ( 
.A(n_8405),
.Y(n_8733)
);

INVx2_ASAP7_75t_SL g8734 ( 
.A(n_8211),
.Y(n_8734)
);

AOI22xp5_ASAP7_75t_L g8735 ( 
.A1(n_8258),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_8735)
);

BUFx6f_ASAP7_75t_L g8736 ( 
.A(n_8224),
.Y(n_8736)
);

AOI22xp33_ASAP7_75t_L g8737 ( 
.A1(n_8527),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_8737)
);

AOI22xp5_ASAP7_75t_L g8738 ( 
.A1(n_8276),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_L g8739 ( 
.A(n_8098),
.B(n_38),
.Y(n_8739)
);

NAND2xp5_ASAP7_75t_L g8740 ( 
.A(n_8101),
.B(n_39),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_L g8741 ( 
.A(n_8133),
.B(n_39),
.Y(n_8741)
);

CKINVDCx20_ASAP7_75t_R g8742 ( 
.A(n_8402),
.Y(n_8742)
);

AND2x2_ASAP7_75t_L g8743 ( 
.A(n_8203),
.B(n_40),
.Y(n_8743)
);

INVx2_ASAP7_75t_L g8744 ( 
.A(n_8312),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_L g8745 ( 
.A(n_8134),
.B(n_40),
.Y(n_8745)
);

CKINVDCx5p33_ASAP7_75t_R g8746 ( 
.A(n_8521),
.Y(n_8746)
);

NAND2xp5_ASAP7_75t_L g8747 ( 
.A(n_8143),
.B(n_8127),
.Y(n_8747)
);

BUFx3_ASAP7_75t_L g8748 ( 
.A(n_8226),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_8315),
.Y(n_8749)
);

BUFx2_ASAP7_75t_L g8750 ( 
.A(n_8229),
.Y(n_8750)
);

INVx2_ASAP7_75t_L g8751 ( 
.A(n_8399),
.Y(n_8751)
);

INVx3_ASAP7_75t_L g8752 ( 
.A(n_8391),
.Y(n_8752)
);

HB1xp67_ASAP7_75t_L g8753 ( 
.A(n_8368),
.Y(n_8753)
);

AND2x4_ASAP7_75t_L g8754 ( 
.A(n_8236),
.B(n_896),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_8107),
.Y(n_8755)
);

OR2x4_ASAP7_75t_L g8756 ( 
.A(n_8157),
.B(n_40),
.Y(n_8756)
);

INVx2_ASAP7_75t_L g8757 ( 
.A(n_8400),
.Y(n_8757)
);

INVx1_ASAP7_75t_L g8758 ( 
.A(n_8122),
.Y(n_8758)
);

INVx8_ASAP7_75t_L g8759 ( 
.A(n_8345),
.Y(n_8759)
);

INVx4_ASAP7_75t_L g8760 ( 
.A(n_8266),
.Y(n_8760)
);

INVx2_ASAP7_75t_SL g8761 ( 
.A(n_8273),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_8144),
.Y(n_8762)
);

INVx2_ASAP7_75t_SL g8763 ( 
.A(n_8287),
.Y(n_8763)
);

INVx1_ASAP7_75t_L g8764 ( 
.A(n_8145),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_L g8765 ( 
.A(n_8317),
.B(n_41),
.Y(n_8765)
);

AND2x4_ASAP7_75t_L g8766 ( 
.A(n_8305),
.B(n_897),
.Y(n_8766)
);

NAND2xp5_ASAP7_75t_L g8767 ( 
.A(n_8355),
.B(n_41),
.Y(n_8767)
);

INVx1_ASAP7_75t_L g8768 ( 
.A(n_8147),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_SL g8769 ( 
.A(n_8284),
.B(n_897),
.Y(n_8769)
);

AND2x4_ASAP7_75t_L g8770 ( 
.A(n_8322),
.B(n_8428),
.Y(n_8770)
);

NOR2xp33_ASAP7_75t_L g8771 ( 
.A(n_8090),
.B(n_898),
.Y(n_8771)
);

NAND2xp5_ASAP7_75t_L g8772 ( 
.A(n_8364),
.B(n_41),
.Y(n_8772)
);

AOI22xp33_ASAP7_75t_L g8773 ( 
.A1(n_8243),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_8773)
);

INVx1_ASAP7_75t_L g8774 ( 
.A(n_8163),
.Y(n_8774)
);

AO22x1_ASAP7_75t_L g8775 ( 
.A1(n_8286),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_8775)
);

NOR3xp33_ASAP7_75t_SL g8776 ( 
.A(n_8499),
.B(n_42),
.C(n_43),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_SL g8777 ( 
.A(n_8302),
.B(n_898),
.Y(n_8777)
);

AOI22xp33_ASAP7_75t_L g8778 ( 
.A1(n_8130),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_8778)
);

NAND2xp5_ASAP7_75t_L g8779 ( 
.A(n_8132),
.B(n_45),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_L g8780 ( 
.A(n_8349),
.B(n_45),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_8182),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_L g8782 ( 
.A(n_8375),
.B(n_46),
.Y(n_8782)
);

INVx1_ASAP7_75t_L g8783 ( 
.A(n_8193),
.Y(n_8783)
);

BUFx3_ASAP7_75t_L g8784 ( 
.A(n_8340),
.Y(n_8784)
);

INVx3_ASAP7_75t_L g8785 ( 
.A(n_8461),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_8216),
.Y(n_8786)
);

BUFx2_ASAP7_75t_L g8787 ( 
.A(n_8363),
.Y(n_8787)
);

INVx1_ASAP7_75t_L g8788 ( 
.A(n_8242),
.Y(n_8788)
);

INVx5_ASAP7_75t_L g8789 ( 
.A(n_8221),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_8389),
.B(n_46),
.Y(n_8790)
);

OR2x2_ASAP7_75t_L g8791 ( 
.A(n_8267),
.B(n_899),
.Y(n_8791)
);

INVx4_ASAP7_75t_L g8792 ( 
.A(n_8363),
.Y(n_8792)
);

NAND2xp5_ASAP7_75t_SL g8793 ( 
.A(n_8319),
.B(n_900),
.Y(n_8793)
);

INVx1_ASAP7_75t_L g8794 ( 
.A(n_8244),
.Y(n_8794)
);

OAI22xp5_ASAP7_75t_SL g8795 ( 
.A1(n_8457),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_8795)
);

A2O1A1Ixp33_ASAP7_75t_L g8796 ( 
.A1(n_8431),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_8796)
);

INVx1_ASAP7_75t_L g8797 ( 
.A(n_8254),
.Y(n_8797)
);

INVx2_ASAP7_75t_L g8798 ( 
.A(n_8409),
.Y(n_8798)
);

CKINVDCx5p33_ASAP7_75t_R g8799 ( 
.A(n_8414),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_8259),
.Y(n_8800)
);

NAND2x1p5_ASAP7_75t_L g8801 ( 
.A(n_8043),
.B(n_900),
.Y(n_8801)
);

NAND2xp5_ASAP7_75t_L g8802 ( 
.A(n_8136),
.B(n_48),
.Y(n_8802)
);

NOR2xp33_ASAP7_75t_L g8803 ( 
.A(n_8277),
.B(n_901),
.Y(n_8803)
);

INVx5_ASAP7_75t_L g8804 ( 
.A(n_8221),
.Y(n_8804)
);

NAND2xp5_ASAP7_75t_L g8805 ( 
.A(n_8215),
.B(n_50),
.Y(n_8805)
);

BUFx2_ASAP7_75t_L g8806 ( 
.A(n_8084),
.Y(n_8806)
);

INVx5_ASAP7_75t_L g8807 ( 
.A(n_8167),
.Y(n_8807)
);

NAND2xp5_ASAP7_75t_L g8808 ( 
.A(n_8223),
.B(n_50),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_8320),
.B(n_50),
.Y(n_8809)
);

AOI22xp33_ASAP7_75t_L g8810 ( 
.A1(n_8274),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_8810)
);

BUFx6f_ASAP7_75t_L g8811 ( 
.A(n_8241),
.Y(n_8811)
);

BUFx3_ASAP7_75t_L g8812 ( 
.A(n_8406),
.Y(n_8812)
);

BUFx2_ASAP7_75t_L g8813 ( 
.A(n_8460),
.Y(n_8813)
);

NAND2xp5_ASAP7_75t_SL g8814 ( 
.A(n_8454),
.B(n_901),
.Y(n_8814)
);

NAND2xp5_ASAP7_75t_SL g8815 ( 
.A(n_8159),
.B(n_902),
.Y(n_8815)
);

NAND2xp5_ASAP7_75t_L g8816 ( 
.A(n_8174),
.B(n_51),
.Y(n_8816)
);

INVx1_ASAP7_75t_L g8817 ( 
.A(n_8262),
.Y(n_8817)
);

NOR3xp33_ASAP7_75t_L g8818 ( 
.A(n_8453),
.B(n_51),
.C(n_52),
.Y(n_8818)
);

NAND2xp5_ASAP7_75t_SL g8819 ( 
.A(n_8416),
.B(n_903),
.Y(n_8819)
);

BUFx6f_ASAP7_75t_L g8820 ( 
.A(n_8024),
.Y(n_8820)
);

BUFx6f_ASAP7_75t_L g8821 ( 
.A(n_8039),
.Y(n_8821)
);

INVx4_ASAP7_75t_L g8822 ( 
.A(n_8227),
.Y(n_8822)
);

NAND2xp5_ASAP7_75t_L g8823 ( 
.A(n_8494),
.B(n_52),
.Y(n_8823)
);

BUFx2_ASAP7_75t_L g8824 ( 
.A(n_8471),
.Y(n_8824)
);

NAND2xp5_ASAP7_75t_L g8825 ( 
.A(n_8366),
.B(n_8439),
.Y(n_8825)
);

NAND2xp5_ASAP7_75t_L g8826 ( 
.A(n_8121),
.B(n_53),
.Y(n_8826)
);

AO22x1_ASAP7_75t_L g8827 ( 
.A1(n_8345),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_8827)
);

INVx2_ASAP7_75t_SL g8828 ( 
.A(n_8455),
.Y(n_8828)
);

INVxp67_ASAP7_75t_L g8829 ( 
.A(n_8336),
.Y(n_8829)
);

AOI22xp33_ASAP7_75t_L g8830 ( 
.A1(n_8404),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_8830)
);

AND2x2_ASAP7_75t_L g8831 ( 
.A(n_8495),
.B(n_54),
.Y(n_8831)
);

NAND2xp5_ASAP7_75t_L g8832 ( 
.A(n_8212),
.B(n_55),
.Y(n_8832)
);

INVx2_ASAP7_75t_SL g8833 ( 
.A(n_8062),
.Y(n_8833)
);

OR2x2_ASAP7_75t_SL g8834 ( 
.A(n_8440),
.B(n_56),
.Y(n_8834)
);

INVx1_ASAP7_75t_L g8835 ( 
.A(n_8269),
.Y(n_8835)
);

AOI22xp5_ASAP7_75t_L g8836 ( 
.A1(n_8433),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_8836)
);

NAND2xp5_ASAP7_75t_SL g8837 ( 
.A(n_8423),
.B(n_903),
.Y(n_8837)
);

CKINVDCx5p33_ASAP7_75t_R g8838 ( 
.A(n_8306),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_8339),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_L g8840 ( 
.A(n_8383),
.B(n_57),
.Y(n_8840)
);

INVx1_ASAP7_75t_L g8841 ( 
.A(n_8341),
.Y(n_8841)
);

AND2x4_ASAP7_75t_L g8842 ( 
.A(n_8501),
.B(n_904),
.Y(n_8842)
);

AOI22xp33_ASAP7_75t_L g8843 ( 
.A1(n_8404),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_8843)
);

NAND2xp5_ASAP7_75t_L g8844 ( 
.A(n_8410),
.B(n_60),
.Y(n_8844)
);

INVx1_ASAP7_75t_L g8845 ( 
.A(n_8347),
.Y(n_8845)
);

AOI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_8140),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_8846)
);

AOI22xp5_ASAP7_75t_L g8847 ( 
.A1(n_8118),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_8847)
);

NAND2xp5_ASAP7_75t_L g8848 ( 
.A(n_8412),
.B(n_61),
.Y(n_8848)
);

AOI22xp33_ASAP7_75t_L g8849 ( 
.A1(n_8404),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_8849)
);

INVx4_ASAP7_75t_L g8850 ( 
.A(n_8408),
.Y(n_8850)
);

INVx2_ASAP7_75t_L g8851 ( 
.A(n_8425),
.Y(n_8851)
);

INVx2_ASAP7_75t_L g8852 ( 
.A(n_8434),
.Y(n_8852)
);

NAND2xp5_ASAP7_75t_SL g8853 ( 
.A(n_8280),
.B(n_904),
.Y(n_8853)
);

NAND2xp5_ASAP7_75t_L g8854 ( 
.A(n_8426),
.B(n_63),
.Y(n_8854)
);

OAI221xp5_ASAP7_75t_L g8855 ( 
.A1(n_8318),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_8855)
);

AND2x2_ASAP7_75t_L g8856 ( 
.A(n_8268),
.B(n_64),
.Y(n_8856)
);

INVx4_ASAP7_75t_L g8857 ( 
.A(n_8408),
.Y(n_8857)
);

INVxp67_ASAP7_75t_L g8858 ( 
.A(n_8352),
.Y(n_8858)
);

INVx1_ASAP7_75t_L g8859 ( 
.A(n_8353),
.Y(n_8859)
);

NAND2xp5_ASAP7_75t_SL g8860 ( 
.A(n_8482),
.B(n_905),
.Y(n_8860)
);

INVx3_ASAP7_75t_L g8861 ( 
.A(n_8390),
.Y(n_8861)
);

BUFx3_ASAP7_75t_L g8862 ( 
.A(n_8487),
.Y(n_8862)
);

BUFx2_ASAP7_75t_L g8863 ( 
.A(n_8360),
.Y(n_8863)
);

OR2x6_ASAP7_75t_L g8864 ( 
.A(n_8415),
.B(n_905),
.Y(n_8864)
);

INVx3_ASAP7_75t_L g8865 ( 
.A(n_8451),
.Y(n_8865)
);

NAND2xp5_ASAP7_75t_L g8866 ( 
.A(n_8459),
.B(n_65),
.Y(n_8866)
);

INVx2_ASAP7_75t_L g8867 ( 
.A(n_8469),
.Y(n_8867)
);

AND2x2_ASAP7_75t_L g8868 ( 
.A(n_8288),
.B(n_65),
.Y(n_8868)
);

INVx1_ASAP7_75t_L g8869 ( 
.A(n_8523),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_8530),
.Y(n_8870)
);

NAND2xp5_ASAP7_75t_SL g8871 ( 
.A(n_8482),
.B(n_906),
.Y(n_8871)
);

INVx5_ASAP7_75t_L g8872 ( 
.A(n_8421),
.Y(n_8872)
);

NAND2xp5_ASAP7_75t_L g8873 ( 
.A(n_8478),
.B(n_66),
.Y(n_8873)
);

A2O1A1Ixp33_ASAP7_75t_L g8874 ( 
.A1(n_8253),
.A2(n_8489),
.B(n_8272),
.C(n_8358),
.Y(n_8874)
);

INVx3_ASAP7_75t_L g8875 ( 
.A(n_8450),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_L g8876 ( 
.A(n_8113),
.B(n_66),
.Y(n_8876)
);

INVx1_ASAP7_75t_L g8877 ( 
.A(n_8496),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_SL g8878 ( 
.A(n_8482),
.B(n_8397),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_8498),
.Y(n_8879)
);

INVx1_ASAP7_75t_L g8880 ( 
.A(n_8407),
.Y(n_8880)
);

INVx5_ASAP7_75t_L g8881 ( 
.A(n_8421),
.Y(n_8881)
);

NAND2xp5_ASAP7_75t_SL g8882 ( 
.A(n_8482),
.B(n_906),
.Y(n_8882)
);

AND2x2_ASAP7_75t_SL g8883 ( 
.A(n_8171),
.B(n_907),
.Y(n_8883)
);

AND2x4_ASAP7_75t_L g8884 ( 
.A(n_8282),
.B(n_8291),
.Y(n_8884)
);

AOI22xp33_ASAP7_75t_L g8885 ( 
.A1(n_8124),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_8885)
);

INVx2_ASAP7_75t_SL g8886 ( 
.A(n_8289),
.Y(n_8886)
);

NAND2xp5_ASAP7_75t_SL g8887 ( 
.A(n_8071),
.B(n_909),
.Y(n_8887)
);

NAND2xp5_ASAP7_75t_L g8888 ( 
.A(n_8137),
.B(n_67),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8470),
.Y(n_8889)
);

INVx2_ASAP7_75t_L g8890 ( 
.A(n_8295),
.Y(n_8890)
);

AND2x6_ASAP7_75t_L g8891 ( 
.A(n_8292),
.B(n_909),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_8492),
.Y(n_8892)
);

OR2x6_ASAP7_75t_L g8893 ( 
.A(n_8110),
.B(n_910),
.Y(n_8893)
);

INVx5_ASAP7_75t_L g8894 ( 
.A(n_8321),
.Y(n_8894)
);

NAND3xp33_ASAP7_75t_SL g8895 ( 
.A(n_8142),
.B(n_68),
.C(n_69),
.Y(n_8895)
);

NAND2xp5_ASAP7_75t_L g8896 ( 
.A(n_8393),
.B(n_68),
.Y(n_8896)
);

AOI22xp5_ASAP7_75t_L g8897 ( 
.A1(n_8148),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_8897)
);

INVxp67_ASAP7_75t_L g8898 ( 
.A(n_8359),
.Y(n_8898)
);

NAND2xp5_ASAP7_75t_SL g8899 ( 
.A(n_8508),
.B(n_910),
.Y(n_8899)
);

BUFx6f_ASAP7_75t_L g8900 ( 
.A(n_8301),
.Y(n_8900)
);

INVx3_ASAP7_75t_L g8901 ( 
.A(n_8372),
.Y(n_8901)
);

INVx2_ASAP7_75t_L g8902 ( 
.A(n_8376),
.Y(n_8902)
);

INVx1_ASAP7_75t_L g8903 ( 
.A(n_8380),
.Y(n_8903)
);

NAND2xp5_ASAP7_75t_L g8904 ( 
.A(n_8394),
.B(n_70),
.Y(n_8904)
);

OAI21xp5_ASAP7_75t_L g8905 ( 
.A1(n_8510),
.A2(n_71),
.B(n_72),
.Y(n_8905)
);

CKINVDCx5p33_ASAP7_75t_R g8906 ( 
.A(n_8195),
.Y(n_8906)
);

NAND2xp5_ASAP7_75t_L g8907 ( 
.A(n_8522),
.B(n_71),
.Y(n_8907)
);

AND2x4_ASAP7_75t_L g8908 ( 
.A(n_8382),
.B(n_911),
.Y(n_8908)
);

INVxp67_ASAP7_75t_L g8909 ( 
.A(n_8463),
.Y(n_8909)
);

INVx5_ASAP7_75t_L g8910 ( 
.A(n_8351),
.Y(n_8910)
);

NOR2xp33_ASAP7_75t_L g8911 ( 
.A(n_8239),
.B(n_911),
.Y(n_8911)
);

INVx1_ASAP7_75t_L g8912 ( 
.A(n_8387),
.Y(n_8912)
);

INVx1_ASAP7_75t_L g8913 ( 
.A(n_8413),
.Y(n_8913)
);

HB1xp67_ASAP7_75t_L g8914 ( 
.A(n_8418),
.Y(n_8914)
);

BUFx4f_ASAP7_75t_L g8915 ( 
.A(n_8373),
.Y(n_8915)
);

AOI22xp5_ASAP7_75t_L g8916 ( 
.A1(n_8422),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_8916)
);

AOI21xp33_ASAP7_75t_L g8917 ( 
.A1(n_8411),
.A2(n_73),
.B(n_74),
.Y(n_8917)
);

NOR2xp33_ASAP7_75t_L g8918 ( 
.A(n_8379),
.B(n_912),
.Y(n_8918)
);

BUFx2_ASAP7_75t_R g8919 ( 
.A(n_8377),
.Y(n_8919)
);

AOI22xp33_ASAP7_75t_L g8920 ( 
.A1(n_8278),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_8920)
);

INVx2_ASAP7_75t_L g8921 ( 
.A(n_8420),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_8430),
.Y(n_8922)
);

INVx1_ASAP7_75t_L g8923 ( 
.A(n_8436),
.Y(n_8923)
);

AND2x4_ASAP7_75t_L g8924 ( 
.A(n_8438),
.B(n_912),
.Y(n_8924)
);

INVx1_ASAP7_75t_L g8925 ( 
.A(n_8464),
.Y(n_8925)
);

INVx1_ASAP7_75t_L g8926 ( 
.A(n_8466),
.Y(n_8926)
);

NOR2xp33_ASAP7_75t_L g8927 ( 
.A(n_8445),
.B(n_914),
.Y(n_8927)
);

NOR2x2_ASAP7_75t_L g8928 ( 
.A(n_8481),
.B(n_8337),
.Y(n_8928)
);

AO22x1_ASAP7_75t_L g8929 ( 
.A1(n_8468),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_8929)
);

NOR2xp33_ASAP7_75t_L g8930 ( 
.A(n_8246),
.B(n_914),
.Y(n_8930)
);

INVx2_ASAP7_75t_L g8931 ( 
.A(n_8488),
.Y(n_8931)
);

BUFx8_ASAP7_75t_L g8932 ( 
.A(n_8491),
.Y(n_8932)
);

BUFx12f_ASAP7_75t_L g8933 ( 
.A(n_8232),
.Y(n_8933)
);

INVx2_ASAP7_75t_SL g8934 ( 
.A(n_8256),
.Y(n_8934)
);

CKINVDCx5p33_ASAP7_75t_R g8935 ( 
.A(n_8497),
.Y(n_8935)
);

INVx2_ASAP7_75t_L g8936 ( 
.A(n_8503),
.Y(n_8936)
);

AOI22xp5_ASAP7_75t_L g8937 ( 
.A1(n_8403),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_8937)
);

INVx2_ASAP7_75t_SL g8938 ( 
.A(n_8367),
.Y(n_8938)
);

CKINVDCx20_ASAP7_75t_R g8939 ( 
.A(n_8261),
.Y(n_8939)
);

INVx1_ASAP7_75t_L g8940 ( 
.A(n_8378),
.Y(n_8940)
);

INVx1_ASAP7_75t_L g8941 ( 
.A(n_8381),
.Y(n_8941)
);

AOI22xp5_ASAP7_75t_L g8942 ( 
.A1(n_8526),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_8942)
);

AOI22xp33_ASAP7_75t_L g8943 ( 
.A1(n_8255),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_8943)
);

NOR2xp33_ASAP7_75t_L g8944 ( 
.A(n_8263),
.B(n_915),
.Y(n_8944)
);

CKINVDCx5p33_ASAP7_75t_R g8945 ( 
.A(n_8506),
.Y(n_8945)
);

OAI21xp33_ASAP7_75t_L g8946 ( 
.A1(n_8194),
.A2(n_78),
.B(n_80),
.Y(n_8946)
);

INVx1_ASAP7_75t_L g8947 ( 
.A(n_8395),
.Y(n_8947)
);

NAND3xp33_ASAP7_75t_SL g8948 ( 
.A(n_8088),
.B(n_80),
.C(n_81),
.Y(n_8948)
);

OR2x2_ASAP7_75t_L g8949 ( 
.A(n_8213),
.B(n_915),
.Y(n_8949)
);

AOI22xp33_ASAP7_75t_L g8950 ( 
.A1(n_8222),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_8950)
);

INVx2_ASAP7_75t_L g8951 ( 
.A(n_8307),
.Y(n_8951)
);

NOR2xp33_ASAP7_75t_L g8952 ( 
.A(n_8264),
.B(n_916),
.Y(n_8952)
);

INVxp67_ASAP7_75t_L g8953 ( 
.A(n_8500),
.Y(n_8953)
);

NAND2xp5_ASAP7_75t_L g8954 ( 
.A(n_8175),
.B(n_8176),
.Y(n_8954)
);

NAND2xp5_ASAP7_75t_L g8955 ( 
.A(n_8189),
.B(n_81),
.Y(n_8955)
);

AO22x1_ASAP7_75t_L g8956 ( 
.A1(n_8371),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_8956)
);

NAND2xp5_ASAP7_75t_L g8957 ( 
.A(n_8191),
.B(n_84),
.Y(n_8957)
);

NAND2xp5_ASAP7_75t_L g8958 ( 
.A(n_8199),
.B(n_8200),
.Y(n_8958)
);

BUFx3_ASAP7_75t_L g8959 ( 
.A(n_8219),
.Y(n_8959)
);

CKINVDCx5p33_ASAP7_75t_R g8960 ( 
.A(n_8504),
.Y(n_8960)
);

INVx2_ASAP7_75t_L g8961 ( 
.A(n_8309),
.Y(n_8961)
);

NAND2x1p5_ASAP7_75t_L g8962 ( 
.A(n_8296),
.B(n_8299),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_8396),
.Y(n_8963)
);

AOI22xp5_ASAP7_75t_L g8964 ( 
.A1(n_8477),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_8964)
);

NAND2xp5_ASAP7_75t_L g8965 ( 
.A(n_8207),
.B(n_85),
.Y(n_8965)
);

NOR2xp33_ASAP7_75t_L g8966 ( 
.A(n_8323),
.B(n_917),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_8210),
.B(n_86),
.Y(n_8967)
);

BUFx6f_ASAP7_75t_L g8968 ( 
.A(n_8374),
.Y(n_8968)
);

INVx1_ASAP7_75t_L g8969 ( 
.A(n_8313),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_8325),
.Y(n_8970)
);

NAND2xp5_ASAP7_75t_SL g8971 ( 
.A(n_8219),
.B(n_918),
.Y(n_8971)
);

INVx1_ASAP7_75t_L g8972 ( 
.A(n_8326),
.Y(n_8972)
);

INVx2_ASAP7_75t_SL g8973 ( 
.A(n_8219),
.Y(n_8973)
);

NAND2xp5_ASAP7_75t_L g8974 ( 
.A(n_8214),
.B(n_86),
.Y(n_8974)
);

INVx1_ASAP7_75t_L g8975 ( 
.A(n_8218),
.Y(n_8975)
);

OR2x2_ASAP7_75t_L g8976 ( 
.A(n_8231),
.B(n_918),
.Y(n_8976)
);

CKINVDCx20_ASAP7_75t_R g8977 ( 
.A(n_8490),
.Y(n_8977)
);

NAND2xp5_ASAP7_75t_SL g8978 ( 
.A(n_8219),
.B(n_919),
.Y(n_8978)
);

NAND2xp5_ASAP7_75t_L g8979 ( 
.A(n_8237),
.B(n_87),
.Y(n_8979)
);

NOR2xp33_ASAP7_75t_R g8980 ( 
.A(n_8271),
.B(n_920),
.Y(n_8980)
);

INVx2_ASAP7_75t_L g8981 ( 
.A(n_8252),
.Y(n_8981)
);

BUFx3_ASAP7_75t_L g8982 ( 
.A(n_8248),
.Y(n_8982)
);

AOI21xp5_ASAP7_75t_L g8983 ( 
.A1(n_8462),
.A2(n_921),
.B(n_920),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_8265),
.Y(n_8984)
);

INVx2_ASAP7_75t_L g8985 ( 
.A(n_8275),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_8279),
.Y(n_8986)
);

BUFx2_ASAP7_75t_L g8987 ( 
.A(n_8283),
.Y(n_8987)
);

NAND2xp5_ASAP7_75t_L g8988 ( 
.A(n_8297),
.B(n_88),
.Y(n_8988)
);

INVx1_ASAP7_75t_L g8989 ( 
.A(n_8298),
.Y(n_8989)
);

INVx1_ASAP7_75t_L g8990 ( 
.A(n_8303),
.Y(n_8990)
);

BUFx3_ASAP7_75t_L g8991 ( 
.A(n_8248),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_8332),
.Y(n_8992)
);

INVx2_ASAP7_75t_SL g8993 ( 
.A(n_8342),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8343),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_8344),
.Y(n_8995)
);

NAND2xp5_ASAP7_75t_L g8996 ( 
.A(n_8346),
.B(n_89),
.Y(n_8996)
);

AND2x6_ASAP7_75t_L g8997 ( 
.A(n_8248),
.B(n_921),
.Y(n_8997)
);

AND2x2_ASAP7_75t_L g8998 ( 
.A(n_8479),
.B(n_89),
.Y(n_8998)
);

BUFx3_ASAP7_75t_L g8999 ( 
.A(n_8248),
.Y(n_8999)
);

NAND2xp5_ASAP7_75t_SL g9000 ( 
.A(n_8138),
.B(n_922),
.Y(n_9000)
);

INVx1_ASAP7_75t_L g9001 ( 
.A(n_8354),
.Y(n_9001)
);

INVx2_ASAP7_75t_L g9002 ( 
.A(n_8356),
.Y(n_9002)
);

INVx1_ASAP7_75t_L g9003 ( 
.A(n_8357),
.Y(n_9003)
);

INVx3_ASAP7_75t_L g9004 ( 
.A(n_8362),
.Y(n_9004)
);

INVx2_ASAP7_75t_L g9005 ( 
.A(n_8365),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8308),
.Y(n_9006)
);

NAND3xp33_ASAP7_75t_SL g9007 ( 
.A(n_8467),
.B(n_89),
.C(n_90),
.Y(n_9007)
);

BUFx6f_ASAP7_75t_L g9008 ( 
.A(n_8442),
.Y(n_9008)
);

NAND2xp5_ASAP7_75t_L g9009 ( 
.A(n_8419),
.B(n_90),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8486),
.Y(n_9010)
);

BUFx6f_ASAP7_75t_L g9011 ( 
.A(n_8427),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8293),
.Y(n_9012)
);

INVx3_ASAP7_75t_L g9013 ( 
.A(n_8429),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8432),
.Y(n_9014)
);

HB1xp67_ASAP7_75t_L g9015 ( 
.A(n_8437),
.Y(n_9015)
);

INVx3_ASAP7_75t_L g9016 ( 
.A(n_8441),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_8443),
.Y(n_9017)
);

INVxp67_ASAP7_75t_L g9018 ( 
.A(n_8447),
.Y(n_9018)
);

INVx2_ASAP7_75t_L g9019 ( 
.A(n_8452),
.Y(n_9019)
);

NAND2xp5_ASAP7_75t_L g9020 ( 
.A(n_8456),
.B(n_90),
.Y(n_9020)
);

BUFx6f_ASAP7_75t_L g9021 ( 
.A(n_8465),
.Y(n_9021)
);

AOI22xp5_ASAP7_75t_L g9022 ( 
.A1(n_8474),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_9022)
);

INVx2_ASAP7_75t_SL g9023 ( 
.A(n_8472),
.Y(n_9023)
);

INVx2_ASAP7_75t_L g9024 ( 
.A(n_8484),
.Y(n_9024)
);

NOR3xp33_ASAP7_75t_SL g9025 ( 
.A(n_8190),
.B(n_91),
.C(n_92),
.Y(n_9025)
);

CKINVDCx5p33_ASAP7_75t_R g9026 ( 
.A(n_8485),
.Y(n_9026)
);

AND2x4_ASAP7_75t_L g9027 ( 
.A(n_8327),
.B(n_922),
.Y(n_9027)
);

AND2x4_ASAP7_75t_L g9028 ( 
.A(n_8369),
.B(n_923),
.Y(n_9028)
);

NAND2xp5_ASAP7_75t_SL g9029 ( 
.A(n_8186),
.B(n_923),
.Y(n_9029)
);

INVx3_ASAP7_75t_L g9030 ( 
.A(n_8206),
.Y(n_9030)
);

NAND2xp5_ASAP7_75t_L g9031 ( 
.A(n_8035),
.B(n_91),
.Y(n_9031)
);

INVxp67_ASAP7_75t_L g9032 ( 
.A(n_8055),
.Y(n_9032)
);

BUFx2_ASAP7_75t_L g9033 ( 
.A(n_8074),
.Y(n_9033)
);

NOR2xp33_ASAP7_75t_L g9034 ( 
.A(n_8031),
.B(n_924),
.Y(n_9034)
);

AOI22xp33_ASAP7_75t_L g9035 ( 
.A1(n_8035),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_L g9036 ( 
.A(n_8035),
.B(n_93),
.Y(n_9036)
);

NAND2xp5_ASAP7_75t_L g9037 ( 
.A(n_8035),
.B(n_94),
.Y(n_9037)
);

INVx2_ASAP7_75t_SL g9038 ( 
.A(n_8051),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8177),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_8177),
.Y(n_9040)
);

BUFx3_ASAP7_75t_L g9041 ( 
.A(n_8051),
.Y(n_9041)
);

NAND2xp5_ASAP7_75t_L g9042 ( 
.A(n_8035),
.B(n_94),
.Y(n_9042)
);

NAND2xp5_ASAP7_75t_SL g9043 ( 
.A(n_8035),
.B(n_924),
.Y(n_9043)
);

NAND2xp5_ASAP7_75t_L g9044 ( 
.A(n_8035),
.B(n_95),
.Y(n_9044)
);

INVx3_ASAP7_75t_L g9045 ( 
.A(n_8206),
.Y(n_9045)
);

CKINVDCx5p33_ASAP7_75t_R g9046 ( 
.A(n_8392),
.Y(n_9046)
);

BUFx6f_ASAP7_75t_L g9047 ( 
.A(n_8392),
.Y(n_9047)
);

BUFx2_ASAP7_75t_L g9048 ( 
.A(n_8074),
.Y(n_9048)
);

NOR2xp33_ASAP7_75t_R g9049 ( 
.A(n_8057),
.B(n_925),
.Y(n_9049)
);

NAND2xp5_ASAP7_75t_L g9050 ( 
.A(n_8035),
.B(n_95),
.Y(n_9050)
);

NAND2xp5_ASAP7_75t_L g9051 ( 
.A(n_8035),
.B(n_96),
.Y(n_9051)
);

AND3x1_ASAP7_75t_L g9052 ( 
.A(n_8035),
.B(n_96),
.C(n_97),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8177),
.Y(n_9053)
);

NOR2xp33_ASAP7_75t_SL g9054 ( 
.A(n_8135),
.B(n_96),
.Y(n_9054)
);

CKINVDCx5p33_ASAP7_75t_R g9055 ( 
.A(n_8392),
.Y(n_9055)
);

NAND2xp5_ASAP7_75t_L g9056 ( 
.A(n_8035),
.B(n_97),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_8177),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_8177),
.Y(n_9058)
);

INVx2_ASAP7_75t_L g9059 ( 
.A(n_8023),
.Y(n_9059)
);

NOR3xp33_ASAP7_75t_SL g9060 ( 
.A(n_8035),
.B(n_97),
.C(n_98),
.Y(n_9060)
);

AOI22xp5_ASAP7_75t_L g9061 ( 
.A1(n_8035),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_9061)
);

AND2x4_ASAP7_75t_SL g9062 ( 
.A(n_8057),
.B(n_925),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_8177),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_8023),
.Y(n_9064)
);

BUFx3_ASAP7_75t_L g9065 ( 
.A(n_8051),
.Y(n_9065)
);

BUFx8_ASAP7_75t_L g9066 ( 
.A(n_8041),
.Y(n_9066)
);

OR2x2_ASAP7_75t_L g9067 ( 
.A(n_8517),
.B(n_926),
.Y(n_9067)
);

AOI22xp33_ASAP7_75t_L g9068 ( 
.A1(n_8035),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_9068)
);

AOI22xp33_ASAP7_75t_L g9069 ( 
.A1(n_8035),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_9069)
);

AND2x2_ASAP7_75t_SL g9070 ( 
.A(n_8035),
.B(n_926),
.Y(n_9070)
);

AOI22xp5_ASAP7_75t_L g9071 ( 
.A1(n_8035),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8177),
.Y(n_9072)
);

INVx5_ASAP7_75t_L g9073 ( 
.A(n_8051),
.Y(n_9073)
);

NAND2x1p5_ASAP7_75t_L g9074 ( 
.A(n_8281),
.B(n_927),
.Y(n_9074)
);

NAND2xp5_ASAP7_75t_L g9075 ( 
.A(n_8035),
.B(n_102),
.Y(n_9075)
);

INVxp67_ASAP7_75t_L g9076 ( 
.A(n_8055),
.Y(n_9076)
);

INVx2_ASAP7_75t_L g9077 ( 
.A(n_8023),
.Y(n_9077)
);

NOR2xp33_ASAP7_75t_R g9078 ( 
.A(n_8057),
.B(n_927),
.Y(n_9078)
);

NAND2xp5_ASAP7_75t_L g9079 ( 
.A(n_8035),
.B(n_102),
.Y(n_9079)
);

BUFx3_ASAP7_75t_L g9080 ( 
.A(n_8051),
.Y(n_9080)
);

NOR2xp33_ASAP7_75t_L g9081 ( 
.A(n_8031),
.B(n_929),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8177),
.Y(n_9082)
);

NOR2xp33_ASAP7_75t_L g9083 ( 
.A(n_8031),
.B(n_930),
.Y(n_9083)
);

BUFx2_ASAP7_75t_L g9084 ( 
.A(n_8074),
.Y(n_9084)
);

INVx2_ASAP7_75t_L g9085 ( 
.A(n_8023),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_8177),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8177),
.Y(n_9087)
);

AND2x4_ASAP7_75t_SL g9088 ( 
.A(n_8057),
.B(n_930),
.Y(n_9088)
);

BUFx3_ASAP7_75t_L g9089 ( 
.A(n_8051),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_8177),
.Y(n_9090)
);

AND2x4_ASAP7_75t_L g9091 ( 
.A(n_8206),
.B(n_931),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_L g9092 ( 
.A(n_8035),
.B(n_103),
.Y(n_9092)
);

INVx2_ASAP7_75t_L g9093 ( 
.A(n_8023),
.Y(n_9093)
);

NAND2xp5_ASAP7_75t_SL g9094 ( 
.A(n_8035),
.B(n_931),
.Y(n_9094)
);

INVx1_ASAP7_75t_L g9095 ( 
.A(n_8177),
.Y(n_9095)
);

NAND2xp5_ASAP7_75t_SL g9096 ( 
.A(n_8035),
.B(n_932),
.Y(n_9096)
);

INVx3_ASAP7_75t_L g9097 ( 
.A(n_8206),
.Y(n_9097)
);

NAND2xp5_ASAP7_75t_L g9098 ( 
.A(n_8035),
.B(n_103),
.Y(n_9098)
);

NAND2xp5_ASAP7_75t_SL g9099 ( 
.A(n_8035),
.B(n_932),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8177),
.Y(n_9100)
);

NOR2xp67_ASAP7_75t_L g9101 ( 
.A(n_8233),
.B(n_104),
.Y(n_9101)
);

INVx1_ASAP7_75t_L g9102 ( 
.A(n_8177),
.Y(n_9102)
);

INVx1_ASAP7_75t_L g9103 ( 
.A(n_8177),
.Y(n_9103)
);

BUFx6f_ASAP7_75t_L g9104 ( 
.A(n_8392),
.Y(n_9104)
);

NOR2xp33_ASAP7_75t_L g9105 ( 
.A(n_8031),
.B(n_933),
.Y(n_9105)
);

NAND2xp5_ASAP7_75t_SL g9106 ( 
.A(n_8035),
.B(n_933),
.Y(n_9106)
);

INVx2_ASAP7_75t_L g9107 ( 
.A(n_8023),
.Y(n_9107)
);

OR2x6_ASAP7_75t_L g9108 ( 
.A(n_8051),
.B(n_934),
.Y(n_9108)
);

AOI22xp33_ASAP7_75t_L g9109 ( 
.A1(n_8035),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_9109)
);

NOR2xp33_ASAP7_75t_R g9110 ( 
.A(n_8057),
.B(n_936),
.Y(n_9110)
);

AOI21xp5_ASAP7_75t_L g9111 ( 
.A1(n_8553),
.A2(n_937),
.B(n_936),
.Y(n_9111)
);

NOR2x1_ASAP7_75t_L g9112 ( 
.A(n_8539),
.B(n_937),
.Y(n_9112)
);

A2O1A1Ixp33_ASAP7_75t_L g9113 ( 
.A1(n_8582),
.A2(n_8729),
.B(n_9036),
.C(n_9031),
.Y(n_9113)
);

AOI21xp5_ASAP7_75t_L g9114 ( 
.A1(n_8630),
.A2(n_939),
.B(n_938),
.Y(n_9114)
);

NOR2xp33_ASAP7_75t_L g9115 ( 
.A(n_8960),
.B(n_938),
.Y(n_9115)
);

AOI221xp5_ASAP7_75t_L g9116 ( 
.A1(n_8719),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.C(n_107),
.Y(n_9116)
);

NOR2xp33_ASAP7_75t_L g9117 ( 
.A(n_8629),
.B(n_940),
.Y(n_9117)
);

AO32x2_ASAP7_75t_L g9118 ( 
.A1(n_8702),
.A2(n_107),
.A3(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_9118)
);

HB1xp67_ASAP7_75t_L g9119 ( 
.A(n_8712),
.Y(n_9119)
);

NOR2xp33_ASAP7_75t_L g9120 ( 
.A(n_9026),
.B(n_941),
.Y(n_9120)
);

AOI21x1_ASAP7_75t_L g9121 ( 
.A1(n_9010),
.A2(n_9006),
.B(n_8878),
.Y(n_9121)
);

NAND2xp5_ASAP7_75t_SL g9122 ( 
.A(n_8968),
.B(n_941),
.Y(n_9122)
);

AOI21xp5_ASAP7_75t_L g9123 ( 
.A1(n_8874),
.A2(n_943),
.B(n_942),
.Y(n_9123)
);

NAND2xp5_ASAP7_75t_L g9124 ( 
.A(n_8992),
.B(n_942),
.Y(n_9124)
);

BUFx3_ASAP7_75t_L g9125 ( 
.A(n_8633),
.Y(n_9125)
);

AOI21xp33_ASAP7_75t_L g9126 ( 
.A1(n_8534),
.A2(n_108),
.B(n_109),
.Y(n_9126)
);

A2O1A1Ixp33_ASAP7_75t_L g9127 ( 
.A1(n_9037),
.A2(n_946),
.B(n_947),
.C(n_945),
.Y(n_9127)
);

OR2x2_ASAP7_75t_L g9128 ( 
.A(n_8625),
.B(n_945),
.Y(n_9128)
);

O2A1O1Ixp33_ASAP7_75t_L g9129 ( 
.A1(n_8659),
.A2(n_9094),
.B(n_9096),
.C(n_9043),
.Y(n_9129)
);

NAND2xp5_ASAP7_75t_L g9130 ( 
.A(n_8995),
.B(n_947),
.Y(n_9130)
);

NAND2xp5_ASAP7_75t_L g9131 ( 
.A(n_9001),
.B(n_948),
.Y(n_9131)
);

INVx2_ASAP7_75t_L g9132 ( 
.A(n_8548),
.Y(n_9132)
);

NAND2x1p5_ASAP7_75t_L g9133 ( 
.A(n_9073),
.B(n_948),
.Y(n_9133)
);

NOR2x1_ASAP7_75t_L g9134 ( 
.A(n_9101),
.B(n_8639),
.Y(n_9134)
);

NOR2xp33_ASAP7_75t_SL g9135 ( 
.A(n_8577),
.B(n_108),
.Y(n_9135)
);

AND2x2_ASAP7_75t_SL g9136 ( 
.A(n_9070),
.B(n_949),
.Y(n_9136)
);

O2A1O1Ixp33_ASAP7_75t_SL g9137 ( 
.A1(n_9099),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_9137)
);

AOI21xp5_ASAP7_75t_L g9138 ( 
.A1(n_8660),
.A2(n_950),
.B(n_949),
.Y(n_9138)
);

BUFx6f_ASAP7_75t_L g9139 ( 
.A(n_8575),
.Y(n_9139)
);

AO21x1_ASAP7_75t_L g9140 ( 
.A1(n_8654),
.A2(n_110),
.B(n_111),
.Y(n_9140)
);

O2A1O1Ixp33_ASAP7_75t_L g9141 ( 
.A1(n_9106),
.A2(n_113),
.B(n_110),
.C(n_112),
.Y(n_9141)
);

AND2x2_ASAP7_75t_L g9142 ( 
.A(n_9015),
.B(n_950),
.Y(n_9142)
);

OAI21xp5_ASAP7_75t_L g9143 ( 
.A1(n_8561),
.A2(n_8543),
.B(n_8542),
.Y(n_9143)
);

NAND2x1p5_ASAP7_75t_L g9144 ( 
.A(n_9073),
.B(n_951),
.Y(n_9144)
);

AOI21xp5_ASAP7_75t_L g9145 ( 
.A1(n_8669),
.A2(n_952),
.B(n_951),
.Y(n_9145)
);

NAND2xp5_ASAP7_75t_L g9146 ( 
.A(n_9003),
.B(n_952),
.Y(n_9146)
);

AOI21xp5_ASAP7_75t_L g9147 ( 
.A1(n_8954),
.A2(n_8958),
.B(n_8747),
.Y(n_9147)
);

AO32x1_ASAP7_75t_L g9148 ( 
.A1(n_8574),
.A2(n_114),
.A3(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_9148)
);

AND2x2_ASAP7_75t_L g9149 ( 
.A(n_8938),
.B(n_954),
.Y(n_9149)
);

OAI22xp5_ASAP7_75t_L g9150 ( 
.A1(n_8593),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_9150)
);

NOR2xp33_ASAP7_75t_L g9151 ( 
.A(n_8829),
.B(n_8858),
.Y(n_9151)
);

BUFx3_ASAP7_75t_L g9152 ( 
.A(n_8656),
.Y(n_9152)
);

AOI21xp5_ASAP7_75t_L g9153 ( 
.A1(n_8638),
.A2(n_955),
.B(n_954),
.Y(n_9153)
);

OAI22xp5_ASAP7_75t_L g9154 ( 
.A1(n_9042),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_9154)
);

AOI21xp5_ASAP7_75t_L g9155 ( 
.A1(n_9012),
.A2(n_956),
.B(n_955),
.Y(n_9155)
);

NOR2xp67_ASAP7_75t_SL g9156 ( 
.A(n_8894),
.B(n_116),
.Y(n_9156)
);

O2A1O1Ixp33_ASAP7_75t_L g9157 ( 
.A1(n_8769),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_8914),
.Y(n_9158)
);

OAI22xp5_ASAP7_75t_L g9159 ( 
.A1(n_9044),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_9159)
);

INVx2_ASAP7_75t_SL g9160 ( 
.A(n_8575),
.Y(n_9160)
);

AOI22xp5_ASAP7_75t_L g9161 ( 
.A1(n_8579),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_9161)
);

OAI21xp5_ASAP7_75t_L g9162 ( 
.A1(n_8636),
.A2(n_120),
.B(n_121),
.Y(n_9162)
);

AND2x2_ASAP7_75t_L g9163 ( 
.A(n_8884),
.B(n_957),
.Y(n_9163)
);

INVx2_ASAP7_75t_SL g9164 ( 
.A(n_8647),
.Y(n_9164)
);

OAI21xp5_ASAP7_75t_L g9165 ( 
.A1(n_8592),
.A2(n_120),
.B(n_122),
.Y(n_9165)
);

NAND2xp5_ASAP7_75t_L g9166 ( 
.A(n_8545),
.B(n_957),
.Y(n_9166)
);

AND2x2_ASAP7_75t_L g9167 ( 
.A(n_8987),
.B(n_8968),
.Y(n_9167)
);

OAI22xp5_ASAP7_75t_L g9168 ( 
.A1(n_9050),
.A2(n_9056),
.B1(n_9075),
.B2(n_9051),
.Y(n_9168)
);

NOR2xp33_ASAP7_75t_L g9169 ( 
.A(n_8898),
.B(n_958),
.Y(n_9169)
);

OAI22xp5_ASAP7_75t_L g9170 ( 
.A1(n_9079),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_9170)
);

INVxp67_ASAP7_75t_L g9171 ( 
.A(n_8665),
.Y(n_9171)
);

NAND2xp5_ASAP7_75t_L g9172 ( 
.A(n_8556),
.B(n_959),
.Y(n_9172)
);

AOI21xp5_ASAP7_75t_L g9173 ( 
.A1(n_9039),
.A2(n_961),
.B(n_959),
.Y(n_9173)
);

INVxp67_ASAP7_75t_L g9174 ( 
.A(n_8578),
.Y(n_9174)
);

BUFx2_ASAP7_75t_L g9175 ( 
.A(n_9033),
.Y(n_9175)
);

AOI22xp5_ASAP7_75t_L g9176 ( 
.A1(n_8911),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_9176)
);

INVx1_ASAP7_75t_L g9177 ( 
.A(n_8679),
.Y(n_9177)
);

NAND2xp5_ASAP7_75t_L g9178 ( 
.A(n_9040),
.B(n_961),
.Y(n_9178)
);

AOI21xp5_ASAP7_75t_L g9179 ( 
.A1(n_9053),
.A2(n_963),
.B(n_962),
.Y(n_9179)
);

AND2x2_ASAP7_75t_L g9180 ( 
.A(n_8998),
.B(n_962),
.Y(n_9180)
);

BUFx3_ASAP7_75t_L g9181 ( 
.A(n_8616),
.Y(n_9181)
);

NAND2xp5_ASAP7_75t_L g9182 ( 
.A(n_9057),
.B(n_963),
.Y(n_9182)
);

AOI21xp5_ASAP7_75t_L g9183 ( 
.A1(n_9058),
.A2(n_965),
.B(n_964),
.Y(n_9183)
);

AO21x1_ASAP7_75t_L g9184 ( 
.A1(n_9092),
.A2(n_9098),
.B(n_8905),
.Y(n_9184)
);

INVxp67_ASAP7_75t_L g9185 ( 
.A(n_9048),
.Y(n_9185)
);

NAND2xp5_ASAP7_75t_SL g9186 ( 
.A(n_9011),
.B(n_964),
.Y(n_9186)
);

NAND2x1p5_ASAP7_75t_L g9187 ( 
.A(n_8703),
.B(n_965),
.Y(n_9187)
);

AOI21xp5_ASAP7_75t_L g9188 ( 
.A1(n_9063),
.A2(n_967),
.B(n_966),
.Y(n_9188)
);

NAND2xp5_ASAP7_75t_L g9189 ( 
.A(n_9072),
.B(n_966),
.Y(n_9189)
);

AOI21xp5_ASAP7_75t_L g9190 ( 
.A1(n_9082),
.A2(n_968),
.B(n_967),
.Y(n_9190)
);

AO21x1_ASAP7_75t_L g9191 ( 
.A1(n_8585),
.A2(n_123),
.B(n_124),
.Y(n_9191)
);

OR2x2_ASAP7_75t_L g9192 ( 
.A(n_8863),
.B(n_968),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_9086),
.B(n_9087),
.Y(n_9193)
);

NAND2xp5_ASAP7_75t_L g9194 ( 
.A(n_9090),
.B(n_969),
.Y(n_9194)
);

NAND2xp5_ASAP7_75t_L g9195 ( 
.A(n_9095),
.B(n_969),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_9100),
.B(n_970),
.Y(n_9196)
);

AOI21x1_ASAP7_75t_L g9197 ( 
.A1(n_8860),
.A2(n_125),
.B(n_126),
.Y(n_9197)
);

NOR2x1_ASAP7_75t_L g9198 ( 
.A(n_9004),
.B(n_970),
.Y(n_9198)
);

NAND2xp5_ASAP7_75t_L g9199 ( 
.A(n_9102),
.B(n_971),
.Y(n_9199)
);

INVx1_ASAP7_75t_L g9200 ( 
.A(n_8680),
.Y(n_9200)
);

INVx2_ASAP7_75t_L g9201 ( 
.A(n_8549),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8686),
.Y(n_9202)
);

AO32x1_ASAP7_75t_L g9203 ( 
.A1(n_8993),
.A2(n_128),
.A3(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_9203)
);

AOI21xp5_ASAP7_75t_L g9204 ( 
.A1(n_9103),
.A2(n_972),
.B(n_971),
.Y(n_9204)
);

INVx2_ASAP7_75t_L g9205 ( 
.A(n_8554),
.Y(n_9205)
);

NOR2xp33_ASAP7_75t_L g9206 ( 
.A(n_8721),
.B(n_972),
.Y(n_9206)
);

OAI321xp33_ASAP7_75t_L g9207 ( 
.A1(n_8855),
.A2(n_129),
.A3(n_131),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_9207)
);

AOI21xp5_ASAP7_75t_L g9208 ( 
.A1(n_8981),
.A2(n_974),
.B(n_973),
.Y(n_9208)
);

INVx1_ASAP7_75t_L g9209 ( 
.A(n_8688),
.Y(n_9209)
);

A2O1A1Ixp33_ASAP7_75t_L g9210 ( 
.A1(n_8771),
.A2(n_974),
.B(n_975),
.C(n_973),
.Y(n_9210)
);

BUFx4f_ASAP7_75t_L g9211 ( 
.A(n_9047),
.Y(n_9211)
);

AOI21xp5_ASAP7_75t_L g9212 ( 
.A1(n_8985),
.A2(n_977),
.B(n_976),
.Y(n_9212)
);

AO22x1_ASAP7_75t_L g9213 ( 
.A1(n_8894),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_9213)
);

AOI21xp5_ASAP7_75t_L g9214 ( 
.A1(n_8880),
.A2(n_977),
.B(n_976),
.Y(n_9214)
);

NOR2xp33_ASAP7_75t_L g9215 ( 
.A(n_8945),
.B(n_978),
.Y(n_9215)
);

INVx4_ASAP7_75t_L g9216 ( 
.A(n_8663),
.Y(n_9216)
);

NOR2xp33_ASAP7_75t_L g9217 ( 
.A(n_8935),
.B(n_8953),
.Y(n_9217)
);

AOI21xp5_ASAP7_75t_L g9218 ( 
.A1(n_8889),
.A2(n_979),
.B(n_978),
.Y(n_9218)
);

OAI21x1_ASAP7_75t_L g9219 ( 
.A1(n_8903),
.A2(n_130),
.B(n_132),
.Y(n_9219)
);

NAND3xp33_ASAP7_75t_L g9220 ( 
.A(n_8624),
.B(n_130),
.C(n_132),
.Y(n_9220)
);

AND2x2_ASAP7_75t_SL g9221 ( 
.A(n_9052),
.B(n_979),
.Y(n_9221)
);

INVx2_ASAP7_75t_L g9222 ( 
.A(n_8559),
.Y(n_9222)
);

OAI321xp33_ASAP7_75t_L g9223 ( 
.A1(n_8795),
.A2(n_134),
.A3(n_136),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_9223)
);

INVx2_ASAP7_75t_L g9224 ( 
.A(n_8588),
.Y(n_9224)
);

INVx2_ASAP7_75t_L g9225 ( 
.A(n_8614),
.Y(n_9225)
);

NAND2x1_ASAP7_75t_L g9226 ( 
.A(n_8973),
.B(n_980),
.Y(n_9226)
);

AOI21xp5_ASAP7_75t_L g9227 ( 
.A1(n_8892),
.A2(n_981),
.B(n_980),
.Y(n_9227)
);

NAND2xp5_ASAP7_75t_L g9228 ( 
.A(n_8940),
.B(n_981),
.Y(n_9228)
);

AOI21xp5_ASAP7_75t_L g9229 ( 
.A1(n_8951),
.A2(n_983),
.B(n_982),
.Y(n_9229)
);

NAND2xp5_ASAP7_75t_L g9230 ( 
.A(n_8941),
.B(n_984),
.Y(n_9230)
);

OAI21xp33_ASAP7_75t_L g9231 ( 
.A1(n_8780),
.A2(n_133),
.B(n_134),
.Y(n_9231)
);

INVx5_ASAP7_75t_L g9232 ( 
.A(n_8997),
.Y(n_9232)
);

OAI21x1_ASAP7_75t_L g9233 ( 
.A1(n_8912),
.A2(n_133),
.B(n_134),
.Y(n_9233)
);

NAND2xp5_ASAP7_75t_L g9234 ( 
.A(n_8947),
.B(n_985),
.Y(n_9234)
);

AOI21xp5_ASAP7_75t_L g9235 ( 
.A1(n_8961),
.A2(n_987),
.B(n_986),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_8690),
.Y(n_9236)
);

AOI21xp5_ASAP7_75t_L g9237 ( 
.A1(n_8705),
.A2(n_8970),
.B(n_8969),
.Y(n_9237)
);

AOI21xp5_ASAP7_75t_L g9238 ( 
.A1(n_8972),
.A2(n_987),
.B(n_986),
.Y(n_9238)
);

A2O1A1Ixp33_ASAP7_75t_L g9239 ( 
.A1(n_8533),
.A2(n_989),
.B(n_990),
.C(n_988),
.Y(n_9239)
);

NAND2xp5_ASAP7_75t_SL g9240 ( 
.A(n_9011),
.B(n_988),
.Y(n_9240)
);

NAND2xp5_ASAP7_75t_L g9241 ( 
.A(n_8963),
.B(n_989),
.Y(n_9241)
);

HB1xp67_ASAP7_75t_L g9242 ( 
.A(n_8551),
.Y(n_9242)
);

BUFx6f_ASAP7_75t_L g9243 ( 
.A(n_8647),
.Y(n_9243)
);

NOR3xp33_ASAP7_75t_L g9244 ( 
.A(n_8895),
.B(n_135),
.C(n_136),
.Y(n_9244)
);

OAI21x1_ASAP7_75t_L g9245 ( 
.A1(n_8913),
.A2(n_135),
.B(n_137),
.Y(n_9245)
);

OAI21xp5_ASAP7_75t_L g9246 ( 
.A1(n_8599),
.A2(n_137),
.B(n_138),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8699),
.Y(n_9247)
);

NAND2xp5_ASAP7_75t_L g9248 ( 
.A(n_8975),
.B(n_991),
.Y(n_9248)
);

NAND2xp5_ASAP7_75t_L g9249 ( 
.A(n_8984),
.B(n_991),
.Y(n_9249)
);

AO21x1_ASAP7_75t_L g9250 ( 
.A1(n_8587),
.A2(n_137),
.B(n_138),
.Y(n_9250)
);

AND2x2_ASAP7_75t_SL g9251 ( 
.A(n_8883),
.B(n_8728),
.Y(n_9251)
);

OAI22xp5_ASAP7_75t_L g9252 ( 
.A1(n_8915),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_9252)
);

OAI21xp5_ASAP7_75t_L g9253 ( 
.A1(n_8601),
.A2(n_139),
.B(n_140),
.Y(n_9253)
);

OAI22xp5_ASAP7_75t_L g9254 ( 
.A1(n_9060),
.A2(n_142),
.B1(n_139),
.B2(n_140),
.Y(n_9254)
);

INVx1_ASAP7_75t_L g9255 ( 
.A(n_8713),
.Y(n_9255)
);

AOI21x1_ASAP7_75t_L g9256 ( 
.A1(n_8871),
.A2(n_142),
.B(n_143),
.Y(n_9256)
);

AOI21xp5_ASAP7_75t_L g9257 ( 
.A1(n_8986),
.A2(n_8990),
.B(n_8989),
.Y(n_9257)
);

NAND3xp33_ASAP7_75t_L g9258 ( 
.A(n_8918),
.B(n_142),
.C(n_143),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_8724),
.Y(n_9259)
);

AND2x2_ASAP7_75t_L g9260 ( 
.A(n_9019),
.B(n_992),
.Y(n_9260)
);

A2O1A1Ixp33_ASAP7_75t_L g9261 ( 
.A1(n_8927),
.A2(n_8946),
.B(n_8687),
.C(n_8930),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_9024),
.B(n_992),
.Y(n_9262)
);

AOI21xp5_ASAP7_75t_L g9263 ( 
.A1(n_8994),
.A2(n_994),
.B(n_993),
.Y(n_9263)
);

AOI21x1_ASAP7_75t_L g9264 ( 
.A1(n_8882),
.A2(n_143),
.B(n_144),
.Y(n_9264)
);

NOR2xp33_ASAP7_75t_SL g9265 ( 
.A(n_8600),
.B(n_144),
.Y(n_9265)
);

A2O1A1Ixp33_ASAP7_75t_L g9266 ( 
.A1(n_9061),
.A2(n_994),
.B(n_995),
.C(n_993),
.Y(n_9266)
);

AOI22xp5_ASAP7_75t_L g9267 ( 
.A1(n_8590),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_9267)
);

AOI22xp5_ASAP7_75t_L g9268 ( 
.A1(n_8603),
.A2(n_8793),
.B1(n_8777),
.B2(n_8803),
.Y(n_9268)
);

NAND2xp5_ASAP7_75t_SL g9269 ( 
.A(n_9021),
.B(n_996),
.Y(n_9269)
);

INVx1_ASAP7_75t_SL g9270 ( 
.A(n_8565),
.Y(n_9270)
);

A2O1A1Ixp33_ASAP7_75t_L g9271 ( 
.A1(n_9071),
.A2(n_8952),
.B(n_8966),
.C(n_8944),
.Y(n_9271)
);

INVx1_ASAP7_75t_L g9272 ( 
.A(n_8727),
.Y(n_9272)
);

NOR2xp33_ASAP7_75t_L g9273 ( 
.A(n_9021),
.B(n_996),
.Y(n_9273)
);

NAND2x1_ASAP7_75t_L g9274 ( 
.A(n_8901),
.B(n_8936),
.Y(n_9274)
);

BUFx12f_ASAP7_75t_L g9275 ( 
.A(n_8560),
.Y(n_9275)
);

NAND2xp5_ASAP7_75t_L g9276 ( 
.A(n_9002),
.B(n_997),
.Y(n_9276)
);

AOI21xp5_ASAP7_75t_L g9277 ( 
.A1(n_9005),
.A2(n_999),
.B(n_998),
.Y(n_9277)
);

OR2x6_ASAP7_75t_L g9278 ( 
.A(n_8759),
.B(n_998),
.Y(n_9278)
);

NOR2xp33_ASAP7_75t_L g9279 ( 
.A(n_9018),
.B(n_999),
.Y(n_9279)
);

NAND2xp5_ASAP7_75t_SL g9280 ( 
.A(n_9008),
.B(n_1000),
.Y(n_9280)
);

AOI21xp5_ASAP7_75t_L g9281 ( 
.A1(n_9014),
.A2(n_1001),
.B(n_1000),
.Y(n_9281)
);

AOI21xp5_ASAP7_75t_L g9282 ( 
.A1(n_9017),
.A2(n_1002),
.B(n_1001),
.Y(n_9282)
);

NOR2xp33_ASAP7_75t_L g9283 ( 
.A(n_8825),
.B(n_1003),
.Y(n_9283)
);

NAND2xp5_ASAP7_75t_L g9284 ( 
.A(n_9013),
.B(n_1003),
.Y(n_9284)
);

INVx2_ASAP7_75t_L g9285 ( 
.A(n_8626),
.Y(n_9285)
);

NAND2xp5_ASAP7_75t_L g9286 ( 
.A(n_9016),
.B(n_1004),
.Y(n_9286)
);

AOI21xp33_ASAP7_75t_L g9287 ( 
.A1(n_8555),
.A2(n_145),
.B(n_146),
.Y(n_9287)
);

INVx3_ASAP7_75t_L g9288 ( 
.A(n_8694),
.Y(n_9288)
);

OAI21xp5_ASAP7_75t_L g9289 ( 
.A1(n_8547),
.A2(n_145),
.B(n_146),
.Y(n_9289)
);

AOI21xp5_ASAP7_75t_L g9290 ( 
.A1(n_8536),
.A2(n_9023),
.B(n_8562),
.Y(n_9290)
);

INVx2_ASAP7_75t_L g9291 ( 
.A(n_8637),
.Y(n_9291)
);

NAND2xp5_ASAP7_75t_SL g9292 ( 
.A(n_9008),
.B(n_1004),
.Y(n_9292)
);

AOI21xp5_ASAP7_75t_L g9293 ( 
.A1(n_8670),
.A2(n_1007),
.B(n_1005),
.Y(n_9293)
);

INVx2_ASAP7_75t_L g9294 ( 
.A(n_8641),
.Y(n_9294)
);

INVx1_ASAP7_75t_L g9295 ( 
.A(n_8755),
.Y(n_9295)
);

INVx2_ASAP7_75t_L g9296 ( 
.A(n_8645),
.Y(n_9296)
);

AOI22xp5_ASAP7_75t_L g9297 ( 
.A1(n_8612),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8715),
.B(n_8620),
.Y(n_9298)
);

NAND2xp5_ASAP7_75t_L g9299 ( 
.A(n_9084),
.B(n_1005),
.Y(n_9299)
);

AOI21xp5_ASAP7_75t_L g9300 ( 
.A1(n_8971),
.A2(n_1009),
.B(n_1008),
.Y(n_9300)
);

AOI21xp5_ASAP7_75t_L g9301 ( 
.A1(n_8978),
.A2(n_8540),
.B(n_8959),
.Y(n_9301)
);

HB1xp67_ASAP7_75t_L g9302 ( 
.A(n_8677),
.Y(n_9302)
);

AOI21xp5_ASAP7_75t_L g9303 ( 
.A1(n_8552),
.A2(n_1009),
.B(n_1008),
.Y(n_9303)
);

AOI21xp5_ASAP7_75t_L g9304 ( 
.A1(n_8982),
.A2(n_1011),
.B(n_1010),
.Y(n_9304)
);

AOI21x1_ASAP7_75t_L g9305 ( 
.A1(n_8853),
.A2(n_147),
.B(n_148),
.Y(n_9305)
);

A2O1A1Ixp33_ASAP7_75t_L g9306 ( 
.A1(n_8809),
.A2(n_1011),
.B(n_1012),
.C(n_1010),
.Y(n_9306)
);

NAND2xp5_ASAP7_75t_L g9307 ( 
.A(n_8586),
.B(n_1012),
.Y(n_9307)
);

O2A1O1Ixp33_ASAP7_75t_L g9308 ( 
.A1(n_9029),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_9308)
);

NAND2xp5_ASAP7_75t_L g9309 ( 
.A(n_9032),
.B(n_1013),
.Y(n_9309)
);

INVx3_ASAP7_75t_L g9310 ( 
.A(n_8694),
.Y(n_9310)
);

OAI21x1_ASAP7_75t_L g9311 ( 
.A1(n_8922),
.A2(n_150),
.B(n_151),
.Y(n_9311)
);

OAI21xp5_ASAP7_75t_L g9312 ( 
.A1(n_8840),
.A2(n_150),
.B(n_151),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_8758),
.Y(n_9313)
);

NOR3xp33_ASAP7_75t_L g9314 ( 
.A(n_9007),
.B(n_151),
.C(n_152),
.Y(n_9314)
);

INVx4_ASAP7_75t_L g9315 ( 
.A(n_8663),
.Y(n_9315)
);

O2A1O1Ixp5_ASAP7_75t_L g9316 ( 
.A1(n_8775),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_9316)
);

OR2x2_ASAP7_75t_L g9317 ( 
.A(n_8902),
.B(n_1013),
.Y(n_9317)
);

A2O1A1Ixp33_ASAP7_75t_L g9318 ( 
.A1(n_8685),
.A2(n_1015),
.B(n_1016),
.C(n_1014),
.Y(n_9318)
);

NOR2x1_ASAP7_75t_L g9319 ( 
.A(n_8991),
.B(n_1014),
.Y(n_9319)
);

BUFx3_ASAP7_75t_L g9320 ( 
.A(n_8550),
.Y(n_9320)
);

INVx3_ASAP7_75t_L g9321 ( 
.A(n_8672),
.Y(n_9321)
);

BUFx6f_ASAP7_75t_L g9322 ( 
.A(n_8672),
.Y(n_9322)
);

NOR2xp33_ASAP7_75t_SL g9323 ( 
.A(n_8838),
.B(n_152),
.Y(n_9323)
);

BUFx6f_ASAP7_75t_L g9324 ( 
.A(n_8736),
.Y(n_9324)
);

A2O1A1Ixp33_ASAP7_75t_L g9325 ( 
.A1(n_8606),
.A2(n_1017),
.B(n_1018),
.C(n_1016),
.Y(n_9325)
);

NOR2xp33_ASAP7_75t_L g9326 ( 
.A(n_8886),
.B(n_8691),
.Y(n_9326)
);

AOI21xp5_ASAP7_75t_L g9327 ( 
.A1(n_8999),
.A2(n_1018),
.B(n_1017),
.Y(n_9327)
);

INVx2_ASAP7_75t_L g9328 ( 
.A(n_8650),
.Y(n_9328)
);

NAND2xp5_ASAP7_75t_L g9329 ( 
.A(n_9076),
.B(n_1019),
.Y(n_9329)
);

AOI21xp5_ASAP7_75t_L g9330 ( 
.A1(n_8887),
.A2(n_1021),
.B(n_1020),
.Y(n_9330)
);

INVx11_ASAP7_75t_L g9331 ( 
.A(n_9066),
.Y(n_9331)
);

AND2x6_ASAP7_75t_L g9332 ( 
.A(n_8942),
.B(n_1020),
.Y(n_9332)
);

INVx3_ASAP7_75t_L g9333 ( 
.A(n_9030),
.Y(n_9333)
);

NAND2xp5_ASAP7_75t_L g9334 ( 
.A(n_8658),
.B(n_1021),
.Y(n_9334)
);

NOR2xp33_ASAP7_75t_L g9335 ( 
.A(n_8906),
.B(n_1022),
.Y(n_9335)
);

OAI21xp5_ASAP7_75t_L g9336 ( 
.A1(n_8844),
.A2(n_153),
.B(n_154),
.Y(n_9336)
);

AOI21xp5_ASAP7_75t_L g9337 ( 
.A1(n_8546),
.A2(n_1023),
.B(n_1022),
.Y(n_9337)
);

AOI21x1_ASAP7_75t_L g9338 ( 
.A1(n_8899),
.A2(n_8564),
.B(n_8708),
.Y(n_9338)
);

BUFx6f_ASAP7_75t_L g9339 ( 
.A(n_8736),
.Y(n_9339)
);

BUFx6f_ASAP7_75t_L g9340 ( 
.A(n_8557),
.Y(n_9340)
);

NAND2xp5_ASAP7_75t_L g9341 ( 
.A(n_8676),
.B(n_1024),
.Y(n_9341)
);

AOI21xp5_ASAP7_75t_L g9342 ( 
.A1(n_8875),
.A2(n_1025),
.B(n_1024),
.Y(n_9342)
);

AOI21xp5_ASAP7_75t_L g9343 ( 
.A1(n_8796),
.A2(n_1026),
.B(n_1025),
.Y(n_9343)
);

NOR3xp33_ASAP7_75t_L g9344 ( 
.A(n_8948),
.B(n_8854),
.C(n_8848),
.Y(n_9344)
);

NAND2x1p5_ASAP7_75t_L g9345 ( 
.A(n_8703),
.B(n_1028),
.Y(n_9345)
);

NAND2xp5_ASAP7_75t_L g9346 ( 
.A(n_8692),
.B(n_1029),
.Y(n_9346)
);

OR2x2_ASAP7_75t_L g9347 ( 
.A(n_8921),
.B(n_1029),
.Y(n_9347)
);

BUFx12f_ASAP7_75t_L g9348 ( 
.A(n_9046),
.Y(n_9348)
);

NAND2xp5_ASAP7_75t_L g9349 ( 
.A(n_9059),
.B(n_1030),
.Y(n_9349)
);

INVx2_ASAP7_75t_L g9350 ( 
.A(n_9064),
.Y(n_9350)
);

AOI21xp5_ASAP7_75t_L g9351 ( 
.A1(n_8605),
.A2(n_1032),
.B(n_1031),
.Y(n_9351)
);

NOR2xp33_ASAP7_75t_L g9352 ( 
.A(n_8919),
.B(n_1032),
.Y(n_9352)
);

NAND2xp5_ASAP7_75t_L g9353 ( 
.A(n_9077),
.B(n_9085),
.Y(n_9353)
);

AOI21xp5_ASAP7_75t_L g9354 ( 
.A1(n_8751),
.A2(n_1034),
.B(n_1033),
.Y(n_9354)
);

AOI21xp5_ASAP7_75t_L g9355 ( 
.A1(n_8757),
.A2(n_1035),
.B(n_1034),
.Y(n_9355)
);

AOI21xp33_ASAP7_75t_L g9356 ( 
.A1(n_8576),
.A2(n_153),
.B(n_155),
.Y(n_9356)
);

NAND2xp5_ASAP7_75t_L g9357 ( 
.A(n_9093),
.B(n_1035),
.Y(n_9357)
);

NAND2xp5_ASAP7_75t_L g9358 ( 
.A(n_9107),
.B(n_1036),
.Y(n_9358)
);

AOI22xp5_ASAP7_75t_L g9359 ( 
.A1(n_8818),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_8798),
.B(n_1036),
.Y(n_9360)
);

AOI21xp5_ASAP7_75t_L g9361 ( 
.A1(n_8851),
.A2(n_1039),
.B(n_1038),
.Y(n_9361)
);

INVx2_ASAP7_75t_L g9362 ( 
.A(n_8852),
.Y(n_9362)
);

AOI21xp5_ASAP7_75t_L g9363 ( 
.A1(n_8827),
.A2(n_1040),
.B(n_1039),
.Y(n_9363)
);

BUFx8_ASAP7_75t_L g9364 ( 
.A(n_9047),
.Y(n_9364)
);

O2A1O1Ixp33_ASAP7_75t_SL g9365 ( 
.A1(n_8866),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_9365)
);

OA22x2_ASAP7_75t_L g9366 ( 
.A1(n_8608),
.A2(n_159),
.B1(n_156),
.B2(n_158),
.Y(n_9366)
);

NOR2xp33_ASAP7_75t_L g9367 ( 
.A(n_8538),
.B(n_1040),
.Y(n_9367)
);

HB1xp67_ASAP7_75t_L g9368 ( 
.A(n_8824),
.Y(n_9368)
);

OAI22xp5_ASAP7_75t_L g9369 ( 
.A1(n_8806),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_9369)
);

NAND2xp5_ASAP7_75t_SL g9370 ( 
.A(n_8828),
.B(n_1041),
.Y(n_9370)
);

INVx3_ASAP7_75t_L g9371 ( 
.A(n_9045),
.Y(n_9371)
);

OR2x6_ASAP7_75t_L g9372 ( 
.A(n_8759),
.B(n_1041),
.Y(n_9372)
);

O2A1O1Ixp33_ASAP7_75t_L g9373 ( 
.A1(n_8873),
.A2(n_161),
.B(n_158),
.C(n_160),
.Y(n_9373)
);

INVx2_ASAP7_75t_L g9374 ( 
.A(n_8931),
.Y(n_9374)
);

AND2x2_ASAP7_75t_L g9375 ( 
.A(n_8667),
.B(n_1042),
.Y(n_9375)
);

NOR2xp33_ASAP7_75t_L g9376 ( 
.A(n_8977),
.B(n_1042),
.Y(n_9376)
);

NAND2xp5_ASAP7_75t_SL g9377 ( 
.A(n_8980),
.B(n_1043),
.Y(n_9377)
);

AOI21x1_ASAP7_75t_L g9378 ( 
.A1(n_8711),
.A2(n_160),
.B(n_161),
.Y(n_9378)
);

AOI22xp5_ASAP7_75t_L g9379 ( 
.A1(n_8939),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_9379)
);

NOR2xp33_ASAP7_75t_L g9380 ( 
.A(n_8821),
.B(n_1043),
.Y(n_9380)
);

OAI21xp5_ASAP7_75t_L g9381 ( 
.A1(n_8896),
.A2(n_162),
.B(n_163),
.Y(n_9381)
);

AOI21x1_ASAP7_75t_L g9382 ( 
.A1(n_8929),
.A2(n_162),
.B(n_163),
.Y(n_9382)
);

NOR2xp33_ASAP7_75t_L g9383 ( 
.A(n_8821),
.B(n_1045),
.Y(n_9383)
);

NAND2xp5_ASAP7_75t_SL g9384 ( 
.A(n_8934),
.B(n_8833),
.Y(n_9384)
);

BUFx12f_ASAP7_75t_L g9385 ( 
.A(n_9055),
.Y(n_9385)
);

BUFx6f_ASAP7_75t_L g9386 ( 
.A(n_9041),
.Y(n_9386)
);

NAND2xp5_ASAP7_75t_L g9387 ( 
.A(n_8909),
.B(n_1045),
.Y(n_9387)
);

NOR2xp33_ASAP7_75t_L g9388 ( 
.A(n_8697),
.B(n_8826),
.Y(n_9388)
);

NAND2xp33_ASAP7_75t_SL g9389 ( 
.A(n_8615),
.B(n_1046),
.Y(n_9389)
);

BUFx3_ASAP7_75t_L g9390 ( 
.A(n_9097),
.Y(n_9390)
);

INVx3_ASAP7_75t_SL g9391 ( 
.A(n_8570),
.Y(n_9391)
);

BUFx2_ASAP7_75t_L g9392 ( 
.A(n_8613),
.Y(n_9392)
);

NAND2xp5_ASAP7_75t_L g9393 ( 
.A(n_8583),
.B(n_1046),
.Y(n_9393)
);

NAND2xp5_ASAP7_75t_L g9394 ( 
.A(n_8558),
.B(n_1047),
.Y(n_9394)
);

NOR2xp67_ASAP7_75t_L g9395 ( 
.A(n_8733),
.B(n_164),
.Y(n_9395)
);

INVx1_ASAP7_75t_L g9396 ( 
.A(n_8762),
.Y(n_9396)
);

AOI21xp5_ASAP7_75t_L g9397 ( 
.A1(n_8962),
.A2(n_1048),
.B(n_1047),
.Y(n_9397)
);

AOI21xp5_ASAP7_75t_L g9398 ( 
.A1(n_8720),
.A2(n_1049),
.B(n_1048),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_SL g9399 ( 
.A(n_8789),
.B(n_1049),
.Y(n_9399)
);

INVx2_ASAP7_75t_L g9400 ( 
.A(n_8701),
.Y(n_9400)
);

NAND2xp5_ASAP7_75t_SL g9401 ( 
.A(n_8789),
.B(n_8804),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_8704),
.Y(n_9402)
);

AOI21xp5_ASAP7_75t_L g9403 ( 
.A1(n_8819),
.A2(n_1051),
.B(n_1050),
.Y(n_9403)
);

BUFx12f_ASAP7_75t_L g9404 ( 
.A(n_9104),
.Y(n_9404)
);

INVxp67_ASAP7_75t_L g9405 ( 
.A(n_8753),
.Y(n_9405)
);

AO22x1_ASAP7_75t_L g9406 ( 
.A1(n_8891),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_9406)
);

OA22x2_ASAP7_75t_L g9407 ( 
.A1(n_8627),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_9407)
);

INVx3_ASAP7_75t_L g9408 ( 
.A(n_8784),
.Y(n_9408)
);

AOI21xp5_ASAP7_75t_L g9409 ( 
.A1(n_8837),
.A2(n_1051),
.B(n_1050),
.Y(n_9409)
);

INVx1_ASAP7_75t_L g9410 ( 
.A(n_8764),
.Y(n_9410)
);

AOI21xp5_ASAP7_75t_L g9411 ( 
.A1(n_8904),
.A2(n_1053),
.B(n_1052),
.Y(n_9411)
);

AOI22xp5_ASAP7_75t_L g9412 ( 
.A1(n_8681),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_9412)
);

NAND2xp5_ASAP7_75t_SL g9413 ( 
.A(n_8804),
.B(n_1052),
.Y(n_9413)
);

AOI21xp5_ASAP7_75t_L g9414 ( 
.A1(n_8890),
.A2(n_1054),
.B(n_1053),
.Y(n_9414)
);

NAND2xp5_ASAP7_75t_SL g9415 ( 
.A(n_8872),
.B(n_1054),
.Y(n_9415)
);

AOI22xp33_ASAP7_75t_L g9416 ( 
.A1(n_8674),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_9416)
);

AO21x1_ASAP7_75t_L g9417 ( 
.A1(n_8983),
.A2(n_167),
.B(n_169),
.Y(n_9417)
);

BUFx6f_ASAP7_75t_L g9418 ( 
.A(n_9065),
.Y(n_9418)
);

O2A1O1Ixp33_ASAP7_75t_SL g9419 ( 
.A1(n_8815),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_9419)
);

O2A1O1Ixp33_ASAP7_75t_L g9420 ( 
.A1(n_8907),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_9420)
);

A2O1A1Ixp33_ASAP7_75t_L g9421 ( 
.A1(n_8617),
.A2(n_1056),
.B(n_1057),
.C(n_1055),
.Y(n_9421)
);

O2A1O1Ixp33_ASAP7_75t_SL g9422 ( 
.A1(n_8876),
.A2(n_173),
.B(n_170),
.C(n_172),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8768),
.Y(n_9423)
);

NAND2x1p5_ASAP7_75t_L g9424 ( 
.A(n_8544),
.B(n_1056),
.Y(n_9424)
);

INVx2_ASAP7_75t_L g9425 ( 
.A(n_8726),
.Y(n_9425)
);

AOI21xp5_ASAP7_75t_L g9426 ( 
.A1(n_8563),
.A2(n_1058),
.B(n_1057),
.Y(n_9426)
);

AOI21xp5_ASAP7_75t_L g9427 ( 
.A1(n_8568),
.A2(n_1060),
.B(n_1059),
.Y(n_9427)
);

AOI21xp5_ASAP7_75t_L g9428 ( 
.A1(n_8584),
.A2(n_1060),
.B(n_1059),
.Y(n_9428)
);

AO22x1_ASAP7_75t_L g9429 ( 
.A1(n_8891),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_9429)
);

AOI22xp33_ASAP7_75t_L g9430 ( 
.A1(n_9035),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_9430)
);

NAND2xp5_ASAP7_75t_SL g9431 ( 
.A(n_8872),
.B(n_1061),
.Y(n_9431)
);

OA22x2_ASAP7_75t_L g9432 ( 
.A1(n_8735),
.A2(n_177),
.B1(n_174),
.B2(n_175),
.Y(n_9432)
);

AOI21xp5_ASAP7_75t_L g9433 ( 
.A1(n_8589),
.A2(n_8596),
.B(n_8591),
.Y(n_9433)
);

NAND2xp5_ASAP7_75t_L g9434 ( 
.A(n_8597),
.B(n_1061),
.Y(n_9434)
);

NAND2xp5_ASAP7_75t_L g9435 ( 
.A(n_8598),
.B(n_1063),
.Y(n_9435)
);

NAND2xp5_ASAP7_75t_L g9436 ( 
.A(n_8604),
.B(n_1063),
.Y(n_9436)
);

INVx4_ASAP7_75t_L g9437 ( 
.A(n_9104),
.Y(n_9437)
);

INVx11_ASAP7_75t_L g9438 ( 
.A(n_8657),
.Y(n_9438)
);

OR2x2_ASAP7_75t_L g9439 ( 
.A(n_8774),
.B(n_1065),
.Y(n_9439)
);

AOI21x1_ASAP7_75t_L g9440 ( 
.A1(n_8695),
.A2(n_177),
.B(n_178),
.Y(n_9440)
);

O2A1O1Ixp5_ASAP7_75t_L g9441 ( 
.A1(n_8956),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_9441)
);

AOI21xp5_ASAP7_75t_L g9442 ( 
.A1(n_8610),
.A2(n_1066),
.B(n_1065),
.Y(n_9442)
);

A2O1A1Ixp33_ASAP7_75t_L g9443 ( 
.A1(n_8776),
.A2(n_8661),
.B(n_9022),
.C(n_8710),
.Y(n_9443)
);

NAND2xp5_ASAP7_75t_L g9444 ( 
.A(n_8623),
.B(n_1066),
.Y(n_9444)
);

OAI21xp33_ASAP7_75t_L g9445 ( 
.A1(n_8738),
.A2(n_179),
.B(n_180),
.Y(n_9445)
);

NOR2xp67_ASAP7_75t_L g9446 ( 
.A(n_8731),
.B(n_179),
.Y(n_9446)
);

AOI21xp33_ASAP7_75t_L g9447 ( 
.A1(n_8581),
.A2(n_180),
.B(n_181),
.Y(n_9447)
);

OAI21xp5_ASAP7_75t_L g9448 ( 
.A1(n_8541),
.A2(n_181),
.B(n_182),
.Y(n_9448)
);

BUFx3_ASAP7_75t_L g9449 ( 
.A(n_9080),
.Y(n_9449)
);

OAI21xp5_ASAP7_75t_L g9450 ( 
.A1(n_8678),
.A2(n_181),
.B(n_182),
.Y(n_9450)
);

INVx1_ASAP7_75t_L g9451 ( 
.A(n_8781),
.Y(n_9451)
);

O2A1O1Ixp33_ASAP7_75t_L g9452 ( 
.A1(n_8888),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_9452)
);

AOI22xp33_ASAP7_75t_L g9453 ( 
.A1(n_9068),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_9453)
);

AOI22xp33_ASAP7_75t_L g9454 ( 
.A1(n_9069),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_9454)
);

AOI21xp5_ASAP7_75t_L g9455 ( 
.A1(n_8631),
.A2(n_1068),
.B(n_1067),
.Y(n_9455)
);

OR2x2_ASAP7_75t_L g9456 ( 
.A(n_8783),
.B(n_1067),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_L g9457 ( 
.A(n_8632),
.B(n_1068),
.Y(n_9457)
);

NOR2xp33_ASAP7_75t_L g9458 ( 
.A(n_8684),
.B(n_1069),
.Y(n_9458)
);

NOR2xp67_ASAP7_75t_L g9459 ( 
.A(n_8752),
.B(n_185),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_8786),
.Y(n_9460)
);

NAND2xp5_ASAP7_75t_L g9461 ( 
.A(n_8634),
.B(n_1069),
.Y(n_9461)
);

HB1xp67_ASAP7_75t_L g9462 ( 
.A(n_8696),
.Y(n_9462)
);

AND2x2_ASAP7_75t_L g9463 ( 
.A(n_8725),
.B(n_1070),
.Y(n_9463)
);

AOI21xp5_ASAP7_75t_L g9464 ( 
.A1(n_8640),
.A2(n_1071),
.B(n_1070),
.Y(n_9464)
);

NOR2x1_ASAP7_75t_R g9465 ( 
.A(n_8807),
.B(n_186),
.Y(n_9465)
);

NAND2xp5_ASAP7_75t_L g9466 ( 
.A(n_8648),
.B(n_1071),
.Y(n_9466)
);

NAND2xp5_ASAP7_75t_L g9467 ( 
.A(n_8649),
.B(n_1072),
.Y(n_9467)
);

AOI21x1_ASAP7_75t_L g9468 ( 
.A1(n_8923),
.A2(n_186),
.B(n_187),
.Y(n_9468)
);

AOI21xp5_ASAP7_75t_L g9469 ( 
.A1(n_8653),
.A2(n_1074),
.B(n_1073),
.Y(n_9469)
);

INVx1_ASAP7_75t_L g9470 ( 
.A(n_8788),
.Y(n_9470)
);

INVx2_ASAP7_75t_L g9471 ( 
.A(n_8744),
.Y(n_9471)
);

A2O1A1Ixp33_ASAP7_75t_L g9472 ( 
.A1(n_8675),
.A2(n_1074),
.B(n_1075),
.C(n_1073),
.Y(n_9472)
);

NAND2xp5_ASAP7_75t_SL g9473 ( 
.A(n_8881),
.B(n_1075),
.Y(n_9473)
);

AND2x2_ASAP7_75t_L g9474 ( 
.A(n_8743),
.B(n_1076),
.Y(n_9474)
);

AOI21xp5_ASAP7_75t_L g9475 ( 
.A1(n_8925),
.A2(n_1077),
.B(n_1076),
.Y(n_9475)
);

NAND2xp5_ASAP7_75t_L g9476 ( 
.A(n_8595),
.B(n_1078),
.Y(n_9476)
);

NAND2xp5_ASAP7_75t_L g9477 ( 
.A(n_8749),
.B(n_1078),
.Y(n_9477)
);

O2A1O1Ixp33_ASAP7_75t_SL g9478 ( 
.A1(n_9000),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_9478)
);

INVx3_ASAP7_75t_L g9479 ( 
.A(n_8760),
.Y(n_9479)
);

AOI21xp5_ASAP7_75t_L g9480 ( 
.A1(n_8926),
.A2(n_1080),
.B(n_1079),
.Y(n_9480)
);

INVx2_ASAP7_75t_L g9481 ( 
.A(n_8867),
.Y(n_9481)
);

AOI21xp5_ASAP7_75t_L g9482 ( 
.A1(n_8864),
.A2(n_1080),
.B(n_1079),
.Y(n_9482)
);

OAI22xp5_ASAP7_75t_L g9483 ( 
.A1(n_9109),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_9483)
);

NAND2xp5_ASAP7_75t_L g9484 ( 
.A(n_8666),
.B(n_1081),
.Y(n_9484)
);

NOR2xp33_ASAP7_75t_L g9485 ( 
.A(n_8756),
.B(n_1081),
.Y(n_9485)
);

NAND2xp5_ASAP7_75t_SL g9486 ( 
.A(n_8881),
.B(n_1082),
.Y(n_9486)
);

AOI21xp5_ASAP7_75t_L g9487 ( 
.A1(n_8864),
.A2(n_1083),
.B(n_1082),
.Y(n_9487)
);

AOI21xp5_ASAP7_75t_L g9488 ( 
.A1(n_8814),
.A2(n_1084),
.B(n_1083),
.Y(n_9488)
);

AOI21xp5_ASAP7_75t_L g9489 ( 
.A1(n_9009),
.A2(n_1085),
.B(n_1084),
.Y(n_9489)
);

INVx4_ASAP7_75t_L g9490 ( 
.A(n_8811),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_8794),
.Y(n_9491)
);

NAND2xp5_ASAP7_75t_L g9492 ( 
.A(n_8732),
.B(n_1088),
.Y(n_9492)
);

AND2x4_ASAP7_75t_L g9493 ( 
.A(n_8621),
.B(n_1089),
.Y(n_9493)
);

BUFx6f_ASAP7_75t_L g9494 ( 
.A(n_9089),
.Y(n_9494)
);

NAND2xp5_ASAP7_75t_L g9495 ( 
.A(n_8739),
.B(n_1089),
.Y(n_9495)
);

O2A1O1Ixp33_ASAP7_75t_L g9496 ( 
.A1(n_8917),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_9496)
);

BUFx6f_ASAP7_75t_L g9497 ( 
.A(n_8748),
.Y(n_9497)
);

BUFx2_ASAP7_75t_L g9498 ( 
.A(n_8820),
.Y(n_9498)
);

INVx1_ASAP7_75t_L g9499 ( 
.A(n_8797),
.Y(n_9499)
);

AOI21xp5_ASAP7_75t_L g9500 ( 
.A1(n_9020),
.A2(n_1091),
.B(n_1090),
.Y(n_9500)
);

OAI22xp5_ASAP7_75t_L g9501 ( 
.A1(n_8594),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_9501)
);

BUFx6f_ASAP7_75t_L g9502 ( 
.A(n_8820),
.Y(n_9502)
);

AOI21xp5_ASAP7_75t_L g9503 ( 
.A1(n_8800),
.A2(n_1092),
.B(n_1090),
.Y(n_9503)
);

CKINVDCx20_ASAP7_75t_R g9504 ( 
.A(n_8742),
.Y(n_9504)
);

NOR2xp33_ASAP7_75t_L g9505 ( 
.A(n_8807),
.B(n_1093),
.Y(n_9505)
);

INVx2_ASAP7_75t_L g9506 ( 
.A(n_8861),
.Y(n_9506)
);

AOI21xp5_ASAP7_75t_L g9507 ( 
.A1(n_8817),
.A2(n_1094),
.B(n_1093),
.Y(n_9507)
);

OAI22xp5_ASAP7_75t_SL g9508 ( 
.A1(n_8668),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_9508)
);

NAND2xp5_ASAP7_75t_L g9509 ( 
.A(n_8740),
.B(n_1094),
.Y(n_9509)
);

AOI21xp5_ASAP7_75t_L g9510 ( 
.A1(n_8835),
.A2(n_1097),
.B(n_1096),
.Y(n_9510)
);

AOI22xp5_ASAP7_75t_L g9511 ( 
.A1(n_9028),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_9511)
);

AND2x2_ASAP7_75t_L g9512 ( 
.A(n_8831),
.B(n_1098),
.Y(n_9512)
);

NAND2xp5_ASAP7_75t_L g9513 ( 
.A(n_8816),
.B(n_1098),
.Y(n_9513)
);

INVx4_ASAP7_75t_L g9514 ( 
.A(n_8811),
.Y(n_9514)
);

NAND2xp5_ASAP7_75t_SL g9515 ( 
.A(n_8900),
.B(n_8910),
.Y(n_9515)
);

NOR2xp67_ASAP7_75t_SL g9516 ( 
.A(n_8910),
.B(n_193),
.Y(n_9516)
);

NAND2xp5_ASAP7_75t_L g9517 ( 
.A(n_8832),
.B(n_1099),
.Y(n_9517)
);

AOI221xp5_ASAP7_75t_L g9518 ( 
.A1(n_8607),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_9518)
);

NOR2xp33_ASAP7_75t_SL g9519 ( 
.A(n_8792),
.B(n_194),
.Y(n_9519)
);

NAND2xp5_ASAP7_75t_L g9520 ( 
.A(n_8644),
.B(n_1100),
.Y(n_9520)
);

OAI22xp5_ASAP7_75t_L g9521 ( 
.A1(n_8737),
.A2(n_8689),
.B1(n_8671),
.B2(n_8850),
.Y(n_9521)
);

AND2x2_ASAP7_75t_L g9522 ( 
.A(n_9034),
.B(n_1100),
.Y(n_9522)
);

AOI22xp5_ASAP7_75t_L g9523 ( 
.A1(n_8846),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_9523)
);

NAND2xp5_ASAP7_75t_L g9524 ( 
.A(n_8652),
.B(n_1101),
.Y(n_9524)
);

AOI21xp5_ASAP7_75t_L g9525 ( 
.A1(n_8839),
.A2(n_1102),
.B(n_1101),
.Y(n_9525)
);

INVxp33_ASAP7_75t_SL g9526 ( 
.A(n_8566),
.Y(n_9526)
);

XOR2xp5_ASAP7_75t_L g9527 ( 
.A(n_8799),
.B(n_195),
.Y(n_9527)
);

INVx2_ASAP7_75t_L g9528 ( 
.A(n_8865),
.Y(n_9528)
);

AOI21xp5_ASAP7_75t_L g9529 ( 
.A1(n_8841),
.A2(n_1103),
.B(n_1102),
.Y(n_9529)
);

AOI21xp5_ASAP7_75t_L g9530 ( 
.A1(n_8845),
.A2(n_1105),
.B(n_1104),
.Y(n_9530)
);

NAND2xp5_ASAP7_75t_L g9531 ( 
.A(n_8955),
.B(n_1104),
.Y(n_9531)
);

BUFx6f_ASAP7_75t_L g9532 ( 
.A(n_8770),
.Y(n_9532)
);

NOR2xp33_ASAP7_75t_L g9533 ( 
.A(n_8812),
.B(n_1105),
.Y(n_9533)
);

NAND2xp5_ASAP7_75t_L g9534 ( 
.A(n_8957),
.B(n_1106),
.Y(n_9534)
);

AND2x2_ASAP7_75t_L g9535 ( 
.A(n_9081),
.B(n_1106),
.Y(n_9535)
);

NAND2xp5_ASAP7_75t_L g9536 ( 
.A(n_8965),
.B(n_1107),
.Y(n_9536)
);

AOI21xp5_ASAP7_75t_L g9537 ( 
.A1(n_8859),
.A2(n_1108),
.B(n_1107),
.Y(n_9537)
);

OAI21x1_ASAP7_75t_L g9538 ( 
.A1(n_8869),
.A2(n_196),
.B(n_197),
.Y(n_9538)
);

BUFx2_ASAP7_75t_L g9539 ( 
.A(n_8862),
.Y(n_9539)
);

BUFx4f_ASAP7_75t_L g9540 ( 
.A(n_8933),
.Y(n_9540)
);

AOI21xp33_ASAP7_75t_L g9541 ( 
.A1(n_8741),
.A2(n_197),
.B(n_198),
.Y(n_9541)
);

NOR2xp33_ASAP7_75t_L g9542 ( 
.A(n_8785),
.B(n_1108),
.Y(n_9542)
);

NAND2xp5_ASAP7_75t_L g9543 ( 
.A(n_8967),
.B(n_1109),
.Y(n_9543)
);

AOI21xp5_ASAP7_75t_L g9544 ( 
.A1(n_8870),
.A2(n_1111),
.B(n_1110),
.Y(n_9544)
);

AOI21xp5_ASAP7_75t_L g9545 ( 
.A1(n_8877),
.A2(n_1112),
.B(n_1111),
.Y(n_9545)
);

O2A1O1Ixp5_ASAP7_75t_L g9546 ( 
.A1(n_8707),
.A2(n_8718),
.B(n_8979),
.C(n_8974),
.Y(n_9546)
);

NOR3xp33_ASAP7_75t_L g9547 ( 
.A(n_8572),
.B(n_198),
.C(n_199),
.Y(n_9547)
);

AOI22x1_ASAP7_75t_L g9548 ( 
.A1(n_8801),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_9548)
);

INVx3_ASAP7_75t_L g9549 ( 
.A(n_8683),
.Y(n_9549)
);

AOI21xp5_ASAP7_75t_L g9550 ( 
.A1(n_8879),
.A2(n_1113),
.B(n_1112),
.Y(n_9550)
);

A2O1A1Ixp33_ASAP7_75t_L g9551 ( 
.A1(n_8836),
.A2(n_1114),
.B(n_1115),
.C(n_1113),
.Y(n_9551)
);

HB1xp67_ASAP7_75t_L g9552 ( 
.A(n_8900),
.Y(n_9552)
);

AOI21xp5_ASAP7_75t_L g9553 ( 
.A1(n_8988),
.A2(n_1115),
.B(n_1114),
.Y(n_9553)
);

NAND2xp5_ASAP7_75t_L g9554 ( 
.A(n_8996),
.B(n_1116),
.Y(n_9554)
);

NAND3xp33_ASAP7_75t_L g9555 ( 
.A(n_8920),
.B(n_200),
.C(n_201),
.Y(n_9555)
);

NAND2xp5_ASAP7_75t_L g9556 ( 
.A(n_8791),
.B(n_1116),
.Y(n_9556)
);

NAND2x1p5_ASAP7_75t_L g9557 ( 
.A(n_8693),
.B(n_8813),
.Y(n_9557)
);

NAND2xp5_ASAP7_75t_L g9558 ( 
.A(n_8745),
.B(n_1117),
.Y(n_9558)
);

NAND2xp5_ASAP7_75t_L g9559 ( 
.A(n_8779),
.B(n_1117),
.Y(n_9559)
);

AOI21xp5_ASAP7_75t_L g9560 ( 
.A1(n_8950),
.A2(n_1119),
.B(n_1118),
.Y(n_9560)
);

NOR3xp33_ASAP7_75t_L g9561 ( 
.A(n_8822),
.B(n_200),
.C(n_201),
.Y(n_9561)
);

NAND2xp5_ASAP7_75t_SL g9562 ( 
.A(n_8611),
.B(n_1118),
.Y(n_9562)
);

NAND2xp5_ASAP7_75t_L g9563 ( 
.A(n_8949),
.B(n_1120),
.Y(n_9563)
);

AND2x2_ASAP7_75t_L g9564 ( 
.A(n_9083),
.B(n_1120),
.Y(n_9564)
);

HB1xp67_ASAP7_75t_L g9565 ( 
.A(n_8750),
.Y(n_9565)
);

AOI21xp5_ASAP7_75t_L g9566 ( 
.A1(n_9027),
.A2(n_1122),
.B(n_1121),
.Y(n_9566)
);

AOI21xp5_ASAP7_75t_L g9567 ( 
.A1(n_8778),
.A2(n_1122),
.B(n_1121),
.Y(n_9567)
);

CKINVDCx20_ASAP7_75t_R g9568 ( 
.A(n_8932),
.Y(n_9568)
);

BUFx4f_ASAP7_75t_L g9569 ( 
.A(n_8646),
.Y(n_9569)
);

NOR2xp33_ASAP7_75t_L g9570 ( 
.A(n_8580),
.B(n_8567),
.Y(n_9570)
);

O2A1O1Ixp33_ASAP7_75t_L g9571 ( 
.A1(n_9025),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_9571)
);

O2A1O1Ixp33_ASAP7_75t_SL g9572 ( 
.A1(n_8642),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_9572)
);

NAND2xp5_ASAP7_75t_L g9573 ( 
.A(n_8976),
.B(n_1123),
.Y(n_9573)
);

AND2x2_ASAP7_75t_L g9574 ( 
.A(n_9105),
.B(n_1123),
.Y(n_9574)
);

NOR2x1p5_ASAP7_75t_SL g9575 ( 
.A(n_9067),
.B(n_1124),
.Y(n_9575)
);

NOR2xp33_ASAP7_75t_L g9576 ( 
.A(n_8787),
.B(n_1124),
.Y(n_9576)
);

HB1xp67_ASAP7_75t_L g9577 ( 
.A(n_8714),
.Y(n_9577)
);

AND2x2_ASAP7_75t_L g9578 ( 
.A(n_8908),
.B(n_1125),
.Y(n_9578)
);

NAND2x1p5_ASAP7_75t_L g9579 ( 
.A(n_8571),
.B(n_1125),
.Y(n_9579)
);

NAND2x1_ASAP7_75t_L g9580 ( 
.A(n_8997),
.B(n_1126),
.Y(n_9580)
);

NOR2xp33_ASAP7_75t_L g9581 ( 
.A(n_8532),
.B(n_1126),
.Y(n_9581)
);

O2A1O1Ixp5_ASAP7_75t_L g9582 ( 
.A1(n_8857),
.A2(n_205),
.B(n_202),
.C(n_204),
.Y(n_9582)
);

AOI21xp5_ASAP7_75t_L g9583 ( 
.A1(n_8885),
.A2(n_1128),
.B(n_1127),
.Y(n_9583)
);

O2A1O1Ixp5_ASAP7_75t_L g9584 ( 
.A1(n_8823),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_9584)
);

AO32x1_ASAP7_75t_L g9585 ( 
.A1(n_9062),
.A2(n_207),
.A3(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_9585)
);

NAND2x1p5_ASAP7_75t_L g9586 ( 
.A(n_8609),
.B(n_1127),
.Y(n_9586)
);

O2A1O1Ixp33_ASAP7_75t_L g9587 ( 
.A1(n_9054),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_9587)
);

OAI21xp5_ASAP7_75t_L g9588 ( 
.A1(n_8916),
.A2(n_207),
.B(n_208),
.Y(n_9588)
);

AOI21xp5_ASAP7_75t_L g9589 ( 
.A1(n_8943),
.A2(n_1130),
.B(n_1129),
.Y(n_9589)
);

INVx2_ASAP7_75t_L g9590 ( 
.A(n_8842),
.Y(n_9590)
);

HB1xp67_ASAP7_75t_L g9591 ( 
.A(n_8734),
.Y(n_9591)
);

A2O1A1Ixp33_ASAP7_75t_L g9592 ( 
.A1(n_8847),
.A2(n_1131),
.B(n_1132),
.C(n_1129),
.Y(n_9592)
);

INVx4_ASAP7_75t_L g9593 ( 
.A(n_8706),
.Y(n_9593)
);

AND2x2_ASAP7_75t_L g9594 ( 
.A(n_8924),
.B(n_1131),
.Y(n_9594)
);

INVx1_ASAP7_75t_L g9595 ( 
.A(n_8602),
.Y(n_9595)
);

INVx2_ASAP7_75t_L g9596 ( 
.A(n_8717),
.Y(n_9596)
);

O2A1O1Ixp33_ASAP7_75t_L g9597 ( 
.A1(n_8802),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_9597)
);

AND2x6_ASAP7_75t_L g9598 ( 
.A(n_8964),
.B(n_1132),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_8618),
.Y(n_9599)
);

AOI21xp5_ASAP7_75t_L g9600 ( 
.A1(n_8716),
.A2(n_1134),
.B(n_1133),
.Y(n_9600)
);

NAND2xp5_ASAP7_75t_L g9601 ( 
.A(n_8937),
.B(n_1134),
.Y(n_9601)
);

OAI21xp5_ASAP7_75t_L g9602 ( 
.A1(n_8897),
.A2(n_209),
.B(n_210),
.Y(n_9602)
);

INVx1_ASAP7_75t_L g9603 ( 
.A(n_8891),
.Y(n_9603)
);

NAND2xp5_ASAP7_75t_L g9604 ( 
.A(n_8765),
.B(n_1135),
.Y(n_9604)
);

INVx1_ASAP7_75t_SL g9605 ( 
.A(n_8761),
.Y(n_9605)
);

OR2x2_ASAP7_75t_L g9606 ( 
.A(n_8767),
.B(n_1135),
.Y(n_9606)
);

AND2x2_ASAP7_75t_L g9607 ( 
.A(n_8856),
.B(n_1136),
.Y(n_9607)
);

AOI21xp5_ASAP7_75t_L g9608 ( 
.A1(n_8772),
.A2(n_1137),
.B(n_1136),
.Y(n_9608)
);

BUFx8_ASAP7_75t_L g9609 ( 
.A(n_8868),
.Y(n_9609)
);

AOI21xp5_ASAP7_75t_L g9610 ( 
.A1(n_8830),
.A2(n_1138),
.B(n_1137),
.Y(n_9610)
);

INVx1_ASAP7_75t_SL g9611 ( 
.A(n_8763),
.Y(n_9611)
);

NOR2xp33_ASAP7_75t_L g9612 ( 
.A(n_8834),
.B(n_1138),
.Y(n_9612)
);

OAI22xp5_ASAP7_75t_L g9613 ( 
.A1(n_8673),
.A2(n_212),
.B1(n_209),
.B2(n_211),
.Y(n_9613)
);

CKINVDCx10_ASAP7_75t_R g9614 ( 
.A(n_8646),
.Y(n_9614)
);

INVxp67_ASAP7_75t_L g9615 ( 
.A(n_8537),
.Y(n_9615)
);

NOR2xp33_ASAP7_75t_L g9616 ( 
.A(n_8805),
.B(n_1139),
.Y(n_9616)
);

AOI21xp5_ASAP7_75t_L g9617 ( 
.A1(n_8843),
.A2(n_8849),
.B(n_8893),
.Y(n_9617)
);

OAI21x1_ASAP7_75t_L g9618 ( 
.A1(n_9074),
.A2(n_211),
.B(n_212),
.Y(n_9618)
);

AOI21xp5_ASAP7_75t_L g9619 ( 
.A1(n_8893),
.A2(n_1140),
.B(n_1139),
.Y(n_9619)
);

NAND2xp5_ASAP7_75t_L g9620 ( 
.A(n_8664),
.B(n_1140),
.Y(n_9620)
);

A2O1A1Ixp33_ASAP7_75t_L g9621 ( 
.A1(n_8773),
.A2(n_1142),
.B(n_1143),
.C(n_1141),
.Y(n_9621)
);

AOI21xp5_ASAP7_75t_L g9622 ( 
.A1(n_8808),
.A2(n_8790),
.B(n_8782),
.Y(n_9622)
);

NAND2xp5_ASAP7_75t_L g9623 ( 
.A(n_8619),
.B(n_1142),
.Y(n_9623)
);

OR2x6_ASAP7_75t_L g9624 ( 
.A(n_8698),
.B(n_1144),
.Y(n_9624)
);

NAND3xp33_ASAP7_75t_L g9625 ( 
.A(n_8810),
.B(n_213),
.C(n_214),
.Y(n_9625)
);

AND2x6_ASAP7_75t_L g9626 ( 
.A(n_8997),
.B(n_1144),
.Y(n_9626)
);

INVx1_ASAP7_75t_L g9627 ( 
.A(n_8730),
.Y(n_9627)
);

NAND2xp5_ASAP7_75t_L g9628 ( 
.A(n_8655),
.B(n_1145),
.Y(n_9628)
);

AOI21xp5_ASAP7_75t_L g9629 ( 
.A1(n_9108),
.A2(n_1146),
.B(n_1145),
.Y(n_9629)
);

AND2x2_ASAP7_75t_SL g9630 ( 
.A(n_9088),
.B(n_1147),
.Y(n_9630)
);

INVx1_ASAP7_75t_L g9631 ( 
.A(n_8754),
.Y(n_9631)
);

BUFx6f_ASAP7_75t_L g9632 ( 
.A(n_8531),
.Y(n_9632)
);

OAI21xp5_ASAP7_75t_L g9633 ( 
.A1(n_8573),
.A2(n_213),
.B(n_214),
.Y(n_9633)
);

OAI22xp33_ASAP7_75t_L g9634 ( 
.A1(n_8698),
.A2(n_1148),
.B1(n_1149),
.B2(n_1147),
.Y(n_9634)
);

AOI21xp5_ASAP7_75t_L g9635 ( 
.A1(n_9108),
.A2(n_1149),
.B(n_1148),
.Y(n_9635)
);

AND2x2_ASAP7_75t_L g9636 ( 
.A(n_8651),
.B(n_1150),
.Y(n_9636)
);

NAND2xp5_ASAP7_75t_L g9637 ( 
.A(n_9038),
.B(n_1150),
.Y(n_9637)
);

AND2x4_ASAP7_75t_L g9638 ( 
.A(n_8700),
.B(n_1151),
.Y(n_9638)
);

OR2x2_ASAP7_75t_L g9639 ( 
.A(n_8635),
.B(n_1152),
.Y(n_9639)
);

NOR2xp33_ASAP7_75t_L g9640 ( 
.A(n_8535),
.B(n_1152),
.Y(n_9640)
);

NOR2xp33_ASAP7_75t_L g9641 ( 
.A(n_8746),
.B(n_8682),
.Y(n_9641)
);

OAI21xp5_ASAP7_75t_L g9642 ( 
.A1(n_8569),
.A2(n_214),
.B(n_215),
.Y(n_9642)
);

A2O1A1Ixp33_ASAP7_75t_L g9643 ( 
.A1(n_8723),
.A2(n_1154),
.B(n_1155),
.C(n_1153),
.Y(n_9643)
);

AND2x2_ASAP7_75t_L g9644 ( 
.A(n_8766),
.B(n_1153),
.Y(n_9644)
);

NOR2xp33_ASAP7_75t_L g9645 ( 
.A(n_8709),
.B(n_1154),
.Y(n_9645)
);

AOI22xp33_ASAP7_75t_L g9646 ( 
.A1(n_9049),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_9646)
);

INVx6_ASAP7_75t_L g9647 ( 
.A(n_9091),
.Y(n_9647)
);

AO21x1_ASAP7_75t_L g9648 ( 
.A1(n_8662),
.A2(n_215),
.B(n_216),
.Y(n_9648)
);

NAND2xp5_ASAP7_75t_L g9649 ( 
.A(n_8700),
.B(n_1155),
.Y(n_9649)
);

NAND2xp5_ASAP7_75t_L g9650 ( 
.A(n_8622),
.B(n_8722),
.Y(n_9650)
);

AOI22xp5_ASAP7_75t_L g9651 ( 
.A1(n_8722),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_9651)
);

AOI21x1_ASAP7_75t_L g9652 ( 
.A1(n_8928),
.A2(n_217),
.B(n_218),
.Y(n_9652)
);

INVx3_ASAP7_75t_L g9653 ( 
.A(n_8643),
.Y(n_9653)
);

O2A1O1Ixp5_ASAP7_75t_L g9654 ( 
.A1(n_9078),
.A2(n_9110),
.B(n_8628),
.C(n_220),
.Y(n_9654)
);

AOI21xp5_ASAP7_75t_L g9655 ( 
.A1(n_8553),
.A2(n_1157),
.B(n_1156),
.Y(n_9655)
);

NAND2xp5_ASAP7_75t_L g9656 ( 
.A(n_8539),
.B(n_1156),
.Y(n_9656)
);

AOI21xp5_ASAP7_75t_L g9657 ( 
.A1(n_8553),
.A2(n_1159),
.B(n_1158),
.Y(n_9657)
);

OAI21xp5_ASAP7_75t_L g9658 ( 
.A1(n_8534),
.A2(n_218),
.B(n_219),
.Y(n_9658)
);

AOI21xp5_ASAP7_75t_L g9659 ( 
.A1(n_8553),
.A2(n_1159),
.B(n_1158),
.Y(n_9659)
);

O2A1O1Ixp33_ASAP7_75t_L g9660 ( 
.A1(n_8659),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_9660)
);

BUFx6f_ASAP7_75t_L g9661 ( 
.A(n_8575),
.Y(n_9661)
);

NAND2xp5_ASAP7_75t_L g9662 ( 
.A(n_8539),
.B(n_1160),
.Y(n_9662)
);

AOI21xp5_ASAP7_75t_L g9663 ( 
.A1(n_8553),
.A2(n_1161),
.B(n_1160),
.Y(n_9663)
);

AOI21xp5_ASAP7_75t_L g9664 ( 
.A1(n_8553),
.A2(n_1162),
.B(n_1161),
.Y(n_9664)
);

NAND2xp5_ASAP7_75t_SL g9665 ( 
.A(n_8539),
.B(n_1162),
.Y(n_9665)
);

AO21x1_ASAP7_75t_L g9666 ( 
.A1(n_8660),
.A2(n_220),
.B(n_221),
.Y(n_9666)
);

BUFx6f_ASAP7_75t_L g9667 ( 
.A(n_8575),
.Y(n_9667)
);

INVx1_ASAP7_75t_SL g9668 ( 
.A(n_8565),
.Y(n_9668)
);

NOR2xp33_ASAP7_75t_L g9669 ( 
.A(n_8539),
.B(n_1163),
.Y(n_9669)
);

AOI22xp33_ASAP7_75t_L g9670 ( 
.A1(n_9070),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_9670)
);

AOI21xp5_ASAP7_75t_L g9671 ( 
.A1(n_8553),
.A2(n_1165),
.B(n_1164),
.Y(n_9671)
);

NAND2xp5_ASAP7_75t_L g9672 ( 
.A(n_8539),
.B(n_1164),
.Y(n_9672)
);

AOI21xp5_ASAP7_75t_L g9673 ( 
.A1(n_8553),
.A2(n_1166),
.B(n_1165),
.Y(n_9673)
);

NOR2xp67_ASAP7_75t_L g9674 ( 
.A(n_9073),
.B(n_222),
.Y(n_9674)
);

A2O1A1Ixp33_ASAP7_75t_L g9675 ( 
.A1(n_8582),
.A2(n_1167),
.B(n_1168),
.C(n_1166),
.Y(n_9675)
);

INVx2_ASAP7_75t_L g9676 ( 
.A(n_8548),
.Y(n_9676)
);

AOI21xp5_ASAP7_75t_L g9677 ( 
.A1(n_8553),
.A2(n_1169),
.B(n_1168),
.Y(n_9677)
);

CKINVDCx8_ASAP7_75t_R g9678 ( 
.A(n_8894),
.Y(n_9678)
);

OAI22xp5_ASAP7_75t_L g9679 ( 
.A1(n_8729),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_9679)
);

AOI21xp5_ASAP7_75t_L g9680 ( 
.A1(n_8553),
.A2(n_1171),
.B(n_1170),
.Y(n_9680)
);

AND2x2_ASAP7_75t_L g9681 ( 
.A(n_8625),
.B(n_1170),
.Y(n_9681)
);

NAND3xp33_ASAP7_75t_SL g9682 ( 
.A(n_8729),
.B(n_223),
.C(n_224),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_8914),
.Y(n_9683)
);

A2O1A1Ixp33_ASAP7_75t_L g9684 ( 
.A1(n_8582),
.A2(n_1172),
.B(n_1173),
.C(n_1171),
.Y(n_9684)
);

AOI21xp5_ASAP7_75t_L g9685 ( 
.A1(n_8553),
.A2(n_1173),
.B(n_1172),
.Y(n_9685)
);

AOI22xp33_ASAP7_75t_L g9686 ( 
.A1(n_9070),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_9686)
);

OR2x6_ASAP7_75t_SL g9687 ( 
.A(n_9026),
.B(n_225),
.Y(n_9687)
);

INVx1_ASAP7_75t_L g9688 ( 
.A(n_8914),
.Y(n_9688)
);

NAND2xp5_ASAP7_75t_L g9689 ( 
.A(n_8539),
.B(n_1174),
.Y(n_9689)
);

INVx11_ASAP7_75t_L g9690 ( 
.A(n_9066),
.Y(n_9690)
);

OAI21xp5_ASAP7_75t_L g9691 ( 
.A1(n_8534),
.A2(n_225),
.B(n_226),
.Y(n_9691)
);

NOR3xp33_ASAP7_75t_L g9692 ( 
.A(n_8895),
.B(n_227),
.C(n_228),
.Y(n_9692)
);

AOI21xp5_ASAP7_75t_L g9693 ( 
.A1(n_8553),
.A2(n_1175),
.B(n_1174),
.Y(n_9693)
);

BUFx4f_ASAP7_75t_L g9694 ( 
.A(n_9047),
.Y(n_9694)
);

NAND2xp5_ASAP7_75t_L g9695 ( 
.A(n_8539),
.B(n_1175),
.Y(n_9695)
);

AOI21xp5_ASAP7_75t_L g9696 ( 
.A1(n_8553),
.A2(n_1177),
.B(n_1176),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_8914),
.Y(n_9697)
);

AOI21xp5_ASAP7_75t_L g9698 ( 
.A1(n_8553),
.A2(n_1177),
.B(n_1176),
.Y(n_9698)
);

NOR3xp33_ASAP7_75t_L g9699 ( 
.A(n_8895),
.B(n_227),
.C(n_229),
.Y(n_9699)
);

NAND2xp5_ASAP7_75t_SL g9700 ( 
.A(n_8539),
.B(n_1178),
.Y(n_9700)
);

A2O1A1Ixp33_ASAP7_75t_L g9701 ( 
.A1(n_8582),
.A2(n_1179),
.B(n_1180),
.C(n_1178),
.Y(n_9701)
);

AND2x2_ASAP7_75t_L g9702 ( 
.A(n_8625),
.B(n_1180),
.Y(n_9702)
);

INVx2_ASAP7_75t_SL g9703 ( 
.A(n_9073),
.Y(n_9703)
);

INVx4_ASAP7_75t_L g9704 ( 
.A(n_9073),
.Y(n_9704)
);

AOI21x1_ASAP7_75t_L g9705 ( 
.A1(n_8553),
.A2(n_229),
.B(n_230),
.Y(n_9705)
);

INVx1_ASAP7_75t_SL g9706 ( 
.A(n_8565),
.Y(n_9706)
);

NAND2xp5_ASAP7_75t_L g9707 ( 
.A(n_8539),
.B(n_1181),
.Y(n_9707)
);

NAND3xp33_ASAP7_75t_SL g9708 ( 
.A(n_8729),
.B(n_229),
.C(n_230),
.Y(n_9708)
);

AOI21xp5_ASAP7_75t_L g9709 ( 
.A1(n_8553),
.A2(n_1182),
.B(n_1181),
.Y(n_9709)
);

INVx2_ASAP7_75t_L g9710 ( 
.A(n_8548),
.Y(n_9710)
);

NAND2xp5_ASAP7_75t_L g9711 ( 
.A(n_8539),
.B(n_1183),
.Y(n_9711)
);

AND2x4_ASAP7_75t_L g9712 ( 
.A(n_9073),
.B(n_1183),
.Y(n_9712)
);

OAI21xp5_ASAP7_75t_L g9713 ( 
.A1(n_8534),
.A2(n_230),
.B(n_231),
.Y(n_9713)
);

NAND2xp5_ASAP7_75t_L g9714 ( 
.A(n_8539),
.B(n_1184),
.Y(n_9714)
);

AOI22xp5_ASAP7_75t_L g9715 ( 
.A1(n_8729),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_9715)
);

AOI21xp5_ASAP7_75t_L g9716 ( 
.A1(n_8553),
.A2(n_1185),
.B(n_1184),
.Y(n_9716)
);

NAND2xp5_ASAP7_75t_L g9717 ( 
.A(n_8539),
.B(n_1186),
.Y(n_9717)
);

NOR2xp33_ASAP7_75t_L g9718 ( 
.A(n_8539),
.B(n_1186),
.Y(n_9718)
);

INVx1_ASAP7_75t_L g9719 ( 
.A(n_8914),
.Y(n_9719)
);

NAND2xp5_ASAP7_75t_L g9720 ( 
.A(n_8539),
.B(n_1188),
.Y(n_9720)
);

NAND2xp5_ASAP7_75t_L g9721 ( 
.A(n_8539),
.B(n_1188),
.Y(n_9721)
);

NAND2xp5_ASAP7_75t_SL g9722 ( 
.A(n_8539),
.B(n_1189),
.Y(n_9722)
);

NAND2xp5_ASAP7_75t_L g9723 ( 
.A(n_8539),
.B(n_1189),
.Y(n_9723)
);

AOI21xp5_ASAP7_75t_L g9724 ( 
.A1(n_8553),
.A2(n_1191),
.B(n_1190),
.Y(n_9724)
);

CKINVDCx5p33_ASAP7_75t_R g9725 ( 
.A(n_8577),
.Y(n_9725)
);

OAI21xp5_ASAP7_75t_L g9726 ( 
.A1(n_8534),
.A2(n_232),
.B(n_233),
.Y(n_9726)
);

INVx1_ASAP7_75t_L g9727 ( 
.A(n_8914),
.Y(n_9727)
);

NAND2xp5_ASAP7_75t_SL g9728 ( 
.A(n_8539),
.B(n_1190),
.Y(n_9728)
);

OAI21xp5_ASAP7_75t_L g9729 ( 
.A1(n_8534),
.A2(n_232),
.B(n_234),
.Y(n_9729)
);

OR2x2_ASAP7_75t_L g9730 ( 
.A(n_8625),
.B(n_1191),
.Y(n_9730)
);

AOI21xp5_ASAP7_75t_L g9731 ( 
.A1(n_8553),
.A2(n_1193),
.B(n_1192),
.Y(n_9731)
);

AOI21xp5_ASAP7_75t_L g9732 ( 
.A1(n_8553),
.A2(n_1193),
.B(n_1192),
.Y(n_9732)
);

NAND2xp5_ASAP7_75t_L g9733 ( 
.A(n_8539),
.B(n_1194),
.Y(n_9733)
);

CKINVDCx5p33_ASAP7_75t_R g9734 ( 
.A(n_8577),
.Y(n_9734)
);

AND2x2_ASAP7_75t_L g9735 ( 
.A(n_8625),
.B(n_1194),
.Y(n_9735)
);

NAND2xp5_ASAP7_75t_SL g9736 ( 
.A(n_8539),
.B(n_1195),
.Y(n_9736)
);

AOI33xp33_ASAP7_75t_L g9737 ( 
.A1(n_8572),
.A2(n_236),
.A3(n_238),
.B1(n_234),
.B2(n_235),
.B3(n_237),
.Y(n_9737)
);

AOI21xp5_ASAP7_75t_L g9738 ( 
.A1(n_8553),
.A2(n_1197),
.B(n_1196),
.Y(n_9738)
);

AND2x4_ASAP7_75t_L g9739 ( 
.A(n_9073),
.B(n_1196),
.Y(n_9739)
);

AOI21xp5_ASAP7_75t_L g9740 ( 
.A1(n_8553),
.A2(n_1200),
.B(n_1199),
.Y(n_9740)
);

AND2x4_ASAP7_75t_L g9741 ( 
.A(n_9073),
.B(n_1199),
.Y(n_9741)
);

AOI21xp5_ASAP7_75t_L g9742 ( 
.A1(n_8553),
.A2(n_1201),
.B(n_1200),
.Y(n_9742)
);

O2A1O1Ixp33_ASAP7_75t_L g9743 ( 
.A1(n_8659),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_9743)
);

OAI22xp5_ASAP7_75t_L g9744 ( 
.A1(n_8729),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_9744)
);

NAND2xp5_ASAP7_75t_L g9745 ( 
.A(n_8539),
.B(n_1201),
.Y(n_9745)
);

OAI22xp5_ASAP7_75t_L g9746 ( 
.A1(n_8729),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_9746)
);

INVx4_ASAP7_75t_L g9747 ( 
.A(n_9073),
.Y(n_9747)
);

INVx2_ASAP7_75t_L g9748 ( 
.A(n_8548),
.Y(n_9748)
);

AOI21xp5_ASAP7_75t_L g9749 ( 
.A1(n_8553),
.A2(n_1203),
.B(n_1202),
.Y(n_9749)
);

NAND2xp5_ASAP7_75t_L g9750 ( 
.A(n_8539),
.B(n_1202),
.Y(n_9750)
);

INVx2_ASAP7_75t_L g9751 ( 
.A(n_8548),
.Y(n_9751)
);

AOI21xp5_ASAP7_75t_L g9752 ( 
.A1(n_8553),
.A2(n_1204),
.B(n_1203),
.Y(n_9752)
);

NAND2xp5_ASAP7_75t_L g9753 ( 
.A(n_8539),
.B(n_1204),
.Y(n_9753)
);

NAND3xp33_ASAP7_75t_SL g9754 ( 
.A(n_8729),
.B(n_238),
.C(n_239),
.Y(n_9754)
);

INVx1_ASAP7_75t_L g9755 ( 
.A(n_8914),
.Y(n_9755)
);

O2A1O1Ixp33_ASAP7_75t_L g9756 ( 
.A1(n_8659),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_9756)
);

NAND2xp5_ASAP7_75t_L g9757 ( 
.A(n_8539),
.B(n_1205),
.Y(n_9757)
);

INVx1_ASAP7_75t_L g9758 ( 
.A(n_8914),
.Y(n_9758)
);

NAND2xp5_ASAP7_75t_L g9759 ( 
.A(n_8539),
.B(n_1205),
.Y(n_9759)
);

A2O1A1Ixp33_ASAP7_75t_L g9760 ( 
.A1(n_8582),
.A2(n_1207),
.B(n_1208),
.C(n_1206),
.Y(n_9760)
);

NOR2xp33_ASAP7_75t_SL g9761 ( 
.A(n_8577),
.B(n_241),
.Y(n_9761)
);

OAI22xp5_ASAP7_75t_L g9762 ( 
.A1(n_8729),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_9762)
);

NAND2xp5_ASAP7_75t_L g9763 ( 
.A(n_8539),
.B(n_1206),
.Y(n_9763)
);

INVx1_ASAP7_75t_L g9764 ( 
.A(n_8914),
.Y(n_9764)
);

BUFx6f_ASAP7_75t_L g9765 ( 
.A(n_8575),
.Y(n_9765)
);

INVx1_ASAP7_75t_L g9766 ( 
.A(n_8914),
.Y(n_9766)
);

NAND2xp5_ASAP7_75t_L g9767 ( 
.A(n_8539),
.B(n_1207),
.Y(n_9767)
);

OAI21xp5_ASAP7_75t_L g9768 ( 
.A1(n_8534),
.A2(n_242),
.B(n_243),
.Y(n_9768)
);

A2O1A1Ixp33_ASAP7_75t_L g9769 ( 
.A1(n_8582),
.A2(n_1210),
.B(n_1211),
.C(n_1209),
.Y(n_9769)
);

AOI21xp5_ASAP7_75t_L g9770 ( 
.A1(n_8553),
.A2(n_1212),
.B(n_1211),
.Y(n_9770)
);

INVx1_ASAP7_75t_L g9771 ( 
.A(n_8914),
.Y(n_9771)
);

NOR3xp33_ASAP7_75t_L g9772 ( 
.A(n_8895),
.B(n_242),
.C(n_243),
.Y(n_9772)
);

NAND2xp5_ASAP7_75t_L g9773 ( 
.A(n_8539),
.B(n_1213),
.Y(n_9773)
);

A2O1A1Ixp33_ASAP7_75t_L g9774 ( 
.A1(n_8582),
.A2(n_1214),
.B(n_1215),
.C(n_1213),
.Y(n_9774)
);

AOI21xp5_ASAP7_75t_L g9775 ( 
.A1(n_8553),
.A2(n_1216),
.B(n_1214),
.Y(n_9775)
);

NAND2xp5_ASAP7_75t_L g9776 ( 
.A(n_9147),
.B(n_1216),
.Y(n_9776)
);

AND2x2_ASAP7_75t_L g9777 ( 
.A(n_9167),
.B(n_1217),
.Y(n_9777)
);

AOI21x1_ASAP7_75t_L g9778 ( 
.A1(n_9705),
.A2(n_244),
.B(n_245),
.Y(n_9778)
);

AOI21xp5_ASAP7_75t_L g9779 ( 
.A1(n_9123),
.A2(n_244),
.B(n_245),
.Y(n_9779)
);

A2O1A1Ixp33_ASAP7_75t_L g9780 ( 
.A1(n_9261),
.A2(n_1218),
.B(n_1219),
.C(n_1217),
.Y(n_9780)
);

OAI21x1_ASAP7_75t_SL g9781 ( 
.A1(n_9162),
.A2(n_244),
.B(n_246),
.Y(n_9781)
);

OAI21x1_ASAP7_75t_L g9782 ( 
.A1(n_9121),
.A2(n_247),
.B(n_248),
.Y(n_9782)
);

BUFx2_ASAP7_75t_L g9783 ( 
.A(n_9175),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9158),
.Y(n_9784)
);

AOI21xp5_ASAP7_75t_L g9785 ( 
.A1(n_9143),
.A2(n_247),
.B(n_248),
.Y(n_9785)
);

INVx1_ASAP7_75t_L g9786 ( 
.A(n_9683),
.Y(n_9786)
);

AND2x2_ASAP7_75t_L g9787 ( 
.A(n_9764),
.B(n_1218),
.Y(n_9787)
);

AOI211x1_ASAP7_75t_L g9788 ( 
.A1(n_9213),
.A2(n_250),
.B(n_247),
.C(n_249),
.Y(n_9788)
);

AO31x2_ASAP7_75t_L g9789 ( 
.A1(n_9666),
.A2(n_9114),
.A3(n_9250),
.B(n_9191),
.Y(n_9789)
);

OR2x2_ASAP7_75t_L g9790 ( 
.A(n_9688),
.B(n_1219),
.Y(n_9790)
);

AOI21xp5_ASAP7_75t_L g9791 ( 
.A1(n_9138),
.A2(n_249),
.B(n_250),
.Y(n_9791)
);

AOI21xp5_ASAP7_75t_L g9792 ( 
.A1(n_9232),
.A2(n_249),
.B(n_250),
.Y(n_9792)
);

AOI21xp5_ASAP7_75t_L g9793 ( 
.A1(n_9232),
.A2(n_251),
.B(n_252),
.Y(n_9793)
);

AOI21xp5_ASAP7_75t_L g9794 ( 
.A1(n_9232),
.A2(n_251),
.B(n_252),
.Y(n_9794)
);

OAI21x1_ASAP7_75t_L g9795 ( 
.A1(n_9433),
.A2(n_252),
.B(n_253),
.Y(n_9795)
);

OAI22xp5_ASAP7_75t_L g9796 ( 
.A1(n_9268),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_9796)
);

AOI21xp5_ASAP7_75t_L g9797 ( 
.A1(n_9257),
.A2(n_253),
.B(n_254),
.Y(n_9797)
);

NAND2xp5_ASAP7_75t_L g9798 ( 
.A(n_9242),
.B(n_1220),
.Y(n_9798)
);

INVx5_ASAP7_75t_L g9799 ( 
.A(n_9626),
.Y(n_9799)
);

AO21x2_ASAP7_75t_L g9800 ( 
.A1(n_9111),
.A2(n_254),
.B(n_255),
.Y(n_9800)
);

OAI21xp5_ASAP7_75t_L g9801 ( 
.A1(n_9271),
.A2(n_255),
.B(n_256),
.Y(n_9801)
);

INVx2_ASAP7_75t_L g9802 ( 
.A(n_9374),
.Y(n_9802)
);

HB1xp67_ASAP7_75t_L g9803 ( 
.A(n_9302),
.Y(n_9803)
);

AOI21x1_ASAP7_75t_L g9804 ( 
.A1(n_9468),
.A2(n_256),
.B(n_257),
.Y(n_9804)
);

OAI21xp5_ASAP7_75t_L g9805 ( 
.A1(n_9113),
.A2(n_256),
.B(n_257),
.Y(n_9805)
);

AOI22xp33_ASAP7_75t_L g9806 ( 
.A1(n_9332),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_9806)
);

AND2x2_ASAP7_75t_L g9807 ( 
.A(n_9766),
.B(n_9697),
.Y(n_9807)
);

OAI21x1_ASAP7_75t_L g9808 ( 
.A1(n_9655),
.A2(n_258),
.B(n_259),
.Y(n_9808)
);

BUFx6f_ASAP7_75t_L g9809 ( 
.A(n_9139),
.Y(n_9809)
);

NAND2xp5_ASAP7_75t_L g9810 ( 
.A(n_9298),
.B(n_1220),
.Y(n_9810)
);

A2O1A1Ixp33_ASAP7_75t_L g9811 ( 
.A1(n_9129),
.A2(n_1222),
.B(n_1223),
.C(n_1221),
.Y(n_9811)
);

AOI21xp5_ASAP7_75t_L g9812 ( 
.A1(n_9165),
.A2(n_258),
.B(n_260),
.Y(n_9812)
);

AOI21x1_ASAP7_75t_L g9813 ( 
.A1(n_9657),
.A2(n_260),
.B(n_261),
.Y(n_9813)
);

OAI21x1_ASAP7_75t_SL g9814 ( 
.A1(n_9140),
.A2(n_260),
.B(n_261),
.Y(n_9814)
);

OAI21xp5_ASAP7_75t_L g9815 ( 
.A1(n_9659),
.A2(n_262),
.B(n_263),
.Y(n_9815)
);

AOI211x1_ASAP7_75t_L g9816 ( 
.A1(n_9406),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_9816)
);

OAI21xp5_ASAP7_75t_L g9817 ( 
.A1(n_9663),
.A2(n_262),
.B(n_263),
.Y(n_9817)
);

INVx2_ASAP7_75t_L g9818 ( 
.A(n_9177),
.Y(n_9818)
);

A2O1A1Ixp33_ASAP7_75t_L g9819 ( 
.A1(n_9367),
.A2(n_1222),
.B(n_1223),
.C(n_1221),
.Y(n_9819)
);

BUFx3_ASAP7_75t_L g9820 ( 
.A(n_9125),
.Y(n_9820)
);

NAND2xp5_ASAP7_75t_SL g9821 ( 
.A(n_9134),
.B(n_1224),
.Y(n_9821)
);

AOI21xp33_ASAP7_75t_L g9822 ( 
.A1(n_9658),
.A2(n_264),
.B(n_265),
.Y(n_9822)
);

AOI21xp33_ASAP7_75t_L g9823 ( 
.A1(n_9691),
.A2(n_264),
.B(n_265),
.Y(n_9823)
);

INVx1_ASAP7_75t_SL g9824 ( 
.A(n_9270),
.Y(n_9824)
);

OAI21xp5_ASAP7_75t_L g9825 ( 
.A1(n_9664),
.A2(n_265),
.B(n_266),
.Y(n_9825)
);

AND2x4_ASAP7_75t_L g9826 ( 
.A(n_9119),
.B(n_1224),
.Y(n_9826)
);

NAND2xp5_ASAP7_75t_L g9827 ( 
.A(n_9193),
.B(n_1225),
.Y(n_9827)
);

AOI21xp5_ASAP7_75t_L g9828 ( 
.A1(n_9770),
.A2(n_266),
.B(n_267),
.Y(n_9828)
);

NOR2x1_ASAP7_75t_SL g9829 ( 
.A(n_9719),
.B(n_1225),
.Y(n_9829)
);

INVx1_ASAP7_75t_L g9830 ( 
.A(n_9727),
.Y(n_9830)
);

AOI21xp33_ASAP7_75t_L g9831 ( 
.A1(n_9713),
.A2(n_266),
.B(n_267),
.Y(n_9831)
);

INVx1_ASAP7_75t_L g9832 ( 
.A(n_9755),
.Y(n_9832)
);

BUFx4_ASAP7_75t_SL g9833 ( 
.A(n_9504),
.Y(n_9833)
);

OAI21x1_ASAP7_75t_L g9834 ( 
.A1(n_9671),
.A2(n_268),
.B(n_269),
.Y(n_9834)
);

OAI21x1_ASAP7_75t_L g9835 ( 
.A1(n_9673),
.A2(n_268),
.B(n_269),
.Y(n_9835)
);

O2A1O1Ixp33_ASAP7_75t_L g9836 ( 
.A1(n_9239),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_9836)
);

AOI21xp5_ASAP7_75t_L g9837 ( 
.A1(n_9775),
.A2(n_270),
.B(n_271),
.Y(n_9837)
);

NAND2x1p5_ASAP7_75t_L g9838 ( 
.A(n_9515),
.B(n_1226),
.Y(n_9838)
);

NAND2xp5_ASAP7_75t_L g9839 ( 
.A(n_9171),
.B(n_9462),
.Y(n_9839)
);

NAND2xp5_ASAP7_75t_SL g9840 ( 
.A(n_9251),
.B(n_1226),
.Y(n_9840)
);

OAI21x1_ASAP7_75t_L g9841 ( 
.A1(n_9677),
.A2(n_271),
.B(n_272),
.Y(n_9841)
);

BUFx2_ASAP7_75t_L g9842 ( 
.A(n_9368),
.Y(n_9842)
);

NAND2xp5_ASAP7_75t_SL g9843 ( 
.A(n_9678),
.B(n_1227),
.Y(n_9843)
);

BUFx12f_ASAP7_75t_L g9844 ( 
.A(n_9364),
.Y(n_9844)
);

CKINVDCx5p33_ASAP7_75t_R g9845 ( 
.A(n_9725),
.Y(n_9845)
);

OAI21xp5_ASAP7_75t_L g9846 ( 
.A1(n_9680),
.A2(n_271),
.B(n_272),
.Y(n_9846)
);

A2O1A1Ixp33_ASAP7_75t_L g9847 ( 
.A1(n_9445),
.A2(n_1228),
.B(n_1229),
.C(n_1227),
.Y(n_9847)
);

OAI21x1_ASAP7_75t_L g9848 ( 
.A1(n_9685),
.A2(n_272),
.B(n_273),
.Y(n_9848)
);

OAI21x1_ASAP7_75t_L g9849 ( 
.A1(n_9693),
.A2(n_273),
.B(n_274),
.Y(n_9849)
);

INVx2_ASAP7_75t_L g9850 ( 
.A(n_9200),
.Y(n_9850)
);

OAI21x1_ASAP7_75t_SL g9851 ( 
.A1(n_9648),
.A2(n_274),
.B(n_275),
.Y(n_9851)
);

OAI21x1_ASAP7_75t_L g9852 ( 
.A1(n_9696),
.A2(n_9709),
.B(n_9698),
.Y(n_9852)
);

AND2x2_ASAP7_75t_L g9853 ( 
.A(n_9771),
.B(n_1228),
.Y(n_9853)
);

NAND2xp5_ASAP7_75t_L g9854 ( 
.A(n_9405),
.B(n_1229),
.Y(n_9854)
);

INVx1_ASAP7_75t_SL g9855 ( 
.A(n_9668),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_9758),
.Y(n_9856)
);

INVx2_ASAP7_75t_SL g9857 ( 
.A(n_9181),
.Y(n_9857)
);

INVx2_ASAP7_75t_L g9858 ( 
.A(n_9202),
.Y(n_9858)
);

AOI21xp5_ASAP7_75t_L g9859 ( 
.A1(n_9716),
.A2(n_9731),
.B(n_9724),
.Y(n_9859)
);

AOI21xp5_ASAP7_75t_L g9860 ( 
.A1(n_9732),
.A2(n_275),
.B(n_276),
.Y(n_9860)
);

OAI21x1_ASAP7_75t_L g9861 ( 
.A1(n_9738),
.A2(n_275),
.B(n_276),
.Y(n_9861)
);

OAI21xp33_ASAP7_75t_SL g9862 ( 
.A1(n_9768),
.A2(n_1232),
.B(n_1231),
.Y(n_9862)
);

INVx2_ASAP7_75t_L g9863 ( 
.A(n_9209),
.Y(n_9863)
);

O2A1O1Ixp5_ASAP7_75t_L g9864 ( 
.A1(n_9726),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_9864)
);

A2O1A1Ixp33_ASAP7_75t_L g9865 ( 
.A1(n_9571),
.A2(n_1233),
.B(n_1234),
.C(n_1232),
.Y(n_9865)
);

AND2x2_ASAP7_75t_L g9866 ( 
.A(n_9552),
.B(n_1233),
.Y(n_9866)
);

O2A1O1Ixp5_ASAP7_75t_L g9867 ( 
.A1(n_9729),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_9867)
);

OAI21x1_ASAP7_75t_L g9868 ( 
.A1(n_9740),
.A2(n_279),
.B(n_280),
.Y(n_9868)
);

BUFx2_ASAP7_75t_L g9869 ( 
.A(n_9174),
.Y(n_9869)
);

NAND2xp5_ASAP7_75t_L g9870 ( 
.A(n_9237),
.B(n_1235),
.Y(n_9870)
);

INVxp67_ASAP7_75t_L g9871 ( 
.A(n_9151),
.Y(n_9871)
);

INVx2_ASAP7_75t_L g9872 ( 
.A(n_9236),
.Y(n_9872)
);

AOI21xp5_ASAP7_75t_L g9873 ( 
.A1(n_9742),
.A2(n_279),
.B(n_280),
.Y(n_9873)
);

AOI21xp5_ASAP7_75t_L g9874 ( 
.A1(n_9749),
.A2(n_9752),
.B(n_9274),
.Y(n_9874)
);

INVx1_ASAP7_75t_SL g9875 ( 
.A(n_9706),
.Y(n_9875)
);

OAI21xp5_ASAP7_75t_L g9876 ( 
.A1(n_9351),
.A2(n_280),
.B(n_281),
.Y(n_9876)
);

NAND2xp5_ASAP7_75t_SL g9877 ( 
.A(n_9184),
.B(n_1235),
.Y(n_9877)
);

AOI21xp5_ASAP7_75t_L g9878 ( 
.A1(n_9343),
.A2(n_281),
.B(n_282),
.Y(n_9878)
);

AOI221xp5_ASAP7_75t_L g9879 ( 
.A1(n_9258),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.C(n_284),
.Y(n_9879)
);

AND2x6_ASAP7_75t_L g9880 ( 
.A(n_9603),
.B(n_1236),
.Y(n_9880)
);

INVx2_ASAP7_75t_L g9881 ( 
.A(n_9247),
.Y(n_9881)
);

NAND2xp5_ASAP7_75t_L g9882 ( 
.A(n_9599),
.B(n_1236),
.Y(n_9882)
);

OAI21x1_ASAP7_75t_L g9883 ( 
.A1(n_9219),
.A2(n_282),
.B(n_283),
.Y(n_9883)
);

CKINVDCx8_ASAP7_75t_R g9884 ( 
.A(n_9614),
.Y(n_9884)
);

NAND2xp5_ASAP7_75t_L g9885 ( 
.A(n_9595),
.B(n_9185),
.Y(n_9885)
);

AND2x2_ASAP7_75t_L g9886 ( 
.A(n_9255),
.B(n_1237),
.Y(n_9886)
);

OAI21x1_ASAP7_75t_L g9887 ( 
.A1(n_9233),
.A2(n_284),
.B(n_285),
.Y(n_9887)
);

BUFx12f_ASAP7_75t_L g9888 ( 
.A(n_9404),
.Y(n_9888)
);

AND2x2_ASAP7_75t_L g9889 ( 
.A(n_9259),
.B(n_1238),
.Y(n_9889)
);

AO21x1_ASAP7_75t_L g9890 ( 
.A1(n_9389),
.A2(n_284),
.B(n_285),
.Y(n_9890)
);

AOI21x1_ASAP7_75t_L g9891 ( 
.A1(n_9382),
.A2(n_285),
.B(n_286),
.Y(n_9891)
);

NAND2xp5_ASAP7_75t_L g9892 ( 
.A(n_9132),
.B(n_1239),
.Y(n_9892)
);

AOI21xp5_ASAP7_75t_L g9893 ( 
.A1(n_9448),
.A2(n_9155),
.B(n_9301),
.Y(n_9893)
);

INVx1_ASAP7_75t_L g9894 ( 
.A(n_9272),
.Y(n_9894)
);

INVx1_ASAP7_75t_L g9895 ( 
.A(n_9295),
.Y(n_9895)
);

BUFx4_ASAP7_75t_SL g9896 ( 
.A(n_9568),
.Y(n_9896)
);

NAND2xp5_ASAP7_75t_L g9897 ( 
.A(n_9201),
.B(n_1239),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_SL g9898 ( 
.A(n_9290),
.B(n_1240),
.Y(n_9898)
);

AO31x2_ASAP7_75t_L g9899 ( 
.A1(n_9417),
.A2(n_288),
.A3(n_286),
.B(n_287),
.Y(n_9899)
);

NOR2xp67_ASAP7_75t_L g9900 ( 
.A(n_9216),
.B(n_286),
.Y(n_9900)
);

NOR2xp33_ASAP7_75t_SL g9901 ( 
.A(n_9526),
.B(n_9734),
.Y(n_9901)
);

OAI21x1_ASAP7_75t_L g9902 ( 
.A1(n_9245),
.A2(n_287),
.B(n_288),
.Y(n_9902)
);

NAND2xp5_ASAP7_75t_L g9903 ( 
.A(n_9205),
.B(n_1241),
.Y(n_9903)
);

OAI21x1_ASAP7_75t_L g9904 ( 
.A1(n_9311),
.A2(n_287),
.B(n_288),
.Y(n_9904)
);

A2O1A1Ixp33_ASAP7_75t_L g9905 ( 
.A1(n_9737),
.A2(n_1245),
.B(n_1246),
.C(n_1243),
.Y(n_9905)
);

OR2x2_ASAP7_75t_L g9906 ( 
.A(n_9313),
.B(n_1243),
.Y(n_9906)
);

INVx2_ASAP7_75t_SL g9907 ( 
.A(n_9320),
.Y(n_9907)
);

BUFx3_ASAP7_75t_L g9908 ( 
.A(n_9152),
.Y(n_9908)
);

AND2x2_ASAP7_75t_L g9909 ( 
.A(n_9396),
.B(n_1245),
.Y(n_9909)
);

NAND2xp5_ASAP7_75t_L g9910 ( 
.A(n_9222),
.B(n_9224),
.Y(n_9910)
);

AND3x4_ASAP7_75t_L g9911 ( 
.A(n_9493),
.B(n_289),
.C(n_290),
.Y(n_9911)
);

NAND2xp5_ASAP7_75t_L g9912 ( 
.A(n_9225),
.B(n_1247),
.Y(n_9912)
);

NAND2xp5_ASAP7_75t_L g9913 ( 
.A(n_9285),
.B(n_1247),
.Y(n_9913)
);

NAND2xp5_ASAP7_75t_L g9914 ( 
.A(n_9291),
.B(n_1248),
.Y(n_9914)
);

OAI21x1_ASAP7_75t_L g9915 ( 
.A1(n_9538),
.A2(n_289),
.B(n_290),
.Y(n_9915)
);

INVx3_ASAP7_75t_L g9916 ( 
.A(n_9139),
.Y(n_9916)
);

OAI21x1_ASAP7_75t_L g9917 ( 
.A1(n_9353),
.A2(n_289),
.B(n_290),
.Y(n_9917)
);

AOI21xp5_ASAP7_75t_L g9918 ( 
.A1(n_9617),
.A2(n_291),
.B(n_292),
.Y(n_9918)
);

AOI21xp5_ASAP7_75t_L g9919 ( 
.A1(n_9148),
.A2(n_291),
.B(n_292),
.Y(n_9919)
);

AOI21xp5_ASAP7_75t_L g9920 ( 
.A1(n_9148),
.A2(n_291),
.B(n_292),
.Y(n_9920)
);

OA21x2_ASAP7_75t_L g9921 ( 
.A1(n_9582),
.A2(n_293),
.B(n_294),
.Y(n_9921)
);

AOI21xp5_ASAP7_75t_L g9922 ( 
.A1(n_9675),
.A2(n_293),
.B(n_294),
.Y(n_9922)
);

INVx2_ASAP7_75t_L g9923 ( 
.A(n_9410),
.Y(n_9923)
);

AOI21x1_ASAP7_75t_L g9924 ( 
.A1(n_9197),
.A2(n_293),
.B(n_294),
.Y(n_9924)
);

INVx2_ASAP7_75t_L g9925 ( 
.A(n_9423),
.Y(n_9925)
);

AND2x2_ASAP7_75t_L g9926 ( 
.A(n_9451),
.B(n_1248),
.Y(n_9926)
);

OAI21x1_ASAP7_75t_L g9927 ( 
.A1(n_9546),
.A2(n_295),
.B(n_296),
.Y(n_9927)
);

INVx1_ASAP7_75t_L g9928 ( 
.A(n_9460),
.Y(n_9928)
);

A2O1A1Ixp33_ASAP7_75t_L g9929 ( 
.A1(n_9450),
.A2(n_1250),
.B(n_1251),
.C(n_1249),
.Y(n_9929)
);

INVx1_ASAP7_75t_L g9930 ( 
.A(n_9470),
.Y(n_9930)
);

NAND2xp5_ASAP7_75t_L g9931 ( 
.A(n_9294),
.B(n_1249),
.Y(n_9931)
);

AOI21xp5_ASAP7_75t_L g9932 ( 
.A1(n_9684),
.A2(n_9760),
.B(n_9701),
.Y(n_9932)
);

AND2x2_ASAP7_75t_L g9933 ( 
.A(n_9491),
.B(n_1250),
.Y(n_9933)
);

NOR2xp33_ASAP7_75t_L g9934 ( 
.A(n_9217),
.B(n_1252),
.Y(n_9934)
);

NAND2xp5_ASAP7_75t_L g9935 ( 
.A(n_9296),
.B(n_1253),
.Y(n_9935)
);

NAND2xp5_ASAP7_75t_L g9936 ( 
.A(n_9328),
.B(n_1254),
.Y(n_9936)
);

BUFx3_ASAP7_75t_L g9937 ( 
.A(n_9324),
.Y(n_9937)
);

NAND2xp5_ASAP7_75t_L g9938 ( 
.A(n_9350),
.B(n_1255),
.Y(n_9938)
);

OAI21x1_ASAP7_75t_L g9939 ( 
.A1(n_9362),
.A2(n_295),
.B(n_296),
.Y(n_9939)
);

OAI22xp5_ASAP7_75t_L g9940 ( 
.A1(n_9670),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_9940)
);

OAI21x1_ASAP7_75t_L g9941 ( 
.A1(n_9676),
.A2(n_297),
.B(n_298),
.Y(n_9941)
);

NAND2xp5_ASAP7_75t_L g9942 ( 
.A(n_9710),
.B(n_1256),
.Y(n_9942)
);

AOI21x1_ASAP7_75t_L g9943 ( 
.A1(n_9256),
.A2(n_297),
.B(n_298),
.Y(n_9943)
);

BUFx4f_ASAP7_75t_L g9944 ( 
.A(n_9275),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_9499),
.Y(n_9945)
);

INVx1_ASAP7_75t_L g9946 ( 
.A(n_9748),
.Y(n_9946)
);

INVx2_ASAP7_75t_L g9947 ( 
.A(n_9751),
.Y(n_9947)
);

INVx4_ASAP7_75t_L g9948 ( 
.A(n_9331),
.Y(n_9948)
);

HB1xp67_ASAP7_75t_L g9949 ( 
.A(n_9577),
.Y(n_9949)
);

AND2x2_ASAP7_75t_SL g9950 ( 
.A(n_9136),
.B(n_298),
.Y(n_9950)
);

AOI21xp5_ASAP7_75t_L g9951 ( 
.A1(n_9769),
.A2(n_299),
.B(n_300),
.Y(n_9951)
);

INVx1_ASAP7_75t_L g9952 ( 
.A(n_9400),
.Y(n_9952)
);

NOR2xp33_ASAP7_75t_L g9953 ( 
.A(n_9388),
.B(n_1257),
.Y(n_9953)
);

OAI21x1_ASAP7_75t_L g9954 ( 
.A1(n_9402),
.A2(n_299),
.B(n_300),
.Y(n_9954)
);

OAI21x1_ASAP7_75t_SL g9955 ( 
.A1(n_9338),
.A2(n_301),
.B(n_302),
.Y(n_9955)
);

OAI21x1_ASAP7_75t_L g9956 ( 
.A1(n_9425),
.A2(n_301),
.B(n_302),
.Y(n_9956)
);

BUFx6f_ASAP7_75t_L g9957 ( 
.A(n_9243),
.Y(n_9957)
);

AOI21xp33_ASAP7_75t_L g9958 ( 
.A1(n_9168),
.A2(n_303),
.B(n_304),
.Y(n_9958)
);

AOI21xp5_ASAP7_75t_L g9959 ( 
.A1(n_9774),
.A2(n_303),
.B(n_304),
.Y(n_9959)
);

INVxp67_ASAP7_75t_L g9960 ( 
.A(n_9565),
.Y(n_9960)
);

AOI21xp5_ASAP7_75t_L g9961 ( 
.A1(n_9203),
.A2(n_9588),
.B(n_9602),
.Y(n_9961)
);

BUFx2_ASAP7_75t_L g9962 ( 
.A(n_9557),
.Y(n_9962)
);

CKINVDCx5p33_ASAP7_75t_R g9963 ( 
.A(n_9348),
.Y(n_9963)
);

AOI21xp33_ASAP7_75t_L g9964 ( 
.A1(n_9496),
.A2(n_303),
.B(n_305),
.Y(n_9964)
);

AND2x2_ASAP7_75t_L g9965 ( 
.A(n_9590),
.B(n_1258),
.Y(n_9965)
);

OAI21xp5_ASAP7_75t_L g9966 ( 
.A1(n_9398),
.A2(n_305),
.B(n_306),
.Y(n_9966)
);

AND2x2_ASAP7_75t_L g9967 ( 
.A(n_9681),
.B(n_1258),
.Y(n_9967)
);

OAI22xp5_ASAP7_75t_L g9968 ( 
.A1(n_9686),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_9968)
);

OAI22xp5_ASAP7_75t_L g9969 ( 
.A1(n_9220),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_9969)
);

NOR2xp67_ASAP7_75t_L g9970 ( 
.A(n_9315),
.B(n_307),
.Y(n_9970)
);

AOI21xp5_ASAP7_75t_L g9971 ( 
.A1(n_9203),
.A2(n_309),
.B(n_310),
.Y(n_9971)
);

AOI21x1_ASAP7_75t_L g9972 ( 
.A1(n_9264),
.A2(n_310),
.B(n_311),
.Y(n_9972)
);

NAND2xp5_ASAP7_75t_L g9973 ( 
.A(n_9471),
.B(n_1259),
.Y(n_9973)
);

AO21x2_ASAP7_75t_L g9974 ( 
.A1(n_9682),
.A2(n_310),
.B(n_311),
.Y(n_9974)
);

INVx2_ASAP7_75t_L g9975 ( 
.A(n_9481),
.Y(n_9975)
);

NAND2xp5_ASAP7_75t_L g9976 ( 
.A(n_9702),
.B(n_1259),
.Y(n_9976)
);

NAND2xp5_ASAP7_75t_L g9977 ( 
.A(n_9735),
.B(n_1260),
.Y(n_9977)
);

AOI21xp5_ASAP7_75t_L g9978 ( 
.A1(n_9289),
.A2(n_311),
.B(n_312),
.Y(n_9978)
);

A2O1A1Ixp33_ASAP7_75t_L g9979 ( 
.A1(n_9443),
.A2(n_1261),
.B(n_1263),
.C(n_1260),
.Y(n_9979)
);

OAI21xp5_ASAP7_75t_L g9980 ( 
.A1(n_9153),
.A2(n_312),
.B(n_313),
.Y(n_9980)
);

OAI21x1_ASAP7_75t_L g9981 ( 
.A1(n_9426),
.A2(n_312),
.B(n_313),
.Y(n_9981)
);

AND2x2_ASAP7_75t_L g9982 ( 
.A(n_9498),
.B(n_1261),
.Y(n_9982)
);

AOI21xp5_ASAP7_75t_L g9983 ( 
.A1(n_9318),
.A2(n_313),
.B(n_314),
.Y(n_9983)
);

AO21x2_ASAP7_75t_L g9984 ( 
.A1(n_9708),
.A2(n_9754),
.B(n_9314),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9317),
.Y(n_9985)
);

OAI21x1_ASAP7_75t_L g9986 ( 
.A1(n_9427),
.A2(n_315),
.B(n_316),
.Y(n_9986)
);

INVx2_ASAP7_75t_SL g9987 ( 
.A(n_9390),
.Y(n_9987)
);

INVx2_ASAP7_75t_SL g9988 ( 
.A(n_9497),
.Y(n_9988)
);

NOR2x1_ASAP7_75t_SL g9989 ( 
.A(n_9278),
.B(n_1263),
.Y(n_9989)
);

AOI21xp5_ASAP7_75t_L g9990 ( 
.A1(n_9207),
.A2(n_315),
.B(n_316),
.Y(n_9990)
);

NAND2xp5_ASAP7_75t_L g9991 ( 
.A(n_9669),
.B(n_1264),
.Y(n_9991)
);

BUFx5_ASAP7_75t_L g9992 ( 
.A(n_9626),
.Y(n_9992)
);

INVx1_ASAP7_75t_SL g9993 ( 
.A(n_9539),
.Y(n_9993)
);

AND2x4_ASAP7_75t_L g9994 ( 
.A(n_9408),
.B(n_1264),
.Y(n_9994)
);

INVx1_ASAP7_75t_L g9995 ( 
.A(n_9347),
.Y(n_9995)
);

OAI21x1_ASAP7_75t_SL g9996 ( 
.A1(n_9305),
.A2(n_315),
.B(n_316),
.Y(n_9996)
);

OAI21x1_ASAP7_75t_L g9997 ( 
.A1(n_9428),
.A2(n_9455),
.B(n_9442),
.Y(n_9997)
);

AOI21xp5_ASAP7_75t_L g9998 ( 
.A1(n_9429),
.A2(n_317),
.B(n_318),
.Y(n_9998)
);

INVx3_ASAP7_75t_L g9999 ( 
.A(n_9243),
.Y(n_9999)
);

NAND2xp5_ASAP7_75t_L g10000 ( 
.A(n_9718),
.B(n_1265),
.Y(n_10000)
);

OAI21x1_ASAP7_75t_L g10001 ( 
.A1(n_9464),
.A2(n_317),
.B(n_318),
.Y(n_10001)
);

NAND2x1p5_ASAP7_75t_L g10002 ( 
.A(n_9384),
.B(n_1265),
.Y(n_10002)
);

OAI21x1_ASAP7_75t_L g10003 ( 
.A1(n_9469),
.A2(n_317),
.B(n_318),
.Y(n_10003)
);

AO21x2_ASAP7_75t_L g10004 ( 
.A1(n_9344),
.A2(n_319),
.B(n_320),
.Y(n_10004)
);

AOI21xp5_ASAP7_75t_L g10005 ( 
.A1(n_9622),
.A2(n_319),
.B(n_320),
.Y(n_10005)
);

OAI21x1_ASAP7_75t_L g10006 ( 
.A1(n_9342),
.A2(n_319),
.B(n_320),
.Y(n_10006)
);

AOI21xp33_ASAP7_75t_L g10007 ( 
.A1(n_9420),
.A2(n_9308),
.B(n_9373),
.Y(n_10007)
);

OAI21x1_ASAP7_75t_L g10008 ( 
.A1(n_9475),
.A2(n_321),
.B(n_322),
.Y(n_10008)
);

AOI21xp5_ASAP7_75t_L g10009 ( 
.A1(n_9567),
.A2(n_321),
.B(n_322),
.Y(n_10009)
);

AOI21xp5_ASAP7_75t_L g10010 ( 
.A1(n_9583),
.A2(n_321),
.B(n_322),
.Y(n_10010)
);

NAND2xp5_ASAP7_75t_L g10011 ( 
.A(n_9283),
.B(n_1266),
.Y(n_10011)
);

AOI221x1_ASAP7_75t_L g10012 ( 
.A1(n_9561),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_326),
.Y(n_10012)
);

NAND2xp5_ASAP7_75t_SL g10013 ( 
.A(n_9112),
.B(n_1267),
.Y(n_10013)
);

INVx1_ASAP7_75t_L g10014 ( 
.A(n_9394),
.Y(n_10014)
);

AOI221xp5_ASAP7_75t_SL g10015 ( 
.A1(n_9508),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_327),
.Y(n_10015)
);

BUFx3_ASAP7_75t_L g10016 ( 
.A(n_9324),
.Y(n_10016)
);

NAND2xp5_ASAP7_75t_L g10017 ( 
.A(n_9117),
.B(n_9128),
.Y(n_10017)
);

INVx1_ASAP7_75t_L g10018 ( 
.A(n_9434),
.Y(n_10018)
);

OAI21xp5_ASAP7_75t_L g10019 ( 
.A1(n_9145),
.A2(n_323),
.B(n_324),
.Y(n_10019)
);

A2O1A1Ixp33_ASAP7_75t_L g10020 ( 
.A1(n_9141),
.A2(n_1268),
.B(n_1269),
.C(n_1267),
.Y(n_10020)
);

BUFx6f_ASAP7_75t_L g10021 ( 
.A(n_9661),
.Y(n_10021)
);

NAND2xp5_ASAP7_75t_L g10022 ( 
.A(n_9730),
.B(n_1268),
.Y(n_10022)
);

BUFx6f_ASAP7_75t_L g10023 ( 
.A(n_9661),
.Y(n_10023)
);

OAI21xp5_ASAP7_75t_SL g10024 ( 
.A1(n_9176),
.A2(n_325),
.B(n_327),
.Y(n_10024)
);

NOR2xp33_ASAP7_75t_R g10025 ( 
.A(n_9211),
.B(n_327),
.Y(n_10025)
);

OAI21xp5_ASAP7_75t_L g10026 ( 
.A1(n_9337),
.A2(n_328),
.B(n_329),
.Y(n_10026)
);

OAI21x1_ASAP7_75t_L g10027 ( 
.A1(n_9480),
.A2(n_328),
.B(n_329),
.Y(n_10027)
);

BUFx2_ASAP7_75t_L g10028 ( 
.A(n_9392),
.Y(n_10028)
);

NOR2xp33_ASAP7_75t_L g10029 ( 
.A(n_9570),
.B(n_1270),
.Y(n_10029)
);

O2A1O1Ixp5_ASAP7_75t_L g10030 ( 
.A1(n_9316),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_10030)
);

OAI21xp5_ASAP7_75t_L g10031 ( 
.A1(n_9293),
.A2(n_330),
.B(n_331),
.Y(n_10031)
);

OAI21x1_ASAP7_75t_L g10032 ( 
.A1(n_9503),
.A2(n_330),
.B(n_331),
.Y(n_10032)
);

AND2x6_ASAP7_75t_L g10033 ( 
.A(n_9319),
.B(n_1271),
.Y(n_10033)
);

OAI21xp5_ASAP7_75t_L g10034 ( 
.A1(n_9303),
.A2(n_331),
.B(n_332),
.Y(n_10034)
);

AOI21xp5_ASAP7_75t_L g10035 ( 
.A1(n_9585),
.A2(n_9330),
.B(n_9414),
.Y(n_10035)
);

AOI21xp5_ASAP7_75t_L g10036 ( 
.A1(n_9585),
.A2(n_332),
.B(n_333),
.Y(n_10036)
);

AOI22xp5_ASAP7_75t_L g10037 ( 
.A1(n_9332),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_10037)
);

NAND2xp5_ASAP7_75t_L g10038 ( 
.A(n_9773),
.B(n_1272),
.Y(n_10038)
);

AND2x2_ASAP7_75t_L g10039 ( 
.A(n_9180),
.B(n_1272),
.Y(n_10039)
);

NAND3xp33_ASAP7_75t_L g10040 ( 
.A(n_9547),
.B(n_9210),
.C(n_9411),
.Y(n_10040)
);

NAND2xp5_ASAP7_75t_SL g10041 ( 
.A(n_9198),
.B(n_1273),
.Y(n_10041)
);

AND2x6_ASAP7_75t_L g10042 ( 
.A(n_9638),
.B(n_1273),
.Y(n_10042)
);

OR2x2_ASAP7_75t_L g10043 ( 
.A(n_9615),
.B(n_9192),
.Y(n_10043)
);

NAND2xp5_ASAP7_75t_L g10044 ( 
.A(n_9656),
.B(n_1274),
.Y(n_10044)
);

O2A1O1Ixp5_ASAP7_75t_L g10045 ( 
.A1(n_9336),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_10045)
);

NAND2xp5_ASAP7_75t_L g10046 ( 
.A(n_9662),
.B(n_1274),
.Y(n_10046)
);

AO31x2_ASAP7_75t_L g10047 ( 
.A1(n_9266),
.A2(n_337),
.A3(n_335),
.B(n_336),
.Y(n_10047)
);

BUFx4f_ASAP7_75t_L g10048 ( 
.A(n_9385),
.Y(n_10048)
);

OAI21x1_ASAP7_75t_L g10049 ( 
.A1(n_9507),
.A2(n_336),
.B(n_337),
.Y(n_10049)
);

NOR2xp67_ASAP7_75t_L g10050 ( 
.A(n_9704),
.B(n_336),
.Y(n_10050)
);

AND2x2_ASAP7_75t_L g10051 ( 
.A(n_9163),
.B(n_1276),
.Y(n_10051)
);

AOI21xp5_ASAP7_75t_L g10052 ( 
.A1(n_9560),
.A2(n_338),
.B(n_339),
.Y(n_10052)
);

BUFx3_ASAP7_75t_L g10053 ( 
.A(n_9339),
.Y(n_10053)
);

BUFx6f_ASAP7_75t_L g10054 ( 
.A(n_9667),
.Y(n_10054)
);

NAND2x1_ASAP7_75t_L g10055 ( 
.A(n_9626),
.B(n_1276),
.Y(n_10055)
);

AOI21x1_ASAP7_75t_L g10056 ( 
.A1(n_9378),
.A2(n_338),
.B(n_339),
.Y(n_10056)
);

OAI21x1_ASAP7_75t_SL g10057 ( 
.A1(n_9363),
.A2(n_338),
.B(n_339),
.Y(n_10057)
);

AOI21x1_ASAP7_75t_L g10058 ( 
.A1(n_9440),
.A2(n_340),
.B(n_341),
.Y(n_10058)
);

OAI22xp33_ASAP7_75t_L g10059 ( 
.A1(n_9359),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_10059)
);

AOI21x1_ASAP7_75t_L g10060 ( 
.A1(n_9665),
.A2(n_340),
.B(n_341),
.Y(n_10060)
);

OAI22x1_ASAP7_75t_L g10061 ( 
.A1(n_9652),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_10061)
);

AND2x2_ASAP7_75t_L g10062 ( 
.A(n_9627),
.B(n_1277),
.Y(n_10062)
);

AOI221xp5_ASAP7_75t_L g10063 ( 
.A1(n_9223),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.C(n_345),
.Y(n_10063)
);

BUFx2_ASAP7_75t_L g10064 ( 
.A(n_9449),
.Y(n_10064)
);

OAI21xp5_ASAP7_75t_L g10065 ( 
.A1(n_9489),
.A2(n_344),
.B(n_345),
.Y(n_10065)
);

OAI22xp5_ASAP7_75t_L g10066 ( 
.A1(n_9523),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_10066)
);

AOI21xp5_ASAP7_75t_L g10067 ( 
.A1(n_9354),
.A2(n_346),
.B(n_348),
.Y(n_10067)
);

NAND2xp5_ASAP7_75t_L g10068 ( 
.A(n_9672),
.B(n_1278),
.Y(n_10068)
);

AND2x4_ASAP7_75t_L g10069 ( 
.A(n_9502),
.B(n_1279),
.Y(n_10069)
);

OAI21xp5_ASAP7_75t_L g10070 ( 
.A1(n_9500),
.A2(n_348),
.B(n_349),
.Y(n_10070)
);

INVx1_ASAP7_75t_L g10071 ( 
.A(n_9435),
.Y(n_10071)
);

OAI21xp5_ASAP7_75t_L g10072 ( 
.A1(n_9553),
.A2(n_348),
.B(n_349),
.Y(n_10072)
);

OAI21x1_ASAP7_75t_SL g10073 ( 
.A1(n_9452),
.A2(n_349),
.B(n_350),
.Y(n_10073)
);

OAI21x1_ASAP7_75t_L g10074 ( 
.A1(n_9510),
.A2(n_350),
.B(n_351),
.Y(n_10074)
);

INVx1_ASAP7_75t_L g10075 ( 
.A(n_9436),
.Y(n_10075)
);

AO31x2_ASAP7_75t_L g10076 ( 
.A1(n_9643),
.A2(n_9551),
.A3(n_9592),
.B(n_9254),
.Y(n_10076)
);

NAND2xp5_ASAP7_75t_L g10077 ( 
.A(n_9689),
.B(n_1280),
.Y(n_10077)
);

OAI22x1_ASAP7_75t_L g10078 ( 
.A1(n_9267),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_10078)
);

CKINVDCx6p67_ASAP7_75t_R g10079 ( 
.A(n_9391),
.Y(n_10079)
);

AOI21x1_ASAP7_75t_L g10080 ( 
.A1(n_9700),
.A2(n_352),
.B(n_353),
.Y(n_10080)
);

OAI21x1_ASAP7_75t_L g10081 ( 
.A1(n_9525),
.A2(n_353),
.B(n_354),
.Y(n_10081)
);

BUFx6f_ASAP7_75t_L g10082 ( 
.A(n_9667),
.Y(n_10082)
);

AOI21xp5_ASAP7_75t_SL g10083 ( 
.A1(n_9587),
.A2(n_1281),
.B(n_1280),
.Y(n_10083)
);

OA22x2_ASAP7_75t_L g10084 ( 
.A1(n_9715),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_10084)
);

NAND2xp5_ASAP7_75t_L g10085 ( 
.A(n_9695),
.B(n_1281),
.Y(n_10085)
);

NAND2xp5_ASAP7_75t_L g10086 ( 
.A(n_9707),
.B(n_1282),
.Y(n_10086)
);

OAI21x1_ASAP7_75t_L g10087 ( 
.A1(n_9529),
.A2(n_354),
.B(n_355),
.Y(n_10087)
);

AND2x4_ASAP7_75t_L g10088 ( 
.A(n_9502),
.B(n_1282),
.Y(n_10088)
);

NAND2x1p5_ASAP7_75t_L g10089 ( 
.A(n_9401),
.B(n_9747),
.Y(n_10089)
);

OAI22x1_ASAP7_75t_L g10090 ( 
.A1(n_9379),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_10090)
);

BUFx2_ASAP7_75t_L g10091 ( 
.A(n_9591),
.Y(n_10091)
);

NOR2xp33_ASAP7_75t_L g10092 ( 
.A(n_9326),
.B(n_1283),
.Y(n_10092)
);

OAI21x1_ASAP7_75t_L g10093 ( 
.A1(n_9530),
.A2(n_356),
.B(n_357),
.Y(n_10093)
);

NAND2xp5_ASAP7_75t_SL g10094 ( 
.A(n_9244),
.B(n_1284),
.Y(n_10094)
);

O2A1O1Ixp5_ASAP7_75t_L g10095 ( 
.A1(n_9381),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_10095)
);

NOR2xp67_ASAP7_75t_L g10096 ( 
.A(n_9703),
.B(n_9549),
.Y(n_10096)
);

NAND2x1p5_ASAP7_75t_L g10097 ( 
.A(n_9479),
.B(n_1284),
.Y(n_10097)
);

AND2x2_ASAP7_75t_L g10098 ( 
.A(n_9260),
.B(n_9262),
.Y(n_10098)
);

AND2x4_ASAP7_75t_L g10099 ( 
.A(n_9333),
.B(n_1285),
.Y(n_10099)
);

BUFx2_ASAP7_75t_L g10100 ( 
.A(n_9497),
.Y(n_10100)
);

OAI21x1_ASAP7_75t_L g10101 ( 
.A1(n_9537),
.A2(n_358),
.B(n_359),
.Y(n_10101)
);

NAND2xp5_ASAP7_75t_L g10102 ( 
.A(n_9711),
.B(n_1286),
.Y(n_10102)
);

A2O1A1Ixp33_ASAP7_75t_L g10103 ( 
.A1(n_9157),
.A2(n_1288),
.B(n_1289),
.C(n_1287),
.Y(n_10103)
);

OAI22xp5_ASAP7_75t_L g10104 ( 
.A1(n_9161),
.A2(n_9412),
.B1(n_9221),
.B2(n_9569),
.Y(n_10104)
);

NAND2xp5_ASAP7_75t_L g10105 ( 
.A(n_9714),
.B(n_1288),
.Y(n_10105)
);

BUFx6f_ASAP7_75t_L g10106 ( 
.A(n_9765),
.Y(n_10106)
);

A2O1A1Ixp33_ASAP7_75t_L g10107 ( 
.A1(n_9660),
.A2(n_1291),
.B(n_1292),
.C(n_1290),
.Y(n_10107)
);

OAI21x1_ASAP7_75t_L g10108 ( 
.A1(n_9544),
.A2(n_358),
.B(n_359),
.Y(n_10108)
);

AND2x4_ASAP7_75t_L g10109 ( 
.A(n_9371),
.B(n_1290),
.Y(n_10109)
);

INVx1_ASAP7_75t_SL g10110 ( 
.A(n_9605),
.Y(n_10110)
);

AND2x2_ASAP7_75t_L g10111 ( 
.A(n_9142),
.B(n_1292),
.Y(n_10111)
);

AND3x2_ASAP7_75t_L g10112 ( 
.A(n_9519),
.B(n_359),
.C(n_360),
.Y(n_10112)
);

INVx2_ASAP7_75t_L g10113 ( 
.A(n_9506),
.Y(n_10113)
);

OA21x2_ASAP7_75t_L g10114 ( 
.A1(n_9584),
.A2(n_9441),
.B(n_9545),
.Y(n_10114)
);

NAND2xp5_ASAP7_75t_L g10115 ( 
.A(n_9717),
.B(n_1293),
.Y(n_10115)
);

O2A1O1Ixp5_ASAP7_75t_L g10116 ( 
.A1(n_9246),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_10116)
);

AOI21xp5_ASAP7_75t_L g10117 ( 
.A1(n_9355),
.A2(n_360),
.B(n_361),
.Y(n_10117)
);

AOI21xp5_ASAP7_75t_L g10118 ( 
.A1(n_9361),
.A2(n_361),
.B(n_362),
.Y(n_10118)
);

NOR2x1_ASAP7_75t_SL g10119 ( 
.A(n_9278),
.B(n_1293),
.Y(n_10119)
);

INVxp67_ASAP7_75t_L g10120 ( 
.A(n_9611),
.Y(n_10120)
);

NOR2x1_ASAP7_75t_L g10121 ( 
.A(n_9166),
.B(n_1294),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_SL g10122 ( 
.A(n_9692),
.B(n_1294),
.Y(n_10122)
);

AOI21xp5_ASAP7_75t_SL g10123 ( 
.A1(n_9306),
.A2(n_1296),
.B(n_1295),
.Y(n_10123)
);

O2A1O1Ixp33_ASAP7_75t_L g10124 ( 
.A1(n_9127),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_10124)
);

OAI21x1_ASAP7_75t_L g10125 ( 
.A1(n_9550),
.A2(n_9179),
.B(n_9173),
.Y(n_10125)
);

OAI21x1_ASAP7_75t_L g10126 ( 
.A1(n_9183),
.A2(n_363),
.B(n_364),
.Y(n_10126)
);

A2O1A1Ixp33_ASAP7_75t_L g10127 ( 
.A1(n_9743),
.A2(n_1297),
.B(n_1298),
.C(n_1295),
.Y(n_10127)
);

INVx2_ASAP7_75t_L g10128 ( 
.A(n_9528),
.Y(n_10128)
);

INVx1_ASAP7_75t_L g10129 ( 
.A(n_9444),
.Y(n_10129)
);

AO31x2_ASAP7_75t_L g10130 ( 
.A1(n_9325),
.A2(n_367),
.A3(n_365),
.B(n_366),
.Y(n_10130)
);

BUFx6f_ASAP7_75t_L g10131 ( 
.A(n_9765),
.Y(n_10131)
);

NAND2xp5_ASAP7_75t_L g10132 ( 
.A(n_9720),
.B(n_1298),
.Y(n_10132)
);

O2A1O1Ixp5_ASAP7_75t_L g10133 ( 
.A1(n_9253),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_10133)
);

AOI21x1_ASAP7_75t_L g10134 ( 
.A1(n_9722),
.A2(n_9736),
.B(n_9728),
.Y(n_10134)
);

OAI21xp5_ASAP7_75t_L g10135 ( 
.A1(n_9610),
.A2(n_367),
.B(n_368),
.Y(n_10135)
);

OAI21x1_ASAP7_75t_L g10136 ( 
.A1(n_9188),
.A2(n_368),
.B(n_369),
.Y(n_10136)
);

AOI21x1_ASAP7_75t_SL g10137 ( 
.A1(n_9649),
.A2(n_1301),
.B(n_1299),
.Y(n_10137)
);

OAI21x1_ASAP7_75t_L g10138 ( 
.A1(n_9190),
.A2(n_369),
.B(n_370),
.Y(n_10138)
);

INVx2_ASAP7_75t_L g10139 ( 
.A(n_9596),
.Y(n_10139)
);

OAI21x1_ASAP7_75t_L g10140 ( 
.A1(n_9204),
.A2(n_369),
.B(n_370),
.Y(n_10140)
);

NAND2x1p5_ASAP7_75t_L g10141 ( 
.A(n_9156),
.B(n_1299),
.Y(n_10141)
);

NAND2xp5_ASAP7_75t_L g10142 ( 
.A(n_9721),
.B(n_1301),
.Y(n_10142)
);

AOI21x1_ASAP7_75t_SL g10143 ( 
.A1(n_9601),
.A2(n_1303),
.B(n_1302),
.Y(n_10143)
);

NAND2xp5_ASAP7_75t_L g10144 ( 
.A(n_9723),
.B(n_1302),
.Y(n_10144)
);

NAND2xp5_ASAP7_75t_L g10145 ( 
.A(n_9733),
.B(n_1303),
.Y(n_10145)
);

A2O1A1Ixp33_ASAP7_75t_L g10146 ( 
.A1(n_9756),
.A2(n_1305),
.B(n_1306),
.C(n_1304),
.Y(n_10146)
);

INVx3_ASAP7_75t_L g10147 ( 
.A(n_9339),
.Y(n_10147)
);

OAI21x1_ASAP7_75t_L g10148 ( 
.A1(n_9214),
.A2(n_370),
.B(n_371),
.Y(n_10148)
);

NAND2xp5_ASAP7_75t_L g10149 ( 
.A(n_9745),
.B(n_1304),
.Y(n_10149)
);

AOI21xp5_ASAP7_75t_L g10150 ( 
.A1(n_9229),
.A2(n_371),
.B(n_372),
.Y(n_10150)
);

OAI21x1_ASAP7_75t_L g10151 ( 
.A1(n_9218),
.A2(n_372),
.B(n_373),
.Y(n_10151)
);

NAND2x1p5_ASAP7_75t_L g10152 ( 
.A(n_9593),
.B(n_1305),
.Y(n_10152)
);

BUFx4f_ASAP7_75t_L g10153 ( 
.A(n_9322),
.Y(n_10153)
);

OAI21xp5_ASAP7_75t_L g10154 ( 
.A1(n_9397),
.A2(n_372),
.B(n_373),
.Y(n_10154)
);

INVx1_ASAP7_75t_L g10155 ( 
.A(n_9457),
.Y(n_10155)
);

AO31x2_ASAP7_75t_L g10156 ( 
.A1(n_9421),
.A2(n_375),
.A3(n_373),
.B(n_374),
.Y(n_10156)
);

OAI21x1_ASAP7_75t_L g10157 ( 
.A1(n_9227),
.A2(n_374),
.B(n_375),
.Y(n_10157)
);

OA21x2_ASAP7_75t_L g10158 ( 
.A1(n_9238),
.A2(n_9282),
.B(n_9281),
.Y(n_10158)
);

AND2x2_ASAP7_75t_L g10159 ( 
.A(n_9149),
.B(n_1307),
.Y(n_10159)
);

BUFx6f_ASAP7_75t_L g10160 ( 
.A(n_9322),
.Y(n_10160)
);

NAND2xp5_ASAP7_75t_L g10161 ( 
.A(n_9750),
.B(n_1307),
.Y(n_10161)
);

OAI21x1_ASAP7_75t_L g10162 ( 
.A1(n_9580),
.A2(n_374),
.B(n_376),
.Y(n_10162)
);

OAI21x1_ASAP7_75t_L g10163 ( 
.A1(n_9235),
.A2(n_376),
.B(n_377),
.Y(n_10163)
);

OAI21xp5_ASAP7_75t_L g10164 ( 
.A1(n_9589),
.A2(n_376),
.B(n_377),
.Y(n_10164)
);

OAI21xp5_ASAP7_75t_L g10165 ( 
.A1(n_9555),
.A2(n_9300),
.B(n_9403),
.Y(n_10165)
);

OAI21xp5_ASAP7_75t_L g10166 ( 
.A1(n_9409),
.A2(n_377),
.B(n_378),
.Y(n_10166)
);

NOR2xp33_ASAP7_75t_L g10167 ( 
.A(n_9215),
.B(n_1308),
.Y(n_10167)
);

A2O1A1Ixp33_ASAP7_75t_L g10168 ( 
.A1(n_9699),
.A2(n_9772),
.B(n_9312),
.C(n_9231),
.Y(n_10168)
);

NAND2xp5_ASAP7_75t_L g10169 ( 
.A(n_9753),
.B(n_1308),
.Y(n_10169)
);

AND2x2_ASAP7_75t_L g10170 ( 
.A(n_9631),
.B(n_1309),
.Y(n_10170)
);

OAI21xp5_ASAP7_75t_L g10171 ( 
.A1(n_9208),
.A2(n_378),
.B(n_379),
.Y(n_10171)
);

OAI22x1_ASAP7_75t_L g10172 ( 
.A1(n_9612),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_10172)
);

OAI21x1_ASAP7_75t_L g10173 ( 
.A1(n_9212),
.A2(n_9277),
.B(n_9263),
.Y(n_10173)
);

NAND2xp5_ASAP7_75t_L g10174 ( 
.A(n_9767),
.B(n_1309),
.Y(n_10174)
);

NAND2xp5_ASAP7_75t_L g10175 ( 
.A(n_9757),
.B(n_1311),
.Y(n_10175)
);

AOI21xp5_ASAP7_75t_L g10176 ( 
.A1(n_9287),
.A2(n_380),
.B(n_381),
.Y(n_10176)
);

OR2x2_ASAP7_75t_L g10177 ( 
.A(n_9284),
.B(n_1312),
.Y(n_10177)
);

NOR2xp67_ASAP7_75t_L g10178 ( 
.A(n_9286),
.B(n_381),
.Y(n_10178)
);

OAI22x1_ASAP7_75t_L g10179 ( 
.A1(n_9562),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_10179)
);

INVx2_ASAP7_75t_L g10180 ( 
.A(n_9461),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_L g10181 ( 
.A(n_9759),
.B(n_1313),
.Y(n_10181)
);

AOI21xp5_ASAP7_75t_SL g10182 ( 
.A1(n_9472),
.A2(n_9621),
.B(n_9597),
.Y(n_10182)
);

NOR2xp33_ASAP7_75t_L g10183 ( 
.A(n_9647),
.B(n_1314),
.Y(n_10183)
);

INVx1_ASAP7_75t_L g10184 ( 
.A(n_9466),
.Y(n_10184)
);

AOI22xp5_ASAP7_75t_L g10185 ( 
.A1(n_9332),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_10185)
);

OAI21xp5_ASAP7_75t_L g10186 ( 
.A1(n_9488),
.A2(n_382),
.B(n_383),
.Y(n_10186)
);

AOI21x1_ASAP7_75t_L g10187 ( 
.A1(n_9516),
.A2(n_9370),
.B(n_9122),
.Y(n_10187)
);

INVx2_ASAP7_75t_SL g10188 ( 
.A(n_9647),
.Y(n_10188)
);

OAI21x1_ASAP7_75t_L g10189 ( 
.A1(n_9477),
.A2(n_384),
.B(n_385),
.Y(n_10189)
);

BUFx2_ASAP7_75t_L g10190 ( 
.A(n_9340),
.Y(n_10190)
);

AOI21x1_ASAP7_75t_L g10191 ( 
.A1(n_9304),
.A2(n_9327),
.B(n_9150),
.Y(n_10191)
);

AND2x4_ASAP7_75t_L g10192 ( 
.A(n_9288),
.B(n_9310),
.Y(n_10192)
);

OA22x2_ASAP7_75t_L g10193 ( 
.A1(n_9642),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_10193)
);

INVx2_ASAP7_75t_L g10194 ( 
.A(n_9467),
.Y(n_10194)
);

OAI22xp5_ASAP7_75t_L g10195 ( 
.A1(n_9377),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_10195)
);

OAI21xp5_ASAP7_75t_L g10196 ( 
.A1(n_9600),
.A2(n_386),
.B(n_388),
.Y(n_10196)
);

OAI21x1_ASAP7_75t_L g10197 ( 
.A1(n_9334),
.A2(n_388),
.B(n_389),
.Y(n_10197)
);

AOI21xp33_ASAP7_75t_L g10198 ( 
.A1(n_9521),
.A2(n_389),
.B(n_390),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_L g10199 ( 
.A(n_9763),
.B(n_1314),
.Y(n_10199)
);

BUFx3_ASAP7_75t_L g10200 ( 
.A(n_9321),
.Y(n_10200)
);

AO31x2_ASAP7_75t_L g10201 ( 
.A1(n_9679),
.A2(n_391),
.A3(n_389),
.B(n_390),
.Y(n_10201)
);

OAI21xp5_ASAP7_75t_L g10202 ( 
.A1(n_9608),
.A2(n_9625),
.B(n_9126),
.Y(n_10202)
);

OAI21xp5_ASAP7_75t_L g10203 ( 
.A1(n_9482),
.A2(n_390),
.B(n_391),
.Y(n_10203)
);

AOI21x1_ASAP7_75t_L g10204 ( 
.A1(n_9280),
.A2(n_9292),
.B(n_9240),
.Y(n_10204)
);

AND2x6_ASAP7_75t_L g10205 ( 
.A(n_9712),
.B(n_9739),
.Y(n_10205)
);

NAND2xp5_ASAP7_75t_L g10206 ( 
.A(n_9206),
.B(n_1315),
.Y(n_10206)
);

INVx1_ASAP7_75t_L g10207 ( 
.A(n_9575),
.Y(n_10207)
);

NAND2xp5_ASAP7_75t_L g10208 ( 
.A(n_9172),
.B(n_1315),
.Y(n_10208)
);

INVx1_ASAP7_75t_L g10209 ( 
.A(n_9341),
.Y(n_10209)
);

AO31x2_ASAP7_75t_L g10210 ( 
.A1(n_9744),
.A2(n_393),
.A3(n_391),
.B(n_392),
.Y(n_10210)
);

AOI21x1_ASAP7_75t_SL g10211 ( 
.A1(n_9307),
.A2(n_1317),
.B(n_1316),
.Y(n_10211)
);

OAI21x1_ASAP7_75t_L g10212 ( 
.A1(n_9346),
.A2(n_392),
.B(n_393),
.Y(n_10212)
);

AOI21xp5_ASAP7_75t_L g10213 ( 
.A1(n_9633),
.A2(n_393),
.B(n_394),
.Y(n_10213)
);

NAND2xp5_ASAP7_75t_L g10214 ( 
.A(n_9178),
.B(n_1316),
.Y(n_10214)
);

OAI21x1_ASAP7_75t_L g10215 ( 
.A1(n_9349),
.A2(n_9358),
.B(n_9357),
.Y(n_10215)
);

NAND2xp5_ASAP7_75t_SL g10216 ( 
.A(n_9532),
.B(n_1317),
.Y(n_10216)
);

NAND2xp5_ASAP7_75t_SL g10217 ( 
.A(n_9532),
.B(n_1318),
.Y(n_10217)
);

INVx2_ASAP7_75t_L g10218 ( 
.A(n_9360),
.Y(n_10218)
);

NAND2xp5_ASAP7_75t_L g10219 ( 
.A(n_9182),
.B(n_1318),
.Y(n_10219)
);

AOI21xp5_ASAP7_75t_L g10220 ( 
.A1(n_9487),
.A2(n_394),
.B(n_395),
.Y(n_10220)
);

OAI21xp33_ASAP7_75t_L g10221 ( 
.A1(n_9297),
.A2(n_394),
.B(n_395),
.Y(n_10221)
);

NAND3xp33_ASAP7_75t_L g10222 ( 
.A(n_9116),
.B(n_395),
.C(n_396),
.Y(n_10222)
);

OAI21x1_ASAP7_75t_L g10223 ( 
.A1(n_9618),
.A2(n_396),
.B(n_397),
.Y(n_10223)
);

NOR2x1_ASAP7_75t_R g10224 ( 
.A(n_9437),
.B(n_396),
.Y(n_10224)
);

NAND2xp5_ASAP7_75t_SL g10225 ( 
.A(n_9632),
.B(n_1319),
.Y(n_10225)
);

A2O1A1Ixp33_ASAP7_75t_L g10226 ( 
.A1(n_9619),
.A2(n_1320),
.B(n_1321),
.C(n_1319),
.Y(n_10226)
);

INVx2_ASAP7_75t_L g10227 ( 
.A(n_9189),
.Y(n_10227)
);

OAI21xp5_ASAP7_75t_L g10228 ( 
.A1(n_9566),
.A2(n_397),
.B(n_398),
.Y(n_10228)
);

OAI21xp5_ASAP7_75t_L g10229 ( 
.A1(n_9416),
.A2(n_397),
.B(n_398),
.Y(n_10229)
);

OR2x6_ASAP7_75t_L g10230 ( 
.A(n_9372),
.B(n_1320),
.Y(n_10230)
);

NAND2xp5_ASAP7_75t_L g10231 ( 
.A(n_9194),
.B(n_1321),
.Y(n_10231)
);

OAI21x1_ASAP7_75t_L g10232 ( 
.A1(n_9226),
.A2(n_9196),
.B(n_9195),
.Y(n_10232)
);

AOI21x1_ASAP7_75t_L g10233 ( 
.A1(n_9186),
.A2(n_398),
.B(n_399),
.Y(n_10233)
);

NAND2xp5_ASAP7_75t_L g10234 ( 
.A(n_9199),
.B(n_1322),
.Y(n_10234)
);

NOR2xp33_ASAP7_75t_SL g10235 ( 
.A(n_9694),
.B(n_399),
.Y(n_10235)
);

OAI21x1_ASAP7_75t_L g10236 ( 
.A1(n_9276),
.A2(n_400),
.B(n_401),
.Y(n_10236)
);

NAND2xp5_ASAP7_75t_L g10237 ( 
.A(n_9124),
.B(n_9130),
.Y(n_10237)
);

OAI21x1_ASAP7_75t_L g10238 ( 
.A1(n_9548),
.A2(n_400),
.B(n_401),
.Y(n_10238)
);

OAI21x1_ASAP7_75t_L g10239 ( 
.A1(n_9131),
.A2(n_400),
.B(n_401),
.Y(n_10239)
);

AND2x4_ASAP7_75t_L g10240 ( 
.A(n_9490),
.B(n_1322),
.Y(n_10240)
);

OAI21x1_ASAP7_75t_L g10241 ( 
.A1(n_9146),
.A2(n_402),
.B(n_403),
.Y(n_10241)
);

NOR2xp33_ASAP7_75t_L g10242 ( 
.A(n_9641),
.B(n_1323),
.Y(n_10242)
);

O2A1O1Ixp5_ASAP7_75t_L g10243 ( 
.A1(n_9746),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_10243)
);

OAI21x1_ASAP7_75t_SL g10244 ( 
.A1(n_9629),
.A2(n_402),
.B(n_403),
.Y(n_10244)
);

AOI21xp5_ASAP7_75t_L g10245 ( 
.A1(n_9137),
.A2(n_404),
.B(n_405),
.Y(n_10245)
);

INVx5_ASAP7_75t_L g10246 ( 
.A(n_9372),
.Y(n_10246)
);

AOI21xp5_ASAP7_75t_L g10247 ( 
.A1(n_9365),
.A2(n_405),
.B(n_406),
.Y(n_10247)
);

OAI21x1_ASAP7_75t_L g10248 ( 
.A1(n_9228),
.A2(n_405),
.B(n_406),
.Y(n_10248)
);

NOR2xp33_ASAP7_75t_L g10249 ( 
.A(n_9115),
.B(n_1323),
.Y(n_10249)
);

AND2x2_ASAP7_75t_L g10250 ( 
.A(n_9375),
.B(n_1324),
.Y(n_10250)
);

AOI21xp5_ASAP7_75t_L g10251 ( 
.A1(n_9422),
.A2(n_406),
.B(n_407),
.Y(n_10251)
);

OAI22xp5_ASAP7_75t_L g10252 ( 
.A1(n_9511),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_10252)
);

BUFx6f_ASAP7_75t_L g10253 ( 
.A(n_9340),
.Y(n_10253)
);

NAND2xp5_ASAP7_75t_L g10254 ( 
.A(n_9230),
.B(n_1324),
.Y(n_10254)
);

OAI21x1_ASAP7_75t_L g10255 ( 
.A1(n_9234),
.A2(n_408),
.B(n_409),
.Y(n_10255)
);

AOI21xp5_ASAP7_75t_L g10256 ( 
.A1(n_9572),
.A2(n_410),
.B(n_411),
.Y(n_10256)
);

AOI21xp5_ASAP7_75t_SL g10257 ( 
.A1(n_9252),
.A2(n_9762),
.B(n_9518),
.Y(n_10257)
);

AOI21x1_ASAP7_75t_L g10258 ( 
.A1(n_9269),
.A2(n_410),
.B(n_411),
.Y(n_10258)
);

AOI21x1_ASAP7_75t_L g10259 ( 
.A1(n_9154),
.A2(n_411),
.B(n_412),
.Y(n_10259)
);

NAND2xp5_ASAP7_75t_L g10260 ( 
.A(n_9241),
.B(n_9248),
.Y(n_10260)
);

OR2x2_ASAP7_75t_L g10261 ( 
.A(n_9556),
.B(n_1325),
.Y(n_10261)
);

NAND2xp5_ASAP7_75t_L g10262 ( 
.A(n_9249),
.B(n_1325),
.Y(n_10262)
);

OAI21x1_ASAP7_75t_L g10263 ( 
.A1(n_9635),
.A2(n_412),
.B(n_413),
.Y(n_10263)
);

AOI21xp5_ASAP7_75t_L g10264 ( 
.A1(n_9483),
.A2(n_412),
.B(n_413),
.Y(n_10264)
);

AOI21x1_ASAP7_75t_L g10265 ( 
.A1(n_9159),
.A2(n_413),
.B(n_414),
.Y(n_10265)
);

AOI21xp5_ASAP7_75t_L g10266 ( 
.A1(n_9356),
.A2(n_414),
.B(n_415),
.Y(n_10266)
);

AOI221xp5_ASAP7_75t_L g10267 ( 
.A1(n_9613),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_10267)
);

NOR2xp33_ASAP7_75t_L g10268 ( 
.A(n_9120),
.B(n_1326),
.Y(n_10268)
);

AO31x2_ASAP7_75t_L g10269 ( 
.A1(n_9170),
.A2(n_417),
.A3(n_415),
.B(n_416),
.Y(n_10269)
);

AOI21xp5_ASAP7_75t_L g10270 ( 
.A1(n_9419),
.A2(n_416),
.B(n_418),
.Y(n_10270)
);

O2A1O1Ixp5_ASAP7_75t_L g10271 ( 
.A1(n_9634),
.A2(n_9431),
.B(n_9473),
.C(n_9415),
.Y(n_10271)
);

OAI22x1_ASAP7_75t_L g10272 ( 
.A1(n_9352),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_10272)
);

OAI22xp5_ASAP7_75t_L g10273 ( 
.A1(n_9430),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_10273)
);

AOI21xp5_ASAP7_75t_L g10274 ( 
.A1(n_9447),
.A2(n_419),
.B(n_420),
.Y(n_10274)
);

AOI21xp5_ASAP7_75t_L g10275 ( 
.A1(n_9478),
.A2(n_421),
.B(n_423),
.Y(n_10275)
);

CKINVDCx5p33_ASAP7_75t_R g10276 ( 
.A(n_9690),
.Y(n_10276)
);

AOI21xp5_ASAP7_75t_L g10277 ( 
.A1(n_9453),
.A2(n_421),
.B(n_423),
.Y(n_10277)
);

AND2x2_ASAP7_75t_L g10278 ( 
.A(n_9463),
.B(n_1326),
.Y(n_10278)
);

NOR2x1_ASAP7_75t_L g10279 ( 
.A(n_9486),
.B(n_1327),
.Y(n_10279)
);

OAI21xp5_ASAP7_75t_L g10280 ( 
.A1(n_9541),
.A2(n_421),
.B(n_423),
.Y(n_10280)
);

AOI21xp5_ASAP7_75t_L g10281 ( 
.A1(n_9454),
.A2(n_424),
.B(n_425),
.Y(n_10281)
);

OA22x2_ASAP7_75t_L g10282 ( 
.A1(n_9624),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_10282)
);

NOR2xp33_ASAP7_75t_L g10283 ( 
.A(n_9323),
.B(n_1328),
.Y(n_10283)
);

NAND2xp5_ASAP7_75t_L g10284 ( 
.A(n_9476),
.B(n_1328),
.Y(n_10284)
);

NAND2xp5_ASAP7_75t_L g10285 ( 
.A(n_9279),
.B(n_9517),
.Y(n_10285)
);

INVx2_ASAP7_75t_SL g10286 ( 
.A(n_9386),
.Y(n_10286)
);

BUFx6f_ASAP7_75t_L g10287 ( 
.A(n_9386),
.Y(n_10287)
);

NOR2xp67_ASAP7_75t_SL g10288 ( 
.A(n_9399),
.B(n_424),
.Y(n_10288)
);

OAI21x1_ASAP7_75t_L g10289 ( 
.A1(n_9637),
.A2(n_425),
.B(n_426),
.Y(n_10289)
);

AOI21x1_ASAP7_75t_L g10290 ( 
.A1(n_9393),
.A2(n_426),
.B(n_427),
.Y(n_10290)
);

INVx2_ASAP7_75t_L g10291 ( 
.A(n_9439),
.Y(n_10291)
);

HB1xp67_ASAP7_75t_L g10292 ( 
.A(n_9299),
.Y(n_10292)
);

NAND2xp5_ASAP7_75t_L g10293 ( 
.A(n_9616),
.B(n_1329),
.Y(n_10293)
);

AOI22xp33_ASAP7_75t_L g10294 ( 
.A1(n_9598),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_10294)
);

NAND2x1_ASAP7_75t_L g10295 ( 
.A(n_9514),
.B(n_1329),
.Y(n_10295)
);

AND2x2_ASAP7_75t_L g10296 ( 
.A(n_9474),
.B(n_1330),
.Y(n_10296)
);

NOR2xp33_ASAP7_75t_L g10297 ( 
.A(n_9376),
.B(n_1330),
.Y(n_10297)
);

AOI21xp5_ASAP7_75t_L g10298 ( 
.A1(n_9366),
.A2(n_428),
.B(n_429),
.Y(n_10298)
);

BUFx3_ASAP7_75t_L g10299 ( 
.A(n_9418),
.Y(n_10299)
);

A2O1A1Ixp33_ASAP7_75t_L g10300 ( 
.A1(n_9458),
.A2(n_1332),
.B(n_1333),
.C(n_1331),
.Y(n_10300)
);

OAI21x1_ASAP7_75t_L g10301 ( 
.A1(n_9424),
.A2(n_428),
.B(n_429),
.Y(n_10301)
);

NAND2xp5_ASAP7_75t_L g10302 ( 
.A(n_9522),
.B(n_1331),
.Y(n_10302)
);

NAND2xp5_ASAP7_75t_L g10303 ( 
.A(n_9535),
.B(n_1333),
.Y(n_10303)
);

OAI21x1_ASAP7_75t_L g10304 ( 
.A1(n_9524),
.A2(n_430),
.B(n_431),
.Y(n_10304)
);

AOI21xp5_ASAP7_75t_L g10305 ( 
.A1(n_9407),
.A2(n_9432),
.B(n_9492),
.Y(n_10305)
);

OAI21x1_ASAP7_75t_L g10306 ( 
.A1(n_9495),
.A2(n_430),
.B(n_431),
.Y(n_10306)
);

AND2x2_ASAP7_75t_L g10307 ( 
.A(n_9607),
.B(n_1334),
.Y(n_10307)
);

OAI21x1_ASAP7_75t_L g10308 ( 
.A1(n_9509),
.A2(n_430),
.B(n_431),
.Y(n_10308)
);

AND2x2_ASAP7_75t_L g10309 ( 
.A(n_9512),
.B(n_1334),
.Y(n_10309)
);

OAI21xp5_ASAP7_75t_L g10310 ( 
.A1(n_9501),
.A2(n_432),
.B(n_433),
.Y(n_10310)
);

AOI21xp5_ASAP7_75t_L g10311 ( 
.A1(n_9513),
.A2(n_432),
.B(n_433),
.Y(n_10311)
);

AO31x2_ASAP7_75t_L g10312 ( 
.A1(n_9369),
.A2(n_435),
.A3(n_432),
.B(n_434),
.Y(n_10312)
);

OAI21xp5_ASAP7_75t_L g10313 ( 
.A1(n_9598),
.A2(n_9534),
.B(n_9531),
.Y(n_10313)
);

INVx2_ASAP7_75t_L g10314 ( 
.A(n_9456),
.Y(n_10314)
);

AND2x2_ASAP7_75t_L g10315 ( 
.A(n_9273),
.B(n_1335),
.Y(n_10315)
);

INVxp67_ASAP7_75t_L g10316 ( 
.A(n_9160),
.Y(n_10316)
);

AOI21xp5_ASAP7_75t_L g10317 ( 
.A1(n_9536),
.A2(n_434),
.B(n_435),
.Y(n_10317)
);

AOI21xp5_ASAP7_75t_L g10318 ( 
.A1(n_9543),
.A2(n_9554),
.B(n_9520),
.Y(n_10318)
);

AOI21x1_ASAP7_75t_L g10319 ( 
.A1(n_9413),
.A2(n_435),
.B(n_436),
.Y(n_10319)
);

NAND2xp5_ASAP7_75t_L g10320 ( 
.A(n_9564),
.B(n_1335),
.Y(n_10320)
);

AND2x2_ASAP7_75t_L g10321 ( 
.A(n_9574),
.B(n_1336),
.Y(n_10321)
);

AO31x2_ASAP7_75t_L g10322 ( 
.A1(n_9558),
.A2(n_438),
.A3(n_436),
.B(n_437),
.Y(n_10322)
);

BUFx3_ASAP7_75t_L g10323 ( 
.A(n_9418),
.Y(n_10323)
);

AOI21xp5_ASAP7_75t_L g10324 ( 
.A1(n_9559),
.A2(n_9624),
.B(n_9604),
.Y(n_10324)
);

AOI21xp5_ASAP7_75t_L g10325 ( 
.A1(n_9135),
.A2(n_436),
.B(n_438),
.Y(n_10325)
);

AOI21xp5_ASAP7_75t_L g10326 ( 
.A1(n_9265),
.A2(n_439),
.B(n_440),
.Y(n_10326)
);

NAND2xp5_ASAP7_75t_L g10327 ( 
.A(n_9563),
.B(n_9573),
.Y(n_10327)
);

INVxp67_ASAP7_75t_L g10328 ( 
.A(n_9164),
.Y(n_10328)
);

INVx2_ASAP7_75t_L g10329 ( 
.A(n_9632),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_9309),
.Y(n_10330)
);

INVx2_ASAP7_75t_L g10331 ( 
.A(n_9329),
.Y(n_10331)
);

NOR2xp33_ASAP7_75t_L g10332 ( 
.A(n_9653),
.B(n_1336),
.Y(n_10332)
);

OA21x2_ASAP7_75t_L g10333 ( 
.A1(n_9620),
.A2(n_439),
.B(n_440),
.Y(n_10333)
);

NAND2xp33_ASAP7_75t_L g10334 ( 
.A(n_9598),
.B(n_439),
.Y(n_10334)
);

NAND2xp5_ASAP7_75t_L g10335 ( 
.A(n_9581),
.B(n_1337),
.Y(n_10335)
);

BUFx10_ASAP7_75t_L g10336 ( 
.A(n_9741),
.Y(n_10336)
);

INVxp67_ASAP7_75t_L g10337 ( 
.A(n_9387),
.Y(n_10337)
);

BUFx6f_ASAP7_75t_L g10338 ( 
.A(n_9494),
.Y(n_10338)
);

NAND2xp5_ASAP7_75t_L g10339 ( 
.A(n_9169),
.B(n_1337),
.Y(n_10339)
);

NAND2xp5_ASAP7_75t_L g10340 ( 
.A(n_9606),
.B(n_1338),
.Y(n_10340)
);

NAND2xp5_ASAP7_75t_L g10341 ( 
.A(n_9484),
.B(n_1338),
.Y(n_10341)
);

OAI22x1_ASAP7_75t_L g10342 ( 
.A1(n_9651),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_10342)
);

OAI21xp5_ASAP7_75t_L g10343 ( 
.A1(n_9654),
.A2(n_441),
.B(n_442),
.Y(n_10343)
);

AND3x4_ASAP7_75t_L g10344 ( 
.A(n_9674),
.B(n_441),
.C(n_443),
.Y(n_10344)
);

NAND2xp5_ASAP7_75t_L g10345 ( 
.A(n_9542),
.B(n_1339),
.Y(n_10345)
);

INVx2_ASAP7_75t_L g10346 ( 
.A(n_9494),
.Y(n_10346)
);

OAI21xp5_ASAP7_75t_L g10347 ( 
.A1(n_9646),
.A2(n_443),
.B(n_444),
.Y(n_10347)
);

NOR2xp33_ASAP7_75t_L g10348 ( 
.A(n_9623),
.B(n_1339),
.Y(n_10348)
);

NAND2x1_ASAP7_75t_L g10349 ( 
.A(n_9446),
.B(n_1340),
.Y(n_10349)
);

HB1xp67_ASAP7_75t_L g10350 ( 
.A(n_9459),
.Y(n_10350)
);

OAI22x1_ASAP7_75t_L g10351 ( 
.A1(n_9187),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_10351)
);

AOI21xp5_ASAP7_75t_SL g10352 ( 
.A1(n_9345),
.A2(n_1341),
.B(n_1340),
.Y(n_10352)
);

INVx3_ASAP7_75t_L g10353 ( 
.A(n_9438),
.Y(n_10353)
);

NAND2xp5_ASAP7_75t_L g10354 ( 
.A(n_9380),
.B(n_1341),
.Y(n_10354)
);

AOI21xp5_ASAP7_75t_SL g10355 ( 
.A1(n_9465),
.A2(n_1343),
.B(n_1342),
.Y(n_10355)
);

OAI21x1_ASAP7_75t_L g10356 ( 
.A1(n_9579),
.A2(n_444),
.B(n_445),
.Y(n_10356)
);

AOI21xp5_ASAP7_75t_L g10357 ( 
.A1(n_9761),
.A2(n_445),
.B(n_446),
.Y(n_10357)
);

NAND2xp5_ASAP7_75t_L g10358 ( 
.A(n_9383),
.B(n_1344),
.Y(n_10358)
);

INVxp67_ASAP7_75t_SL g10359 ( 
.A(n_9395),
.Y(n_10359)
);

AND2x2_ASAP7_75t_L g10360 ( 
.A(n_9485),
.B(n_9578),
.Y(n_10360)
);

A2O1A1Ixp33_ASAP7_75t_L g10361 ( 
.A1(n_9505),
.A2(n_1346),
.B(n_1347),
.C(n_1345),
.Y(n_10361)
);

OAI21xp5_ASAP7_75t_L g10362 ( 
.A1(n_9628),
.A2(n_446),
.B(n_447),
.Y(n_10362)
);

OAI21x1_ASAP7_75t_L g10363 ( 
.A1(n_9586),
.A2(n_446),
.B(n_447),
.Y(n_10363)
);

AO31x2_ASAP7_75t_L g10364 ( 
.A1(n_9645),
.A2(n_450),
.A3(n_448),
.B(n_449),
.Y(n_10364)
);

AO21x1_ASAP7_75t_L g10365 ( 
.A1(n_9335),
.A2(n_448),
.B(n_449),
.Y(n_10365)
);

INVx1_ASAP7_75t_L g10366 ( 
.A(n_9118),
.Y(n_10366)
);

INVx2_ASAP7_75t_L g10367 ( 
.A(n_9650),
.Y(n_10367)
);

NOR2x1_ASAP7_75t_SL g10368 ( 
.A(n_9639),
.B(n_1348),
.Y(n_10368)
);

AOI21xp5_ASAP7_75t_L g10369 ( 
.A1(n_9133),
.A2(n_9144),
.B(n_9540),
.Y(n_10369)
);

NAND2xp5_ASAP7_75t_L g10370 ( 
.A(n_9576),
.B(n_1349),
.Y(n_10370)
);

AOI22xp33_ASAP7_75t_L g10371 ( 
.A1(n_9640),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_10371)
);

OAI21xp5_ASAP7_75t_L g10372 ( 
.A1(n_9533),
.A2(n_450),
.B(n_451),
.Y(n_10372)
);

AOI21xp5_ASAP7_75t_L g10373 ( 
.A1(n_9118),
.A2(n_452),
.B(n_453),
.Y(n_10373)
);

INVx1_ASAP7_75t_L g10374 ( 
.A(n_9594),
.Y(n_10374)
);

CKINVDCx20_ASAP7_75t_R g10375 ( 
.A(n_9609),
.Y(n_10375)
);

NAND2xp5_ASAP7_75t_L g10376 ( 
.A(n_9636),
.B(n_1349),
.Y(n_10376)
);

NOR2xp33_ASAP7_75t_L g10377 ( 
.A(n_9871),
.B(n_9687),
.Y(n_10377)
);

OR2x6_ASAP7_75t_L g10378 ( 
.A(n_9874),
.B(n_9644),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_9894),
.Y(n_10379)
);

NAND3xp33_ASAP7_75t_SL g10380 ( 
.A(n_9785),
.B(n_9527),
.C(n_9630),
.Y(n_10380)
);

AOI21xp5_ASAP7_75t_L g10381 ( 
.A1(n_9859),
.A2(n_9893),
.B(n_9932),
.Y(n_10381)
);

AOI21xp5_ASAP7_75t_L g10382 ( 
.A1(n_10334),
.A2(n_452),
.B(n_453),
.Y(n_10382)
);

OAI21x1_ASAP7_75t_L g10383 ( 
.A1(n_9852),
.A2(n_452),
.B(n_453),
.Y(n_10383)
);

OAI21x1_ASAP7_75t_L g10384 ( 
.A1(n_9997),
.A2(n_454),
.B(n_455),
.Y(n_10384)
);

NAND3xp33_ASAP7_75t_L g10385 ( 
.A(n_10005),
.B(n_454),
.C(n_455),
.Y(n_10385)
);

INVx1_ASAP7_75t_L g10386 ( 
.A(n_9895),
.Y(n_10386)
);

NAND3xp33_ASAP7_75t_L g10387 ( 
.A(n_10040),
.B(n_454),
.C(n_456),
.Y(n_10387)
);

BUFx12f_ASAP7_75t_L g10388 ( 
.A(n_9844),
.Y(n_10388)
);

OAI22xp5_ASAP7_75t_L g10389 ( 
.A1(n_10037),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_10389)
);

AO31x2_ASAP7_75t_L g10390 ( 
.A1(n_10012),
.A2(n_459),
.A3(n_456),
.B(n_458),
.Y(n_10390)
);

OAI21xp5_ASAP7_75t_L g10391 ( 
.A1(n_9978),
.A2(n_458),
.B(n_459),
.Y(n_10391)
);

OAI21xp5_ASAP7_75t_L g10392 ( 
.A1(n_9812),
.A2(n_459),
.B(n_460),
.Y(n_10392)
);

OAI21xp5_ASAP7_75t_L g10393 ( 
.A1(n_9779),
.A2(n_460),
.B(n_461),
.Y(n_10393)
);

OAI21x1_ASAP7_75t_SL g10394 ( 
.A1(n_10373),
.A2(n_460),
.B(n_461),
.Y(n_10394)
);

INVx2_ASAP7_75t_L g10395 ( 
.A(n_9818),
.Y(n_10395)
);

AOI21xp5_ASAP7_75t_L g10396 ( 
.A1(n_10182),
.A2(n_461),
.B(n_462),
.Y(n_10396)
);

AOI21xp5_ASAP7_75t_L g10397 ( 
.A1(n_9805),
.A2(n_462),
.B(n_463),
.Y(n_10397)
);

AO21x1_ASAP7_75t_L g10398 ( 
.A1(n_9877),
.A2(n_462),
.B(n_463),
.Y(n_10398)
);

NOR2xp67_ASAP7_75t_L g10399 ( 
.A(n_9784),
.B(n_463),
.Y(n_10399)
);

OAI21xp5_ASAP7_75t_L g10400 ( 
.A1(n_9918),
.A2(n_464),
.B(n_465),
.Y(n_10400)
);

AOI21xp5_ASAP7_75t_L g10401 ( 
.A1(n_10165),
.A2(n_464),
.B(n_465),
.Y(n_10401)
);

AOI21xp5_ASAP7_75t_L g10402 ( 
.A1(n_10007),
.A2(n_464),
.B(n_466),
.Y(n_10402)
);

NAND2xp5_ASAP7_75t_L g10403 ( 
.A(n_9803),
.B(n_1351),
.Y(n_10403)
);

AOI21xp5_ASAP7_75t_L g10404 ( 
.A1(n_10202),
.A2(n_466),
.B(n_467),
.Y(n_10404)
);

OAI21xp5_ASAP7_75t_L g10405 ( 
.A1(n_10213),
.A2(n_467),
.B(n_468),
.Y(n_10405)
);

INVx1_ASAP7_75t_L g10406 ( 
.A(n_9928),
.Y(n_10406)
);

AOI21x1_ASAP7_75t_L g10407 ( 
.A1(n_9776),
.A2(n_468),
.B(n_469),
.Y(n_10407)
);

A2O1A1Ixp33_ASAP7_75t_L g10408 ( 
.A1(n_9836),
.A2(n_9801),
.B(n_10124),
.C(n_10168),
.Y(n_10408)
);

NAND2xp5_ASAP7_75t_L g10409 ( 
.A(n_9839),
.B(n_1351),
.Y(n_10409)
);

AOI21xp5_ASAP7_75t_L g10410 ( 
.A1(n_10257),
.A2(n_468),
.B(n_469),
.Y(n_10410)
);

AOI21xp5_ASAP7_75t_L g10411 ( 
.A1(n_9961),
.A2(n_470),
.B(n_471),
.Y(n_10411)
);

NOR2x1_ASAP7_75t_L g10412 ( 
.A(n_10014),
.B(n_470),
.Y(n_10412)
);

AOI21xp5_ASAP7_75t_L g10413 ( 
.A1(n_9815),
.A2(n_470),
.B(n_471),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_9930),
.Y(n_10414)
);

OA21x2_ASAP7_75t_L g10415 ( 
.A1(n_9782),
.A2(n_1354),
.B(n_1353),
.Y(n_10415)
);

BUFx4_ASAP7_75t_SL g10416 ( 
.A(n_10375),
.Y(n_10416)
);

INVx1_ASAP7_75t_L g10417 ( 
.A(n_9850),
.Y(n_10417)
);

OAI21xp5_ASAP7_75t_L g10418 ( 
.A1(n_9791),
.A2(n_471),
.B(n_472),
.Y(n_10418)
);

NAND2xp5_ASAP7_75t_L g10419 ( 
.A(n_9949),
.B(n_1355),
.Y(n_10419)
);

INVx1_ASAP7_75t_L g10420 ( 
.A(n_9858),
.Y(n_10420)
);

OR2x2_ASAP7_75t_L g10421 ( 
.A(n_9786),
.B(n_1355),
.Y(n_10421)
);

NAND2xp5_ASAP7_75t_L g10422 ( 
.A(n_9842),
.B(n_1356),
.Y(n_10422)
);

INVx1_ASAP7_75t_L g10423 ( 
.A(n_9863),
.Y(n_10423)
);

OAI21xp5_ASAP7_75t_L g10424 ( 
.A1(n_9828),
.A2(n_473),
.B(n_474),
.Y(n_10424)
);

INVx1_ASAP7_75t_L g10425 ( 
.A(n_9872),
.Y(n_10425)
);

BUFx6f_ASAP7_75t_L g10426 ( 
.A(n_10160),
.Y(n_10426)
);

NAND3xp33_ASAP7_75t_L g10427 ( 
.A(n_9879),
.B(n_473),
.C(n_474),
.Y(n_10427)
);

OAI21x1_ASAP7_75t_L g10428 ( 
.A1(n_10125),
.A2(n_474),
.B(n_475),
.Y(n_10428)
);

INVx1_ASAP7_75t_L g10429 ( 
.A(n_9881),
.Y(n_10429)
);

NOR2x1_ASAP7_75t_SL g10430 ( 
.A(n_9799),
.B(n_1356),
.Y(n_10430)
);

NAND2xp5_ASAP7_75t_L g10431 ( 
.A(n_9960),
.B(n_1357),
.Y(n_10431)
);

OAI21x1_ASAP7_75t_L g10432 ( 
.A1(n_10173),
.A2(n_475),
.B(n_476),
.Y(n_10432)
);

BUFx2_ASAP7_75t_L g10433 ( 
.A(n_10091),
.Y(n_10433)
);

OAI21x1_ASAP7_75t_L g10434 ( 
.A1(n_9927),
.A2(n_475),
.B(n_476),
.Y(n_10434)
);

OAI21x1_ASAP7_75t_L g10435 ( 
.A1(n_9795),
.A2(n_476),
.B(n_477),
.Y(n_10435)
);

OAI21x1_ASAP7_75t_L g10436 ( 
.A1(n_9778),
.A2(n_9804),
.B(n_10215),
.Y(n_10436)
);

OAI22xp5_ASAP7_75t_L g10437 ( 
.A1(n_10185),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_10437)
);

AO31x2_ASAP7_75t_L g10438 ( 
.A1(n_9919),
.A2(n_481),
.A3(n_478),
.B(n_480),
.Y(n_10438)
);

INVx3_ASAP7_75t_L g10439 ( 
.A(n_9820),
.Y(n_10439)
);

AND2x4_ASAP7_75t_SL g10440 ( 
.A(n_10079),
.B(n_1357),
.Y(n_10440)
);

OAI22xp5_ASAP7_75t_L g10441 ( 
.A1(n_9905),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_10441)
);

NAND2xp5_ASAP7_75t_L g10442 ( 
.A(n_9807),
.B(n_1358),
.Y(n_10442)
);

AOI21xp5_ASAP7_75t_L g10443 ( 
.A1(n_9817),
.A2(n_481),
.B(n_482),
.Y(n_10443)
);

AOI22xp5_ASAP7_75t_L g10444 ( 
.A1(n_9984),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_10444)
);

NAND2xp5_ASAP7_75t_L g10445 ( 
.A(n_10292),
.B(n_1359),
.Y(n_10445)
);

INVx2_ASAP7_75t_SL g10446 ( 
.A(n_9908),
.Y(n_10446)
);

AND2x2_ASAP7_75t_L g10447 ( 
.A(n_9783),
.B(n_1359),
.Y(n_10447)
);

OAI21x1_ASAP7_75t_L g10448 ( 
.A1(n_10207),
.A2(n_483),
.B(n_484),
.Y(n_10448)
);

NAND2xp5_ASAP7_75t_L g10449 ( 
.A(n_9830),
.B(n_1360),
.Y(n_10449)
);

OAI21x1_ASAP7_75t_L g10450 ( 
.A1(n_10232),
.A2(n_9887),
.B(n_9883),
.Y(n_10450)
);

INVx1_ASAP7_75t_L g10451 ( 
.A(n_9923),
.Y(n_10451)
);

AOI21xp5_ASAP7_75t_L g10452 ( 
.A1(n_9825),
.A2(n_484),
.B(n_485),
.Y(n_10452)
);

AOI22xp5_ASAP7_75t_L g10453 ( 
.A1(n_10024),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_10453)
);

NAND2xp5_ASAP7_75t_L g10454 ( 
.A(n_9832),
.B(n_1360),
.Y(n_10454)
);

OA21x2_ASAP7_75t_L g10455 ( 
.A1(n_9870),
.A2(n_1362),
.B(n_1361),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_9925),
.Y(n_10456)
);

INVx2_ASAP7_75t_L g10457 ( 
.A(n_9945),
.Y(n_10457)
);

NAND3xp33_ASAP7_75t_L g10458 ( 
.A(n_9819),
.B(n_486),
.C(n_487),
.Y(n_10458)
);

AOI21xp5_ASAP7_75t_L g10459 ( 
.A1(n_9846),
.A2(n_486),
.B(n_487),
.Y(n_10459)
);

AOI21xp5_ASAP7_75t_L g10460 ( 
.A1(n_10158),
.A2(n_488),
.B(n_489),
.Y(n_10460)
);

BUFx4f_ASAP7_75t_L g10461 ( 
.A(n_10253),
.Y(n_10461)
);

INVx1_ASAP7_75t_L g10462 ( 
.A(n_9856),
.Y(n_10462)
);

OAI22xp5_ASAP7_75t_L g10463 ( 
.A1(n_9806),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_10463)
);

AOI21xp5_ASAP7_75t_L g10464 ( 
.A1(n_9876),
.A2(n_490),
.B(n_491),
.Y(n_10464)
);

AOI211x1_ASAP7_75t_L g10465 ( 
.A1(n_10365),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_10465)
);

INVx3_ASAP7_75t_L g10466 ( 
.A(n_10200),
.Y(n_10466)
);

INVx1_ASAP7_75t_L g10467 ( 
.A(n_9946),
.Y(n_10467)
);

NAND2xp5_ASAP7_75t_L g10468 ( 
.A(n_10367),
.B(n_1361),
.Y(n_10468)
);

NOR2xp67_ASAP7_75t_L g10469 ( 
.A(n_9799),
.B(n_491),
.Y(n_10469)
);

BUFx3_ASAP7_75t_L g10470 ( 
.A(n_10253),
.Y(n_10470)
);

NAND2xp5_ASAP7_75t_SL g10471 ( 
.A(n_9992),
.B(n_1362),
.Y(n_10471)
);

OAI21x1_ASAP7_75t_SL g10472 ( 
.A1(n_9829),
.A2(n_9890),
.B(n_9955),
.Y(n_10472)
);

OAI21x1_ASAP7_75t_L g10473 ( 
.A1(n_9902),
.A2(n_9915),
.B(n_9904),
.Y(n_10473)
);

AOI21xp5_ASAP7_75t_SL g10474 ( 
.A1(n_9929),
.A2(n_492),
.B(n_493),
.Y(n_10474)
);

BUFx3_ASAP7_75t_L g10475 ( 
.A(n_10287),
.Y(n_10475)
);

NAND2xp5_ASAP7_75t_L g10476 ( 
.A(n_10218),
.B(n_1363),
.Y(n_10476)
);

OAI21xp5_ASAP7_75t_L g10477 ( 
.A1(n_9837),
.A2(n_492),
.B(n_493),
.Y(n_10477)
);

AOI21xp5_ASAP7_75t_L g10478 ( 
.A1(n_10123),
.A2(n_493),
.B(n_494),
.Y(n_10478)
);

NAND2xp5_ASAP7_75t_L g10479 ( 
.A(n_10180),
.B(n_1363),
.Y(n_10479)
);

NAND2xp5_ASAP7_75t_L g10480 ( 
.A(n_10194),
.B(n_1364),
.Y(n_10480)
);

NAND2xp5_ASAP7_75t_L g10481 ( 
.A(n_10209),
.B(n_1364),
.Y(n_10481)
);

INVx4_ASAP7_75t_L g10482 ( 
.A(n_10287),
.Y(n_10482)
);

OAI22xp5_ASAP7_75t_L g10483 ( 
.A1(n_10294),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_10483)
);

AOI221xp5_ASAP7_75t_SL g10484 ( 
.A1(n_10325),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.C(n_497),
.Y(n_10484)
);

OAI21xp5_ASAP7_75t_L g10485 ( 
.A1(n_9860),
.A2(n_495),
.B(n_496),
.Y(n_10485)
);

OAI21x1_ASAP7_75t_L g10486 ( 
.A1(n_10035),
.A2(n_497),
.B(n_498),
.Y(n_10486)
);

OAI21x1_ASAP7_75t_L g10487 ( 
.A1(n_9813),
.A2(n_497),
.B(n_498),
.Y(n_10487)
);

AOI21x1_ASAP7_75t_SL g10488 ( 
.A1(n_10206),
.A2(n_10000),
.B(n_9991),
.Y(n_10488)
);

AND2x6_ASAP7_75t_SL g10489 ( 
.A(n_10297),
.B(n_498),
.Y(n_10489)
);

NAND2xp5_ASAP7_75t_L g10490 ( 
.A(n_10227),
.B(n_1365),
.Y(n_10490)
);

AOI21xp5_ASAP7_75t_L g10491 ( 
.A1(n_10171),
.A2(n_499),
.B(n_500),
.Y(n_10491)
);

A2O1A1Ixp33_ASAP7_75t_L g10492 ( 
.A1(n_9979),
.A2(n_1366),
.B(n_1367),
.C(n_1365),
.Y(n_10492)
);

O2A1O1Ixp33_ASAP7_75t_L g10493 ( 
.A1(n_9811),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_10493)
);

AOI21xp5_ASAP7_75t_L g10494 ( 
.A1(n_9966),
.A2(n_500),
.B(n_501),
.Y(n_10494)
);

INVx1_ASAP7_75t_L g10495 ( 
.A(n_9952),
.Y(n_10495)
);

AO31x2_ASAP7_75t_L g10496 ( 
.A1(n_9920),
.A2(n_503),
.A3(n_501),
.B(n_502),
.Y(n_10496)
);

INVx1_ASAP7_75t_L g10497 ( 
.A(n_9802),
.Y(n_10497)
);

OAI21x1_ASAP7_75t_L g10498 ( 
.A1(n_9808),
.A2(n_502),
.B(n_503),
.Y(n_10498)
);

OAI21xp5_ASAP7_75t_L g10499 ( 
.A1(n_9873),
.A2(n_502),
.B(n_504),
.Y(n_10499)
);

AOI21xp5_ASAP7_75t_L g10500 ( 
.A1(n_9980),
.A2(n_504),
.B(n_505),
.Y(n_10500)
);

OAI21xp5_ASAP7_75t_L g10501 ( 
.A1(n_9878),
.A2(n_504),
.B(n_505),
.Y(n_10501)
);

AOI21xp5_ASAP7_75t_L g10502 ( 
.A1(n_10019),
.A2(n_506),
.B(n_507),
.Y(n_10502)
);

OAI21xp33_ASAP7_75t_L g10503 ( 
.A1(n_10300),
.A2(n_506),
.B(n_507),
.Y(n_10503)
);

INVx1_ASAP7_75t_L g10504 ( 
.A(n_9947),
.Y(n_10504)
);

INVx1_ASAP7_75t_L g10505 ( 
.A(n_9975),
.Y(n_10505)
);

NOR2xp33_ASAP7_75t_L g10506 ( 
.A(n_10285),
.B(n_1370),
.Y(n_10506)
);

NOR2xp33_ASAP7_75t_L g10507 ( 
.A(n_10017),
.B(n_9824),
.Y(n_10507)
);

NAND2xp5_ASAP7_75t_L g10508 ( 
.A(n_10018),
.B(n_1370),
.Y(n_10508)
);

NAND2x1p5_ASAP7_75t_L g10509 ( 
.A(n_9962),
.B(n_1372),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9910),
.Y(n_10510)
);

OA21x2_ASAP7_75t_L g10511 ( 
.A1(n_9917),
.A2(n_1373),
.B(n_1372),
.Y(n_10511)
);

A2O1A1Ixp33_ASAP7_75t_L g10512 ( 
.A1(n_9922),
.A2(n_1374),
.B(n_1375),
.C(n_1373),
.Y(n_10512)
);

A2O1A1Ixp33_ASAP7_75t_L g10513 ( 
.A1(n_9951),
.A2(n_1375),
.B(n_1376),
.C(n_1374),
.Y(n_10513)
);

OR2x2_ASAP7_75t_L g10514 ( 
.A(n_10043),
.B(n_10291),
.Y(n_10514)
);

NAND2xp5_ASAP7_75t_L g10515 ( 
.A(n_10071),
.B(n_1376),
.Y(n_10515)
);

AOI21xp5_ASAP7_75t_L g10516 ( 
.A1(n_9822),
.A2(n_9831),
.B(n_9823),
.Y(n_10516)
);

INVx2_ASAP7_75t_L g10517 ( 
.A(n_10139),
.Y(n_10517)
);

OAI21x1_ASAP7_75t_L g10518 ( 
.A1(n_9834),
.A2(n_506),
.B(n_507),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_L g10519 ( 
.A(n_10075),
.B(n_1377),
.Y(n_10519)
);

INVx2_ASAP7_75t_L g10520 ( 
.A(n_10113),
.Y(n_10520)
);

INVx3_ASAP7_75t_L g10521 ( 
.A(n_9809),
.Y(n_10521)
);

A2O1A1Ixp33_ASAP7_75t_L g10522 ( 
.A1(n_9959),
.A2(n_1378),
.B(n_1379),
.C(n_1377),
.Y(n_10522)
);

OAI21x1_ASAP7_75t_L g10523 ( 
.A1(n_9835),
.A2(n_508),
.B(n_509),
.Y(n_10523)
);

AOI21xp5_ASAP7_75t_L g10524 ( 
.A1(n_9983),
.A2(n_508),
.B(n_509),
.Y(n_10524)
);

AOI21xp5_ASAP7_75t_L g10525 ( 
.A1(n_10083),
.A2(n_508),
.B(n_509),
.Y(n_10525)
);

INVxp67_ASAP7_75t_L g10526 ( 
.A(n_9869),
.Y(n_10526)
);

AOI31xp67_ASAP7_75t_L g10527 ( 
.A1(n_9898),
.A2(n_512),
.A3(n_510),
.B(n_511),
.Y(n_10527)
);

INVx2_ASAP7_75t_L g10528 ( 
.A(n_10128),
.Y(n_10528)
);

AOI21xp5_ASAP7_75t_L g10529 ( 
.A1(n_10198),
.A2(n_510),
.B(n_512),
.Y(n_10529)
);

INVx1_ASAP7_75t_L g10530 ( 
.A(n_9985),
.Y(n_10530)
);

AND2x4_ASAP7_75t_L g10531 ( 
.A(n_9993),
.B(n_1378),
.Y(n_10531)
);

OAI21x1_ASAP7_75t_L g10532 ( 
.A1(n_9841),
.A2(n_512),
.B(n_513),
.Y(n_10532)
);

A2O1A1Ixp33_ASAP7_75t_L g10533 ( 
.A1(n_10221),
.A2(n_1380),
.B(n_1381),
.C(n_1379),
.Y(n_10533)
);

INVx2_ASAP7_75t_SL g10534 ( 
.A(n_10064),
.Y(n_10534)
);

OA21x2_ASAP7_75t_L g10535 ( 
.A1(n_10239),
.A2(n_1381),
.B(n_1380),
.Y(n_10535)
);

NOR2xp33_ASAP7_75t_L g10536 ( 
.A(n_9855),
.B(n_1382),
.Y(n_10536)
);

NAND2xp5_ASAP7_75t_L g10537 ( 
.A(n_10129),
.B(n_1382),
.Y(n_10537)
);

INVx3_ASAP7_75t_SL g10538 ( 
.A(n_9845),
.Y(n_10538)
);

NAND2xp5_ASAP7_75t_L g10539 ( 
.A(n_10155),
.B(n_10184),
.Y(n_10539)
);

A2O1A1Ixp33_ASAP7_75t_L g10540 ( 
.A1(n_10271),
.A2(n_1384),
.B(n_1385),
.C(n_1383),
.Y(n_10540)
);

NAND2xp5_ASAP7_75t_L g10541 ( 
.A(n_10314),
.B(n_1383),
.Y(n_10541)
);

NAND2xp5_ASAP7_75t_SL g10542 ( 
.A(n_9992),
.B(n_1386),
.Y(n_10542)
);

OAI21x1_ASAP7_75t_L g10543 ( 
.A1(n_9848),
.A2(n_513),
.B(n_514),
.Y(n_10543)
);

NAND2xp5_ASAP7_75t_L g10544 ( 
.A(n_10331),
.B(n_1386),
.Y(n_10544)
);

NAND2xp5_ASAP7_75t_L g10545 ( 
.A(n_10337),
.B(n_1387),
.Y(n_10545)
);

OAI21x1_ASAP7_75t_L g10546 ( 
.A1(n_9849),
.A2(n_513),
.B(n_514),
.Y(n_10546)
);

AOI31xp67_ASAP7_75t_L g10547 ( 
.A1(n_9840),
.A2(n_516),
.A3(n_514),
.B(n_515),
.Y(n_10547)
);

OAI21xp5_ASAP7_75t_L g10548 ( 
.A1(n_10067),
.A2(n_515),
.B(n_516),
.Y(n_10548)
);

NAND2xp5_ASAP7_75t_L g10549 ( 
.A(n_10330),
.B(n_1387),
.Y(n_10549)
);

OAI22xp5_ASAP7_75t_L g10550 ( 
.A1(n_10222),
.A2(n_9847),
.B1(n_9780),
.B2(n_9865),
.Y(n_10550)
);

OAI21x1_ASAP7_75t_SL g10551 ( 
.A1(n_10134),
.A2(n_515),
.B(n_517),
.Y(n_10551)
);

AND2x2_ASAP7_75t_L g10552 ( 
.A(n_10028),
.B(n_1389),
.Y(n_10552)
);

NAND2xp5_ASAP7_75t_SL g10553 ( 
.A(n_9992),
.B(n_1390),
.Y(n_10553)
);

O2A1O1Ixp5_ASAP7_75t_SL g10554 ( 
.A1(n_9958),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_10554)
);

NAND2xp5_ASAP7_75t_L g10555 ( 
.A(n_9995),
.B(n_1390),
.Y(n_10555)
);

AND2x2_ASAP7_75t_L g10556 ( 
.A(n_10098),
.B(n_1391),
.Y(n_10556)
);

INVx3_ASAP7_75t_L g10557 ( 
.A(n_9809),
.Y(n_10557)
);

OAI21x1_ASAP7_75t_L g10558 ( 
.A1(n_9861),
.A2(n_518),
.B(n_519),
.Y(n_10558)
);

AO32x2_ASAP7_75t_L g10559 ( 
.A1(n_9796),
.A2(n_10104),
.A3(n_10252),
.B1(n_9969),
.B2(n_10066),
.Y(n_10559)
);

INVx2_ASAP7_75t_SL g10560 ( 
.A(n_9857),
.Y(n_10560)
);

OAI22xp5_ASAP7_75t_L g10561 ( 
.A1(n_10246),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_10561)
);

OAI21x1_ASAP7_75t_L g10562 ( 
.A1(n_9868),
.A2(n_520),
.B(n_521),
.Y(n_10562)
);

AND2x2_ASAP7_75t_L g10563 ( 
.A(n_9875),
.B(n_1391),
.Y(n_10563)
);

INVx1_ASAP7_75t_L g10564 ( 
.A(n_9885),
.Y(n_10564)
);

NOR2xp33_ASAP7_75t_L g10565 ( 
.A(n_10327),
.B(n_1392),
.Y(n_10565)
);

INVxp67_ASAP7_75t_L g10566 ( 
.A(n_10350),
.Y(n_10566)
);

OAI22xp5_ASAP7_75t_L g10567 ( 
.A1(n_10246),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_10567)
);

INVx2_ASAP7_75t_L g10568 ( 
.A(n_9798),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_9906),
.Y(n_10569)
);

AOI21xp5_ASAP7_75t_L g10570 ( 
.A1(n_10065),
.A2(n_521),
.B(n_522),
.Y(n_10570)
);

AOI21x1_ASAP7_75t_L g10571 ( 
.A1(n_9891),
.A2(n_522),
.B(n_523),
.Y(n_10571)
);

OAI21xp5_ASAP7_75t_L g10572 ( 
.A1(n_10117),
.A2(n_523),
.B(n_524),
.Y(n_10572)
);

INVx2_ASAP7_75t_L g10573 ( 
.A(n_9790),
.Y(n_10573)
);

AND2x2_ASAP7_75t_L g10574 ( 
.A(n_10100),
.B(n_1392),
.Y(n_10574)
);

AO31x2_ASAP7_75t_L g10575 ( 
.A1(n_9971),
.A2(n_526),
.A3(n_524),
.B(n_525),
.Y(n_10575)
);

NAND3xp33_ASAP7_75t_SL g10576 ( 
.A(n_10372),
.B(n_524),
.C(n_526),
.Y(n_10576)
);

AOI21xp5_ASAP7_75t_L g10577 ( 
.A1(n_10070),
.A2(n_526),
.B(n_527),
.Y(n_10577)
);

OAI21x1_ASAP7_75t_L g10578 ( 
.A1(n_9981),
.A2(n_527),
.B(n_528),
.Y(n_10578)
);

NOR2xp33_ASAP7_75t_L g10579 ( 
.A(n_10237),
.B(n_1393),
.Y(n_10579)
);

BUFx8_ASAP7_75t_SL g10580 ( 
.A(n_10276),
.Y(n_10580)
);

AOI21xp5_ASAP7_75t_L g10581 ( 
.A1(n_10072),
.A2(n_527),
.B(n_528),
.Y(n_10581)
);

AND2x2_ASAP7_75t_L g10582 ( 
.A(n_10360),
.B(n_10190),
.Y(n_10582)
);

AOI22xp5_ASAP7_75t_L g10583 ( 
.A1(n_9862),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_10583)
);

BUFx2_ASAP7_75t_L g10584 ( 
.A(n_10089),
.Y(n_10584)
);

NAND3x1_ASAP7_75t_L g10585 ( 
.A(n_10249),
.B(n_529),
.C(n_530),
.Y(n_10585)
);

AOI21xp5_ASAP7_75t_L g10586 ( 
.A1(n_10196),
.A2(n_529),
.B(n_530),
.Y(n_10586)
);

AOI21xp5_ASAP7_75t_L g10587 ( 
.A1(n_10164),
.A2(n_531),
.B(n_532),
.Y(n_10587)
);

AND2x4_ASAP7_75t_L g10588 ( 
.A(n_10096),
.B(n_1393),
.Y(n_10588)
);

O2A1O1Ixp5_ASAP7_75t_L g10589 ( 
.A1(n_9998),
.A2(n_533),
.B(n_531),
.C(n_532),
.Y(n_10589)
);

AOI22x1_ASAP7_75t_L g10590 ( 
.A1(n_10061),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_10590)
);

OAI21xp5_ASAP7_75t_L g10591 ( 
.A1(n_10118),
.A2(n_533),
.B(n_534),
.Y(n_10591)
);

CKINVDCx20_ASAP7_75t_R g10592 ( 
.A(n_9963),
.Y(n_10592)
);

AOI221x1_ASAP7_75t_L g10593 ( 
.A1(n_10172),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.C(n_537),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_10322),
.Y(n_10594)
);

O2A1O1Ixp5_ASAP7_75t_L g10595 ( 
.A1(n_10203),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_10595)
);

OAI21x1_ASAP7_75t_L g10596 ( 
.A1(n_9986),
.A2(n_535),
.B(n_536),
.Y(n_10596)
);

AO31x2_ASAP7_75t_L g10597 ( 
.A1(n_10036),
.A2(n_539),
.A3(n_537),
.B(n_538),
.Y(n_10597)
);

NAND2xp5_ASAP7_75t_L g10598 ( 
.A(n_10318),
.B(n_1394),
.Y(n_10598)
);

NAND2xp33_ASAP7_75t_R g10599 ( 
.A(n_10025),
.B(n_538),
.Y(n_10599)
);

OAI21x1_ASAP7_75t_SL g10600 ( 
.A1(n_10204),
.A2(n_538),
.B(n_539),
.Y(n_10600)
);

INVx2_ASAP7_75t_L g10601 ( 
.A(n_9787),
.Y(n_10601)
);

OAI21x1_ASAP7_75t_L g10602 ( 
.A1(n_10001),
.A2(n_539),
.B(n_540),
.Y(n_10602)
);

NAND3x1_ASAP7_75t_L g10603 ( 
.A(n_10268),
.B(n_540),
.C(n_541),
.Y(n_10603)
);

AO21x1_ASAP7_75t_L g10604 ( 
.A1(n_10366),
.A2(n_540),
.B(n_541),
.Y(n_10604)
);

INVx1_ASAP7_75t_SL g10605 ( 
.A(n_9833),
.Y(n_10605)
);

OAI21x1_ASAP7_75t_L g10606 ( 
.A1(n_10003),
.A2(n_541),
.B(n_542),
.Y(n_10606)
);

AOI21xp5_ASAP7_75t_L g10607 ( 
.A1(n_10154),
.A2(n_542),
.B(n_543),
.Y(n_10607)
);

NAND2xp5_ASAP7_75t_SL g10608 ( 
.A(n_9992),
.B(n_1394),
.Y(n_10608)
);

AOI21xp5_ASAP7_75t_L g10609 ( 
.A1(n_10135),
.A2(n_542),
.B(n_543),
.Y(n_10609)
);

INVxp67_ASAP7_75t_L g10610 ( 
.A(n_10110),
.Y(n_10610)
);

AOI21xp5_ASAP7_75t_L g10611 ( 
.A1(n_10034),
.A2(n_543),
.B(n_544),
.Y(n_10611)
);

AO21x1_ASAP7_75t_L g10612 ( 
.A1(n_10247),
.A2(n_544),
.B(n_545),
.Y(n_10612)
);

INVx1_ASAP7_75t_L g10613 ( 
.A(n_10322),
.Y(n_10613)
);

BUFx3_ASAP7_75t_L g10614 ( 
.A(n_10338),
.Y(n_10614)
);

BUFx2_ASAP7_75t_L g10615 ( 
.A(n_10120),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_9886),
.Y(n_10616)
);

INVx1_ASAP7_75t_L g10617 ( 
.A(n_9889),
.Y(n_10617)
);

AOI21xp5_ASAP7_75t_SL g10618 ( 
.A1(n_10103),
.A2(n_544),
.B(n_545),
.Y(n_10618)
);

NAND2xp33_ASAP7_75t_L g10619 ( 
.A(n_10033),
.B(n_546),
.Y(n_10619)
);

OAI21x1_ASAP7_75t_L g10620 ( 
.A1(n_10006),
.A2(n_546),
.B(n_547),
.Y(n_10620)
);

OAI21x1_ASAP7_75t_L g10621 ( 
.A1(n_10008),
.A2(n_546),
.B(n_548),
.Y(n_10621)
);

AND2x4_ASAP7_75t_L g10622 ( 
.A(n_9907),
.B(n_1395),
.Y(n_10622)
);

NAND2xp5_ASAP7_75t_L g10623 ( 
.A(n_10260),
.B(n_10313),
.Y(n_10623)
);

A2O1A1Ixp33_ASAP7_75t_L g10624 ( 
.A1(n_10228),
.A2(n_10010),
.B(n_10009),
.C(n_10186),
.Y(n_10624)
);

OAI21x1_ASAP7_75t_L g10625 ( 
.A1(n_10027),
.A2(n_548),
.B(n_549),
.Y(n_10625)
);

AO21x1_ASAP7_75t_L g10626 ( 
.A1(n_10251),
.A2(n_10256),
.B(n_9821),
.Y(n_10626)
);

OR2x2_ASAP7_75t_L g10627 ( 
.A(n_9854),
.B(n_10374),
.Y(n_10627)
);

AOI21x1_ASAP7_75t_L g10628 ( 
.A1(n_10290),
.A2(n_548),
.B(n_549),
.Y(n_10628)
);

AOI21xp5_ASAP7_75t_L g10629 ( 
.A1(n_10026),
.A2(n_549),
.B(n_550),
.Y(n_10629)
);

AOI21xp5_ASAP7_75t_L g10630 ( 
.A1(n_10094),
.A2(n_10122),
.B(n_9867),
.Y(n_10630)
);

OAI21x1_ASAP7_75t_L g10631 ( 
.A1(n_10032),
.A2(n_550),
.B(n_551),
.Y(n_10631)
);

OAI21x1_ASAP7_75t_L g10632 ( 
.A1(n_10049),
.A2(n_550),
.B(n_551),
.Y(n_10632)
);

OAI21xp5_ASAP7_75t_L g10633 ( 
.A1(n_10150),
.A2(n_551),
.B(n_552),
.Y(n_10633)
);

NAND2x1p5_ASAP7_75t_L g10634 ( 
.A(n_9987),
.B(n_1396),
.Y(n_10634)
);

NAND3x1_ASAP7_75t_L g10635 ( 
.A(n_10167),
.B(n_552),
.C(n_553),
.Y(n_10635)
);

AOI21xp5_ASAP7_75t_L g10636 ( 
.A1(n_9864),
.A2(n_552),
.B(n_553),
.Y(n_10636)
);

A2O1A1Ixp33_ASAP7_75t_L g10637 ( 
.A1(n_10166),
.A2(n_1398),
.B(n_1399),
.C(n_1397),
.Y(n_10637)
);

AOI21xp5_ASAP7_75t_L g10638 ( 
.A1(n_10031),
.A2(n_554),
.B(n_555),
.Y(n_10638)
);

INVx4_ASAP7_75t_L g10639 ( 
.A(n_10338),
.Y(n_10639)
);

AO31x2_ASAP7_75t_L g10640 ( 
.A1(n_10020),
.A2(n_556),
.A3(n_554),
.B(n_555),
.Y(n_10640)
);

OAI21x1_ASAP7_75t_L g10641 ( 
.A1(n_10074),
.A2(n_554),
.B(n_555),
.Y(n_10641)
);

AOI21xp5_ASAP7_75t_L g10642 ( 
.A1(n_9964),
.A2(n_556),
.B(n_557),
.Y(n_10642)
);

NAND2xp5_ASAP7_75t_L g10643 ( 
.A(n_10324),
.B(n_9827),
.Y(n_10643)
);

BUFx6f_ASAP7_75t_L g10644 ( 
.A(n_10160),
.Y(n_10644)
);

INVx1_ASAP7_75t_L g10645 ( 
.A(n_9909),
.Y(n_10645)
);

NAND2xp5_ASAP7_75t_L g10646 ( 
.A(n_9810),
.B(n_1397),
.Y(n_10646)
);

BUFx2_ASAP7_75t_L g10647 ( 
.A(n_10346),
.Y(n_10647)
);

AOI21xp5_ASAP7_75t_L g10648 ( 
.A1(n_10114),
.A2(n_557),
.B(n_558),
.Y(n_10648)
);

OAI22xp5_ASAP7_75t_L g10649 ( 
.A1(n_10107),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_10649)
);

AO21x1_ASAP7_75t_L g10650 ( 
.A1(n_10283),
.A2(n_558),
.B(n_559),
.Y(n_10650)
);

AOI21xp5_ASAP7_75t_L g10651 ( 
.A1(n_9797),
.A2(n_559),
.B(n_560),
.Y(n_10651)
);

OAI21x1_ASAP7_75t_L g10652 ( 
.A1(n_10081),
.A2(n_560),
.B(n_561),
.Y(n_10652)
);

NAND2xp5_ASAP7_75t_L g10653 ( 
.A(n_9853),
.B(n_1399),
.Y(n_10653)
);

INVx1_ASAP7_75t_L g10654 ( 
.A(n_9926),
.Y(n_10654)
);

OAI21x1_ASAP7_75t_L g10655 ( 
.A1(n_10087),
.A2(n_561),
.B(n_562),
.Y(n_10655)
);

NAND2xp5_ASAP7_75t_SL g10656 ( 
.A(n_10187),
.B(n_1401),
.Y(n_10656)
);

OAI21x1_ASAP7_75t_L g10657 ( 
.A1(n_10093),
.A2(n_10108),
.B(n_10101),
.Y(n_10657)
);

NAND2xp5_ASAP7_75t_L g10658 ( 
.A(n_10305),
.B(n_10121),
.Y(n_10658)
);

OAI21x1_ASAP7_75t_L g10659 ( 
.A1(n_10126),
.A2(n_562),
.B(n_563),
.Y(n_10659)
);

NAND2xp5_ASAP7_75t_L g10660 ( 
.A(n_10029),
.B(n_1401),
.Y(n_10660)
);

NAND2xp5_ASAP7_75t_L g10661 ( 
.A(n_10092),
.B(n_1402),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_9933),
.Y(n_10662)
);

OA21x2_ASAP7_75t_L g10663 ( 
.A1(n_10241),
.A2(n_1404),
.B(n_1403),
.Y(n_10663)
);

OAI21x1_ASAP7_75t_L g10664 ( 
.A1(n_10136),
.A2(n_562),
.B(n_563),
.Y(n_10664)
);

AOI221x1_ASAP7_75t_L g10665 ( 
.A1(n_10272),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.C(n_567),
.Y(n_10665)
);

AOI21xp5_ASAP7_75t_L g10666 ( 
.A1(n_10229),
.A2(n_564),
.B(n_565),
.Y(n_10666)
);

NAND2xp5_ASAP7_75t_L g10667 ( 
.A(n_10011),
.B(n_1403),
.Y(n_10667)
);

HB1xp67_ASAP7_75t_L g10668 ( 
.A(n_9892),
.Y(n_10668)
);

NOR2xp33_ASAP7_75t_L g10669 ( 
.A(n_9934),
.B(n_1404),
.Y(n_10669)
);

INVx2_ASAP7_75t_L g10670 ( 
.A(n_10329),
.Y(n_10670)
);

OAI21xp5_ASAP7_75t_L g10671 ( 
.A1(n_10220),
.A2(n_564),
.B(n_565),
.Y(n_10671)
);

AOI21xp5_ASAP7_75t_SL g10672 ( 
.A1(n_10127),
.A2(n_566),
.B(n_567),
.Y(n_10672)
);

NOR2xp33_ASAP7_75t_L g10673 ( 
.A(n_9953),
.B(n_1405),
.Y(n_10673)
);

NAND2x1p5_ASAP7_75t_L g10674 ( 
.A(n_10055),
.B(n_9944),
.Y(n_10674)
);

AOI221x1_ASAP7_75t_L g10675 ( 
.A1(n_10078),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.C(n_569),
.Y(n_10675)
);

AOI21xp5_ASAP7_75t_L g10676 ( 
.A1(n_10052),
.A2(n_568),
.B(n_569),
.Y(n_10676)
);

NAND2xp5_ASAP7_75t_L g10677 ( 
.A(n_10022),
.B(n_1405),
.Y(n_10677)
);

OAI21xp33_ASAP7_75t_L g10678 ( 
.A1(n_10361),
.A2(n_570),
.B(n_571),
.Y(n_10678)
);

OAI21x1_ASAP7_75t_L g10679 ( 
.A1(n_10138),
.A2(n_10148),
.B(n_10140),
.Y(n_10679)
);

NAND2xp5_ASAP7_75t_SL g10680 ( 
.A(n_9950),
.B(n_1406),
.Y(n_10680)
);

AOI21xp5_ASAP7_75t_L g10681 ( 
.A1(n_10045),
.A2(n_570),
.B(n_571),
.Y(n_10681)
);

NAND2xp5_ASAP7_75t_L g10682 ( 
.A(n_10348),
.B(n_1406),
.Y(n_10682)
);

NOR2xp33_ASAP7_75t_L g10683 ( 
.A(n_10188),
.B(n_10335),
.Y(n_10683)
);

BUFx6f_ASAP7_75t_L g10684 ( 
.A(n_9957),
.Y(n_10684)
);

AOI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_10095),
.A2(n_570),
.B(n_572),
.Y(n_10685)
);

NAND2xp5_ASAP7_75t_L g10686 ( 
.A(n_10038),
.B(n_1407),
.Y(n_10686)
);

AND2x2_ASAP7_75t_L g10687 ( 
.A(n_9777),
.B(n_1407),
.Y(n_10687)
);

OAI21x1_ASAP7_75t_L g10688 ( 
.A1(n_10151),
.A2(n_572),
.B(n_573),
.Y(n_10688)
);

AO31x2_ASAP7_75t_L g10689 ( 
.A1(n_10146),
.A2(n_574),
.A3(n_572),
.B(n_573),
.Y(n_10689)
);

AND2x2_ASAP7_75t_L g10690 ( 
.A(n_10192),
.B(n_1408),
.Y(n_10690)
);

AOI31xp67_ASAP7_75t_L g10691 ( 
.A1(n_10193),
.A2(n_576),
.A3(n_574),
.B(n_575),
.Y(n_10691)
);

AOI21xp5_ASAP7_75t_L g10692 ( 
.A1(n_10116),
.A2(n_574),
.B(n_575),
.Y(n_10692)
);

OAI21xp5_ASAP7_75t_L g10693 ( 
.A1(n_10176),
.A2(n_575),
.B(n_576),
.Y(n_10693)
);

AOI21xp5_ASAP7_75t_L g10694 ( 
.A1(n_10133),
.A2(n_577),
.B(n_578),
.Y(n_10694)
);

AO31x2_ASAP7_75t_L g10695 ( 
.A1(n_10226),
.A2(n_579),
.A3(n_577),
.B(n_578),
.Y(n_10695)
);

AOI21xp5_ASAP7_75t_L g10696 ( 
.A1(n_10030),
.A2(n_579),
.B(n_580),
.Y(n_10696)
);

INVx1_ASAP7_75t_SL g10697 ( 
.A(n_9937),
.Y(n_10697)
);

OAI21x1_ASAP7_75t_L g10698 ( 
.A1(n_10157),
.A2(n_579),
.B(n_580),
.Y(n_10698)
);

AND2x2_ASAP7_75t_L g10699 ( 
.A(n_9988),
.B(n_1408),
.Y(n_10699)
);

AO21x1_ASAP7_75t_L g10700 ( 
.A1(n_10013),
.A2(n_580),
.B(n_581),
.Y(n_10700)
);

AOI21xp33_ASAP7_75t_L g10701 ( 
.A1(n_9800),
.A2(n_582),
.B(n_583),
.Y(n_10701)
);

AOI21xp5_ASAP7_75t_L g10702 ( 
.A1(n_10310),
.A2(n_582),
.B(n_583),
.Y(n_10702)
);

NAND2xp5_ASAP7_75t_L g10703 ( 
.A(n_10044),
.B(n_1409),
.Y(n_10703)
);

INVx4_ASAP7_75t_L g10704 ( 
.A(n_9957),
.Y(n_10704)
);

NAND2xp5_ASAP7_75t_L g10705 ( 
.A(n_10046),
.B(n_1411),
.Y(n_10705)
);

AOI21xp5_ASAP7_75t_L g10706 ( 
.A1(n_10041),
.A2(n_582),
.B(n_583),
.Y(n_10706)
);

AOI21xp5_ASAP7_75t_L g10707 ( 
.A1(n_10245),
.A2(n_584),
.B(n_585),
.Y(n_10707)
);

INVx2_ASAP7_75t_L g10708 ( 
.A(n_9897),
.Y(n_10708)
);

AND2x2_ASAP7_75t_SL g10709 ( 
.A(n_10048),
.B(n_584),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_9903),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_SL g10711 ( 
.A(n_10369),
.B(n_1411),
.Y(n_10711)
);

NAND2xp5_ASAP7_75t_L g10712 ( 
.A(n_10068),
.B(n_1412),
.Y(n_10712)
);

AOI21xp5_ASAP7_75t_L g10713 ( 
.A1(n_10063),
.A2(n_584),
.B(n_585),
.Y(n_10713)
);

BUFx2_ASAP7_75t_L g10714 ( 
.A(n_9888),
.Y(n_10714)
);

NOR2xp67_ASAP7_75t_L g10715 ( 
.A(n_10316),
.B(n_585),
.Y(n_10715)
);

CKINVDCx16_ASAP7_75t_R g10716 ( 
.A(n_9901),
.Y(n_10716)
);

O2A1O1Ixp5_ASAP7_75t_SL g10717 ( 
.A1(n_10362),
.A2(n_588),
.B(n_586),
.C(n_587),
.Y(n_10717)
);

OAI22x1_ASAP7_75t_L g10718 ( 
.A1(n_9911),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_10718)
);

AND3x1_ASAP7_75t_L g10719 ( 
.A(n_10235),
.B(n_586),
.C(n_587),
.Y(n_10719)
);

AND2x2_ASAP7_75t_L g10720 ( 
.A(n_10147),
.B(n_1413),
.Y(n_10720)
);

OAI21x1_ASAP7_75t_L g10721 ( 
.A1(n_9939),
.A2(n_588),
.B(n_589),
.Y(n_10721)
);

NAND2xp5_ASAP7_75t_SL g10722 ( 
.A(n_10015),
.B(n_1413),
.Y(n_10722)
);

AOI22xp5_ASAP7_75t_L g10723 ( 
.A1(n_10059),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_10723)
);

NAND3xp33_ASAP7_75t_L g10724 ( 
.A(n_10266),
.B(n_589),
.C(n_590),
.Y(n_10724)
);

OAI21x1_ASAP7_75t_L g10725 ( 
.A1(n_9941),
.A2(n_590),
.B(n_591),
.Y(n_10725)
);

CKINVDCx20_ASAP7_75t_R g10726 ( 
.A(n_9884),
.Y(n_10726)
);

BUFx3_ASAP7_75t_L g10727 ( 
.A(n_10299),
.Y(n_10727)
);

AOI21xp5_ASAP7_75t_L g10728 ( 
.A1(n_10347),
.A2(n_591),
.B(n_592),
.Y(n_10728)
);

OAI21x1_ASAP7_75t_L g10729 ( 
.A1(n_9954),
.A2(n_592),
.B(n_593),
.Y(n_10729)
);

INVx1_ASAP7_75t_L g10730 ( 
.A(n_9912),
.Y(n_10730)
);

OAI21xp5_ASAP7_75t_L g10731 ( 
.A1(n_10274),
.A2(n_593),
.B(n_594),
.Y(n_10731)
);

NAND2xp5_ASAP7_75t_SL g10732 ( 
.A(n_10343),
.B(n_10178),
.Y(n_10732)
);

AOI21x1_ASAP7_75t_L g10733 ( 
.A1(n_9924),
.A2(n_593),
.B(n_594),
.Y(n_10733)
);

AOI21x1_ASAP7_75t_L g10734 ( 
.A1(n_9943),
.A2(n_594),
.B(n_595),
.Y(n_10734)
);

AND2x2_ASAP7_75t_L g10735 ( 
.A(n_10328),
.B(n_1414),
.Y(n_10735)
);

NAND2xp33_ASAP7_75t_SL g10736 ( 
.A(n_10288),
.B(n_10344),
.Y(n_10736)
);

AOI21xp5_ASAP7_75t_L g10737 ( 
.A1(n_10270),
.A2(n_596),
.B(n_597),
.Y(n_10737)
);

BUFx2_ASAP7_75t_L g10738 ( 
.A(n_10323),
.Y(n_10738)
);

OAI21xp33_ASAP7_75t_L g10739 ( 
.A1(n_10326),
.A2(n_596),
.B(n_597),
.Y(n_10739)
);

OA21x2_ASAP7_75t_L g10740 ( 
.A1(n_10248),
.A2(n_1415),
.B(n_1414),
.Y(n_10740)
);

OAI21xp5_ASAP7_75t_L g10741 ( 
.A1(n_10311),
.A2(n_596),
.B(n_598),
.Y(n_10741)
);

OAI21x1_ASAP7_75t_L g10742 ( 
.A1(n_9956),
.A2(n_598),
.B(n_599),
.Y(n_10742)
);

INVx1_ASAP7_75t_L g10743 ( 
.A(n_9913),
.Y(n_10743)
);

NAND2xp5_ASAP7_75t_L g10744 ( 
.A(n_10077),
.B(n_1415),
.Y(n_10744)
);

INVx2_ASAP7_75t_L g10745 ( 
.A(n_9914),
.Y(n_10745)
);

AOI21xp5_ASAP7_75t_L g10746 ( 
.A1(n_10275),
.A2(n_598),
.B(n_600),
.Y(n_10746)
);

OAI22xp5_ASAP7_75t_L g10747 ( 
.A1(n_10230),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_10747)
);

AOI21x1_ASAP7_75t_SL g10748 ( 
.A1(n_10208),
.A2(n_600),
.B(n_601),
.Y(n_10748)
);

NAND2xp5_ASAP7_75t_L g10749 ( 
.A(n_10085),
.B(n_1416),
.Y(n_10749)
);

BUFx3_ASAP7_75t_L g10750 ( 
.A(n_10016),
.Y(n_10750)
);

AOI21xp5_ASAP7_75t_L g10751 ( 
.A1(n_10243),
.A2(n_601),
.B(n_602),
.Y(n_10751)
);

CKINVDCx20_ASAP7_75t_R g10752 ( 
.A(n_9948),
.Y(n_10752)
);

INVx1_ASAP7_75t_L g10753 ( 
.A(n_9931),
.Y(n_10753)
);

INVx1_ASAP7_75t_L g10754 ( 
.A(n_9935),
.Y(n_10754)
);

A2O1A1Ixp33_ASAP7_75t_L g10755 ( 
.A1(n_10357),
.A2(n_1417),
.B(n_1418),
.C(n_1416),
.Y(n_10755)
);

INVx1_ASAP7_75t_L g10756 ( 
.A(n_9936),
.Y(n_10756)
);

NAND2xp5_ASAP7_75t_L g10757 ( 
.A(n_10086),
.B(n_1417),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_L g10758 ( 
.A(n_10102),
.B(n_1418),
.Y(n_10758)
);

AO21x1_ASAP7_75t_L g10759 ( 
.A1(n_9792),
.A2(n_9794),
.B(n_9793),
.Y(n_10759)
);

NAND2xp33_ASAP7_75t_L g10760 ( 
.A(n_10033),
.B(n_602),
.Y(n_10760)
);

HB1xp67_ASAP7_75t_L g10761 ( 
.A(n_9938),
.Y(n_10761)
);

AOI21xp5_ASAP7_75t_L g10762 ( 
.A1(n_10280),
.A2(n_603),
.B(n_604),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_9942),
.Y(n_10763)
);

BUFx3_ASAP7_75t_L g10764 ( 
.A(n_10053),
.Y(n_10764)
);

OAI22xp5_ASAP7_75t_L g10765 ( 
.A1(n_10230),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_10765)
);

INVx1_ASAP7_75t_L g10766 ( 
.A(n_9973),
.Y(n_10766)
);

AND2x2_ASAP7_75t_L g10767 ( 
.A(n_10315),
.B(n_1419),
.Y(n_10767)
);

AO21x1_ASAP7_75t_L g10768 ( 
.A1(n_9990),
.A2(n_604),
.B(n_605),
.Y(n_10768)
);

NOR2xp33_ASAP7_75t_L g10769 ( 
.A(n_10354),
.B(n_10358),
.Y(n_10769)
);

BUFx6f_ASAP7_75t_L g10770 ( 
.A(n_10021),
.Y(n_10770)
);

NAND2xp5_ASAP7_75t_L g10771 ( 
.A(n_10105),
.B(n_1419),
.Y(n_10771)
);

NAND2xp5_ASAP7_75t_L g10772 ( 
.A(n_10115),
.B(n_1420),
.Y(n_10772)
);

CKINVDCx11_ASAP7_75t_R g10773 ( 
.A(n_10336),
.Y(n_10773)
);

OAI21x1_ASAP7_75t_L g10774 ( 
.A1(n_9972),
.A2(n_10056),
.B(n_10058),
.Y(n_10774)
);

NAND2x1p5_ASAP7_75t_L g10775 ( 
.A(n_10153),
.B(n_1420),
.Y(n_10775)
);

OAI21xp5_ASAP7_75t_L g10776 ( 
.A1(n_10317),
.A2(n_605),
.B(n_606),
.Y(n_10776)
);

NAND2xp5_ASAP7_75t_L g10777 ( 
.A(n_10132),
.B(n_1422),
.Y(n_10777)
);

CKINVDCx6p67_ASAP7_75t_R g10778 ( 
.A(n_10042),
.Y(n_10778)
);

NAND2xp5_ASAP7_75t_L g10779 ( 
.A(n_10142),
.B(n_1423),
.Y(n_10779)
);

INVx1_ASAP7_75t_L g10780 ( 
.A(n_10333),
.Y(n_10780)
);

NAND2xp5_ASAP7_75t_L g10781 ( 
.A(n_10144),
.B(n_1423),
.Y(n_10781)
);

NAND2xp5_ASAP7_75t_L g10782 ( 
.A(n_10145),
.B(n_1424),
.Y(n_10782)
);

INVx1_ASAP7_75t_L g10783 ( 
.A(n_9899),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_L g10784 ( 
.A(n_10149),
.B(n_1424),
.Y(n_10784)
);

INVx1_ASAP7_75t_L g10785 ( 
.A(n_9899),
.Y(n_10785)
);

OAI22xp5_ASAP7_75t_L g10786 ( 
.A1(n_10084),
.A2(n_10141),
.B1(n_10267),
.B2(n_10002),
.Y(n_10786)
);

AOI21xp5_ASAP7_75t_L g10787 ( 
.A1(n_10277),
.A2(n_606),
.B(n_607),
.Y(n_10787)
);

AO31x2_ASAP7_75t_L g10788 ( 
.A1(n_10342),
.A2(n_608),
.A3(n_606),
.B(n_607),
.Y(n_10788)
);

O2A1O1Ixp33_ASAP7_75t_L g10789 ( 
.A1(n_10073),
.A2(n_609),
.B(n_607),
.C(n_608),
.Y(n_10789)
);

NAND2x1_ASAP7_75t_L g10790 ( 
.A(n_9880),
.B(n_1425),
.Y(n_10790)
);

AOI21xp5_ASAP7_75t_L g10791 ( 
.A1(n_10281),
.A2(n_608),
.B(n_609),
.Y(n_10791)
);

NAND2xp5_ASAP7_75t_L g10792 ( 
.A(n_10161),
.B(n_1425),
.Y(n_10792)
);

INVx1_ASAP7_75t_L g10793 ( 
.A(n_10189),
.Y(n_10793)
);

AOI21xp5_ASAP7_75t_L g10794 ( 
.A1(n_9974),
.A2(n_609),
.B(n_610),
.Y(n_10794)
);

AOI21xp5_ASAP7_75t_L g10795 ( 
.A1(n_10264),
.A2(n_610),
.B(n_611),
.Y(n_10795)
);

INVx2_ASAP7_75t_L g10796 ( 
.A(n_9916),
.Y(n_10796)
);

NAND2xp5_ASAP7_75t_L g10797 ( 
.A(n_10169),
.B(n_1426),
.Y(n_10797)
);

NAND2x1p5_ASAP7_75t_L g10798 ( 
.A(n_9999),
.B(n_1426),
.Y(n_10798)
);

O2A1O1Ixp5_ASAP7_75t_SL g10799 ( 
.A1(n_10225),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_10799)
);

O2A1O1Ixp33_ASAP7_75t_L g10800 ( 
.A1(n_9781),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_10800)
);

AOI21xp5_ASAP7_75t_SL g10801 ( 
.A1(n_9989),
.A2(n_613),
.B(n_614),
.Y(n_10801)
);

OAI21xp5_ASAP7_75t_SL g10802 ( 
.A1(n_10112),
.A2(n_614),
.B(n_615),
.Y(n_10802)
);

AOI21xp5_ASAP7_75t_L g10803 ( 
.A1(n_10352),
.A2(n_614),
.B(n_615),
.Y(n_10803)
);

AOI21xp5_ASAP7_75t_L g10804 ( 
.A1(n_10004),
.A2(n_615),
.B(n_616),
.Y(n_10804)
);

NAND2xp5_ASAP7_75t_L g10805 ( 
.A(n_10174),
.B(n_1427),
.Y(n_10805)
);

NAND2xp5_ASAP7_75t_L g10806 ( 
.A(n_10175),
.B(n_1427),
.Y(n_10806)
);

OAI21xp5_ASAP7_75t_SL g10807 ( 
.A1(n_10298),
.A2(n_616),
.B(n_617),
.Y(n_10807)
);

OAI22xp5_ASAP7_75t_L g10808 ( 
.A1(n_9788),
.A2(n_618),
.B1(n_616),
.B2(n_617),
.Y(n_10808)
);

BUFx2_ASAP7_75t_L g10809 ( 
.A(n_10359),
.Y(n_10809)
);

AOI21xp5_ASAP7_75t_L g10810 ( 
.A1(n_9921),
.A2(n_617),
.B(n_618),
.Y(n_10810)
);

AND2x2_ASAP7_75t_SL g10811 ( 
.A(n_9826),
.B(n_618),
.Y(n_10811)
);

AND2x2_ASAP7_75t_L g10812 ( 
.A(n_9866),
.B(n_1428),
.Y(n_10812)
);

INVxp67_ASAP7_75t_SL g10813 ( 
.A(n_10163),
.Y(n_10813)
);

NAND2xp5_ASAP7_75t_L g10814 ( 
.A(n_10181),
.B(n_1428),
.Y(n_10814)
);

HB1xp67_ASAP7_75t_L g10815 ( 
.A(n_9789),
.Y(n_10815)
);

OAI21xp5_ASAP7_75t_L g10816 ( 
.A1(n_10191),
.A2(n_619),
.B(n_620),
.Y(n_10816)
);

BUFx8_ASAP7_75t_L g10817 ( 
.A(n_10042),
.Y(n_10817)
);

AOI21x1_ASAP7_75t_L g10818 ( 
.A1(n_10060),
.A2(n_619),
.B(n_620),
.Y(n_10818)
);

OAI21x1_ASAP7_75t_L g10819 ( 
.A1(n_10223),
.A2(n_620),
.B(n_621),
.Y(n_10819)
);

OAI21x1_ASAP7_75t_L g10820 ( 
.A1(n_10197),
.A2(n_621),
.B(n_622),
.Y(n_10820)
);

BUFx2_ASAP7_75t_L g10821 ( 
.A(n_10205),
.Y(n_10821)
);

OAI21x1_ASAP7_75t_L g10822 ( 
.A1(n_10212),
.A2(n_10263),
.B(n_10162),
.Y(n_10822)
);

AND2x2_ASAP7_75t_L g10823 ( 
.A(n_9982),
.B(n_1430),
.Y(n_10823)
);

AOI21xp5_ASAP7_75t_L g10824 ( 
.A1(n_9940),
.A2(n_621),
.B(n_622),
.Y(n_10824)
);

INVx1_ASAP7_75t_L g10825 ( 
.A(n_10236),
.Y(n_10825)
);

AND2x4_ASAP7_75t_L g10826 ( 
.A(n_10286),
.B(n_1431),
.Y(n_10826)
);

AOI21x1_ASAP7_75t_L g10827 ( 
.A1(n_10080),
.A2(n_623),
.B(n_624),
.Y(n_10827)
);

AO31x2_ASAP7_75t_L g10828 ( 
.A1(n_10179),
.A2(n_625),
.A3(n_623),
.B(n_624),
.Y(n_10828)
);

AO31x2_ASAP7_75t_L g10829 ( 
.A1(n_10090),
.A2(n_626),
.A3(n_623),
.B(n_625),
.Y(n_10829)
);

NOR2xp33_ASAP7_75t_L g10830 ( 
.A(n_10242),
.B(n_1431),
.Y(n_10830)
);

AOI21xp5_ASAP7_75t_L g10831 ( 
.A1(n_9968),
.A2(n_626),
.B(n_627),
.Y(n_10831)
);

OAI21x1_ASAP7_75t_L g10832 ( 
.A1(n_10255),
.A2(n_626),
.B(n_627),
.Y(n_10832)
);

NAND2x1_ASAP7_75t_L g10833 ( 
.A(n_9880),
.B(n_1432),
.Y(n_10833)
);

O2A1O1Ixp33_ASAP7_75t_L g10834 ( 
.A1(n_10195),
.A2(n_629),
.B(n_627),
.C(n_628),
.Y(n_10834)
);

O2A1O1Ixp5_ASAP7_75t_SL g10835 ( 
.A1(n_10216),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_10835)
);

AND2x2_ASAP7_75t_L g10836 ( 
.A(n_10159),
.B(n_1433),
.Y(n_10836)
);

NAND2xp5_ASAP7_75t_L g10837 ( 
.A(n_10199),
.B(n_1434),
.Y(n_10837)
);

AOI21xp5_ASAP7_75t_L g10838 ( 
.A1(n_10273),
.A2(n_628),
.B(n_629),
.Y(n_10838)
);

INVx1_ASAP7_75t_L g10839 ( 
.A(n_10364),
.Y(n_10839)
);

AOI21xp5_ASAP7_75t_L g10840 ( 
.A1(n_10238),
.A2(n_630),
.B(n_631),
.Y(n_10840)
);

BUFx6f_ASAP7_75t_L g10841 ( 
.A(n_10021),
.Y(n_10841)
);

O2A1O1Ixp33_ASAP7_75t_L g10842 ( 
.A1(n_10244),
.A2(n_633),
.B(n_631),
.C(n_632),
.Y(n_10842)
);

NOR2xp33_ASAP7_75t_L g10843 ( 
.A(n_10293),
.B(n_1435),
.Y(n_10843)
);

NAND2xp5_ASAP7_75t_L g10844 ( 
.A(n_10214),
.B(n_1435),
.Y(n_10844)
);

AOI21xp5_ASAP7_75t_L g10845 ( 
.A1(n_9814),
.A2(n_9851),
.B(n_10217),
.Y(n_10845)
);

AOI21x1_ASAP7_75t_L g10846 ( 
.A1(n_10259),
.A2(n_632),
.B(n_633),
.Y(n_10846)
);

OAI21x1_ASAP7_75t_L g10847 ( 
.A1(n_10436),
.A2(n_10137),
.B(n_10143),
.Y(n_10847)
);

OA21x2_ASAP7_75t_L g10848 ( 
.A1(n_10643),
.A2(n_10306),
.B(n_10304),
.Y(n_10848)
);

AO21x2_ASAP7_75t_L g10849 ( 
.A1(n_10815),
.A2(n_10780),
.B(n_10613),
.Y(n_10849)
);

OAI21x1_ASAP7_75t_L g10850 ( 
.A1(n_10381),
.A2(n_10211),
.B(n_9996),
.Y(n_10850)
);

BUFx2_ASAP7_75t_L g10851 ( 
.A(n_10809),
.Y(n_10851)
);

INVx2_ASAP7_75t_L g10852 ( 
.A(n_10379),
.Y(n_10852)
);

NAND2xp5_ASAP7_75t_L g10853 ( 
.A(n_10564),
.B(n_10339),
.Y(n_10853)
);

INVx2_ASAP7_75t_L g10854 ( 
.A(n_10386),
.Y(n_10854)
);

NAND2x1p5_ASAP7_75t_L g10855 ( 
.A(n_10821),
.B(n_10353),
.Y(n_10855)
);

INVx2_ASAP7_75t_L g10856 ( 
.A(n_10406),
.Y(n_10856)
);

AO21x2_ASAP7_75t_L g10857 ( 
.A1(n_10594),
.A2(n_10231),
.B(n_10219),
.Y(n_10857)
);

NAND2xp5_ASAP7_75t_L g10858 ( 
.A(n_10510),
.B(n_9789),
.Y(n_10858)
);

AOI21xp5_ASAP7_75t_L g10859 ( 
.A1(n_10408),
.A2(n_10279),
.B(n_10057),
.Y(n_10859)
);

OAI21x1_ASAP7_75t_SL g10860 ( 
.A1(n_10604),
.A2(n_10119),
.B(n_10368),
.Y(n_10860)
);

BUFx6f_ASAP7_75t_L g10861 ( 
.A(n_10580),
.Y(n_10861)
);

INVx1_ASAP7_75t_L g10862 ( 
.A(n_10414),
.Y(n_10862)
);

BUFx3_ASAP7_75t_L g10863 ( 
.A(n_10388),
.Y(n_10863)
);

AOI21x1_ASAP7_75t_L g10864 ( 
.A1(n_10656),
.A2(n_10265),
.B(n_9882),
.Y(n_10864)
);

INVx1_ASAP7_75t_L g10865 ( 
.A(n_10462),
.Y(n_10865)
);

NAND2x1p5_ASAP7_75t_L g10866 ( 
.A(n_10615),
.B(n_10295),
.Y(n_10866)
);

OAI21xp5_ASAP7_75t_L g10867 ( 
.A1(n_10401),
.A2(n_10345),
.B(n_10308),
.Y(n_10867)
);

NAND2x1p5_ASAP7_75t_L g10868 ( 
.A(n_10433),
.B(n_10023),
.Y(n_10868)
);

OA21x2_ASAP7_75t_L g10869 ( 
.A1(n_10623),
.A2(n_10289),
.B(n_10341),
.Y(n_10869)
);

OAI21x1_ASAP7_75t_L g10870 ( 
.A1(n_10450),
.A2(n_10258),
.B(n_10233),
.Y(n_10870)
);

OR2x2_ASAP7_75t_L g10871 ( 
.A(n_10514),
.B(n_10177),
.Y(n_10871)
);

OA21x2_ASAP7_75t_L g10872 ( 
.A1(n_10839),
.A2(n_10340),
.B(n_10254),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_10417),
.Y(n_10873)
);

AND2x4_ASAP7_75t_L g10874 ( 
.A(n_10534),
.B(n_10023),
.Y(n_10874)
);

INVx3_ASAP7_75t_L g10875 ( 
.A(n_10482),
.Y(n_10875)
);

INVxp67_ASAP7_75t_SL g10876 ( 
.A(n_10566),
.Y(n_10876)
);

AND2x2_ASAP7_75t_L g10877 ( 
.A(n_10526),
.B(n_10321),
.Y(n_10877)
);

OAI21x1_ASAP7_75t_SL g10878 ( 
.A1(n_10430),
.A2(n_10319),
.B(n_10262),
.Y(n_10878)
);

OAI21xp5_ASAP7_75t_L g10879 ( 
.A1(n_10404),
.A2(n_10234),
.B(n_10284),
.Y(n_10879)
);

BUFx6f_ASAP7_75t_L g10880 ( 
.A(n_10426),
.Y(n_10880)
);

OAI21x1_ASAP7_75t_L g10881 ( 
.A1(n_10774),
.A2(n_10301),
.B(n_10356),
.Y(n_10881)
);

OR2x2_ASAP7_75t_L g10882 ( 
.A(n_10420),
.B(n_10261),
.Y(n_10882)
);

INVx4_ASAP7_75t_L g10883 ( 
.A(n_10538),
.Y(n_10883)
);

OAI21x1_ASAP7_75t_L g10884 ( 
.A1(n_10473),
.A2(n_10363),
.B(n_9838),
.Y(n_10884)
);

AND2x4_ASAP7_75t_L g10885 ( 
.A(n_10584),
.B(n_10054),
.Y(n_10885)
);

HB1xp67_ASAP7_75t_L g10886 ( 
.A(n_10793),
.Y(n_10886)
);

OAI21x1_ASAP7_75t_L g10887 ( 
.A1(n_10657),
.A2(n_10349),
.B(n_10152),
.Y(n_10887)
);

OAI21x1_ASAP7_75t_L g10888 ( 
.A1(n_10679),
.A2(n_10097),
.B(n_10282),
.Y(n_10888)
);

INVxp67_ASAP7_75t_L g10889 ( 
.A(n_10668),
.Y(n_10889)
);

AOI22xp5_ASAP7_75t_L g10890 ( 
.A1(n_10550),
.A2(n_10042),
.B1(n_9880),
.B2(n_10033),
.Y(n_10890)
);

INVx2_ASAP7_75t_L g10891 ( 
.A(n_10395),
.Y(n_10891)
);

NOR2xp33_ASAP7_75t_L g10892 ( 
.A(n_10716),
.B(n_10376),
.Y(n_10892)
);

AND2x4_ASAP7_75t_L g10893 ( 
.A(n_10647),
.B(n_10054),
.Y(n_10893)
);

OAI21x1_ASAP7_75t_L g10894 ( 
.A1(n_10432),
.A2(n_9970),
.B(n_9900),
.Y(n_10894)
);

AOI22xp33_ASAP7_75t_L g10895 ( 
.A1(n_10380),
.A2(n_10332),
.B1(n_10371),
.B2(n_10370),
.Y(n_10895)
);

OAI22xp5_ASAP7_75t_L g10896 ( 
.A1(n_10458),
.A2(n_9816),
.B1(n_9843),
.B2(n_10355),
.Y(n_10896)
);

OA21x2_ASAP7_75t_L g10897 ( 
.A1(n_10486),
.A2(n_10303),
.B(n_10302),
.Y(n_10897)
);

INVxp67_ASAP7_75t_SL g10898 ( 
.A(n_10761),
.Y(n_10898)
);

NAND2xp5_ASAP7_75t_L g10899 ( 
.A(n_10568),
.B(n_9976),
.Y(n_10899)
);

AOI21xp5_ASAP7_75t_L g10900 ( 
.A1(n_10624),
.A2(n_10351),
.B(n_9977),
.Y(n_10900)
);

AOI22xp5_ASAP7_75t_L g10901 ( 
.A1(n_10619),
.A2(n_10205),
.B1(n_10183),
.B2(n_10050),
.Y(n_10901)
);

INVx1_ASAP7_75t_SL g10902 ( 
.A(n_10605),
.Y(n_10902)
);

NOR2xp67_ASAP7_75t_L g10903 ( 
.A(n_10658),
.B(n_10598),
.Y(n_10903)
);

AND2x4_ASAP7_75t_L g10904 ( 
.A(n_10670),
.B(n_10082),
.Y(n_10904)
);

CKINVDCx5p33_ASAP7_75t_R g10905 ( 
.A(n_10416),
.Y(n_10905)
);

OAI21x1_ASAP7_75t_L g10906 ( 
.A1(n_10383),
.A2(n_10170),
.B(n_10062),
.Y(n_10906)
);

OR2x2_ASAP7_75t_L g10907 ( 
.A(n_10423),
.B(n_10320),
.Y(n_10907)
);

CKINVDCx20_ASAP7_75t_R g10908 ( 
.A(n_10592),
.Y(n_10908)
);

OAI22xp5_ASAP7_75t_L g10909 ( 
.A1(n_10637),
.A2(n_10082),
.B1(n_10131),
.B2(n_10106),
.Y(n_10909)
);

INVx1_ASAP7_75t_L g10910 ( 
.A(n_10425),
.Y(n_10910)
);

INVx5_ASAP7_75t_L g10911 ( 
.A(n_10489),
.Y(n_10911)
);

BUFx6f_ASAP7_75t_L g10912 ( 
.A(n_10426),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_10429),
.Y(n_10913)
);

AOI22x1_ASAP7_75t_L g10914 ( 
.A1(n_10396),
.A2(n_10240),
.B1(n_10088),
.B2(n_10069),
.Y(n_10914)
);

AOI21xp5_ASAP7_75t_L g10915 ( 
.A1(n_10397),
.A2(n_10494),
.B(n_10630),
.Y(n_10915)
);

NAND3xp33_ASAP7_75t_L g10916 ( 
.A(n_10411),
.B(n_9965),
.C(n_9967),
.Y(n_10916)
);

OA21x2_ASAP7_75t_L g10917 ( 
.A1(n_10783),
.A2(n_10785),
.B(n_10822),
.Y(n_10917)
);

OR2x6_ASAP7_75t_L g10918 ( 
.A(n_10674),
.B(n_10106),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_10451),
.Y(n_10919)
);

INVx1_ASAP7_75t_L g10920 ( 
.A(n_10456),
.Y(n_10920)
);

OR2x6_ASAP7_75t_L g10921 ( 
.A(n_10378),
.B(n_10131),
.Y(n_10921)
);

OA21x2_ASAP7_75t_L g10922 ( 
.A1(n_10539),
.A2(n_10111),
.B(n_10039),
.Y(n_10922)
);

BUFx2_ASAP7_75t_L g10923 ( 
.A(n_10738),
.Y(n_10923)
);

CKINVDCx5p33_ASAP7_75t_R g10924 ( 
.A(n_10726),
.Y(n_10924)
);

OAI21x1_ASAP7_75t_L g10925 ( 
.A1(n_10460),
.A2(n_10051),
.B(n_10250),
.Y(n_10925)
);

INVx2_ASAP7_75t_L g10926 ( 
.A(n_10457),
.Y(n_10926)
);

OAI21x1_ASAP7_75t_L g10927 ( 
.A1(n_10384),
.A2(n_10296),
.B(n_10278),
.Y(n_10927)
);

OA21x2_ASAP7_75t_L g10928 ( 
.A1(n_10428),
.A2(n_10309),
.B(n_10307),
.Y(n_10928)
);

AND2x4_ASAP7_75t_L g10929 ( 
.A(n_10530),
.B(n_10099),
.Y(n_10929)
);

INVx1_ASAP7_75t_L g10930 ( 
.A(n_10467),
.Y(n_10930)
);

INVx1_ASAP7_75t_SL g10931 ( 
.A(n_10773),
.Y(n_10931)
);

AND2x4_ASAP7_75t_L g10932 ( 
.A(n_10569),
.B(n_10109),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_10495),
.Y(n_10933)
);

INVx1_ASAP7_75t_L g10934 ( 
.A(n_10497),
.Y(n_10934)
);

BUFx10_ASAP7_75t_L g10935 ( 
.A(n_10440),
.Y(n_10935)
);

CKINVDCx16_ASAP7_75t_R g10936 ( 
.A(n_10599),
.Y(n_10936)
);

OAI21x1_ASAP7_75t_L g10937 ( 
.A1(n_10648),
.A2(n_10156),
.B(n_10130),
.Y(n_10937)
);

OAI21x1_ASAP7_75t_L g10938 ( 
.A1(n_10434),
.A2(n_10156),
.B(n_10130),
.Y(n_10938)
);

BUFx3_ASAP7_75t_L g10939 ( 
.A(n_10752),
.Y(n_10939)
);

BUFx3_ASAP7_75t_L g10940 ( 
.A(n_10727),
.Y(n_10940)
);

BUFx3_ASAP7_75t_L g10941 ( 
.A(n_10750),
.Y(n_10941)
);

OAI21x1_ASAP7_75t_L g10942 ( 
.A1(n_10810),
.A2(n_9896),
.B(n_10047),
.Y(n_10942)
);

INVx1_ASAP7_75t_L g10943 ( 
.A(n_10504),
.Y(n_10943)
);

OAI21x1_ASAP7_75t_L g10944 ( 
.A1(n_10825),
.A2(n_10047),
.B(n_10364),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_10505),
.Y(n_10945)
);

OA21x2_ASAP7_75t_L g10946 ( 
.A1(n_10816),
.A2(n_9994),
.B(n_10269),
.Y(n_10946)
);

INVx6_ASAP7_75t_L g10947 ( 
.A(n_10639),
.Y(n_10947)
);

INVx1_ASAP7_75t_L g10948 ( 
.A(n_10517),
.Y(n_10948)
);

INVx2_ASAP7_75t_L g10949 ( 
.A(n_10520),
.Y(n_10949)
);

INVx2_ASAP7_75t_L g10950 ( 
.A(n_10528),
.Y(n_10950)
);

INVx1_ASAP7_75t_L g10951 ( 
.A(n_10573),
.Y(n_10951)
);

AOI22x1_ASAP7_75t_L g10952 ( 
.A1(n_10410),
.A2(n_10224),
.B1(n_10076),
.B2(n_10269),
.Y(n_10952)
);

OAI21x1_ASAP7_75t_L g10953 ( 
.A1(n_10813),
.A2(n_10210),
.B(n_10201),
.Y(n_10953)
);

INVx2_ASAP7_75t_L g10954 ( 
.A(n_10796),
.Y(n_10954)
);

NAND2xp5_ASAP7_75t_L g10955 ( 
.A(n_10708),
.B(n_10076),
.Y(n_10955)
);

AOI22xp33_ASAP7_75t_L g10956 ( 
.A1(n_10576),
.A2(n_10205),
.B1(n_10210),
.B2(n_10201),
.Y(n_10956)
);

INVx3_ASAP7_75t_L g10957 ( 
.A(n_10470),
.Y(n_10957)
);

NOR2xp33_ASAP7_75t_L g10958 ( 
.A(n_10710),
.B(n_1436),
.Y(n_10958)
);

OAI21x1_ASAP7_75t_L g10959 ( 
.A1(n_10571),
.A2(n_10312),
.B(n_632),
.Y(n_10959)
);

BUFx12f_ASAP7_75t_L g10960 ( 
.A(n_10714),
.Y(n_10960)
);

INVx1_ASAP7_75t_L g10961 ( 
.A(n_10627),
.Y(n_10961)
);

AND2x2_ASAP7_75t_L g10962 ( 
.A(n_10582),
.B(n_10312),
.Y(n_10962)
);

OAI21x1_ASAP7_75t_L g10963 ( 
.A1(n_10733),
.A2(n_633),
.B(n_634),
.Y(n_10963)
);

AO21x1_ASAP7_75t_L g10964 ( 
.A1(n_10760),
.A2(n_634),
.B(n_635),
.Y(n_10964)
);

O2A1O1Ixp33_ASAP7_75t_L g10965 ( 
.A1(n_10540),
.A2(n_636),
.B(n_634),
.C(n_635),
.Y(n_10965)
);

OAI21x1_ASAP7_75t_L g10966 ( 
.A1(n_10734),
.A2(n_636),
.B(n_637),
.Y(n_10966)
);

INVx2_ASAP7_75t_L g10967 ( 
.A(n_10745),
.Y(n_10967)
);

OA21x2_ASAP7_75t_L g10968 ( 
.A1(n_10730),
.A2(n_636),
.B(n_637),
.Y(n_10968)
);

OAI22xp5_ASAP7_75t_L g10969 ( 
.A1(n_10492),
.A2(n_10453),
.B1(n_10427),
.B2(n_10583),
.Y(n_10969)
);

INVx3_ASAP7_75t_L g10970 ( 
.A(n_10475),
.Y(n_10970)
);

INVx1_ASAP7_75t_L g10971 ( 
.A(n_10743),
.Y(n_10971)
);

NAND2xp5_ASAP7_75t_L g10972 ( 
.A(n_10753),
.B(n_1436),
.Y(n_10972)
);

HB1xp67_ASAP7_75t_L g10973 ( 
.A(n_10754),
.Y(n_10973)
);

NAND2xp5_ASAP7_75t_L g10974 ( 
.A(n_10756),
.B(n_1437),
.Y(n_10974)
);

OAI21x1_ASAP7_75t_L g10975 ( 
.A1(n_10487),
.A2(n_637),
.B(n_638),
.Y(n_10975)
);

AND2x2_ASAP7_75t_L g10976 ( 
.A(n_10439),
.B(n_638),
.Y(n_10976)
);

O2A1O1Ixp33_ASAP7_75t_L g10977 ( 
.A1(n_10722),
.A2(n_640),
.B(n_638),
.C(n_639),
.Y(n_10977)
);

OAI21x1_ASAP7_75t_SL g10978 ( 
.A1(n_10650),
.A2(n_639),
.B(n_640),
.Y(n_10978)
);

OAI21xp5_ASAP7_75t_L g10979 ( 
.A1(n_10402),
.A2(n_1439),
.B(n_1438),
.Y(n_10979)
);

OAI21xp5_ASAP7_75t_L g10980 ( 
.A1(n_10500),
.A2(n_1439),
.B(n_1438),
.Y(n_10980)
);

NAND2xp5_ASAP7_75t_L g10981 ( 
.A(n_10763),
.B(n_1440),
.Y(n_10981)
);

AOI22x1_ASAP7_75t_L g10982 ( 
.A1(n_10718),
.A2(n_642),
.B1(n_639),
.B2(n_641),
.Y(n_10982)
);

AOI22x1_ASAP7_75t_L g10983 ( 
.A1(n_10525),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_10983)
);

AO21x1_ASAP7_75t_L g10984 ( 
.A1(n_10680),
.A2(n_10736),
.B(n_10802),
.Y(n_10984)
);

NOR2xp33_ASAP7_75t_L g10985 ( 
.A(n_10766),
.B(n_1440),
.Y(n_10985)
);

AOI22xp33_ASAP7_75t_L g10986 ( 
.A1(n_10626),
.A2(n_1442),
.B1(n_1443),
.B2(n_1441),
.Y(n_10986)
);

AOI21x1_ASAP7_75t_L g10987 ( 
.A1(n_10399),
.A2(n_641),
.B(n_643),
.Y(n_10987)
);

OAI21x1_ASAP7_75t_L g10988 ( 
.A1(n_10435),
.A2(n_643),
.B(n_644),
.Y(n_10988)
);

INVx2_ASAP7_75t_L g10989 ( 
.A(n_10616),
.Y(n_10989)
);

OAI21x1_ASAP7_75t_L g10990 ( 
.A1(n_10846),
.A2(n_644),
.B(n_645),
.Y(n_10990)
);

AO222x2_ASAP7_75t_L g10991 ( 
.A1(n_10585),
.A2(n_646),
.B1(n_648),
.B2(n_644),
.C1(n_645),
.C2(n_647),
.Y(n_10991)
);

INVx1_ASAP7_75t_L g10992 ( 
.A(n_10617),
.Y(n_10992)
);

OAI21x1_ASAP7_75t_SL g10993 ( 
.A1(n_10398),
.A2(n_645),
.B(n_646),
.Y(n_10993)
);

OA21x2_ASAP7_75t_L g10994 ( 
.A1(n_10403),
.A2(n_10454),
.B(n_10449),
.Y(n_10994)
);

INVx1_ASAP7_75t_L g10995 ( 
.A(n_10645),
.Y(n_10995)
);

AOI22xp5_ASAP7_75t_L g10996 ( 
.A1(n_10503),
.A2(n_1442),
.B1(n_1443),
.B2(n_1441),
.Y(n_10996)
);

NOR2xp33_ASAP7_75t_L g10997 ( 
.A(n_10610),
.B(n_1444),
.Y(n_10997)
);

INVx2_ASAP7_75t_L g10998 ( 
.A(n_10654),
.Y(n_10998)
);

AND2x2_ASAP7_75t_L g10999 ( 
.A(n_10466),
.B(n_646),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_10662),
.Y(n_11000)
);

NAND2xp5_ASAP7_75t_L g11001 ( 
.A(n_10507),
.B(n_1445),
.Y(n_11001)
);

CKINVDCx16_ASAP7_75t_R g11002 ( 
.A(n_10764),
.Y(n_11002)
);

OAI21x1_ASAP7_75t_L g11003 ( 
.A1(n_10721),
.A2(n_647),
.B(n_648),
.Y(n_11003)
);

NAND2xp5_ASAP7_75t_L g11004 ( 
.A(n_10601),
.B(n_1446),
.Y(n_11004)
);

NOR2xp67_ASAP7_75t_L g11005 ( 
.A(n_10560),
.B(n_647),
.Y(n_11005)
);

AOI21x1_ASAP7_75t_L g11006 ( 
.A1(n_10407),
.A2(n_648),
.B(n_649),
.Y(n_11006)
);

NAND2xp5_ASAP7_75t_L g11007 ( 
.A(n_10409),
.B(n_1446),
.Y(n_11007)
);

OAI21x1_ASAP7_75t_L g11008 ( 
.A1(n_10725),
.A2(n_649),
.B(n_650),
.Y(n_11008)
);

AO21x2_ASAP7_75t_L g11009 ( 
.A1(n_10600),
.A2(n_650),
.B(n_651),
.Y(n_11009)
);

NOR2xp33_ASAP7_75t_L g11010 ( 
.A(n_10506),
.B(n_10660),
.Y(n_11010)
);

OAI21x1_ASAP7_75t_L g11011 ( 
.A1(n_10729),
.A2(n_651),
.B(n_652),
.Y(n_11011)
);

INVx1_ASAP7_75t_L g11012 ( 
.A(n_10421),
.Y(n_11012)
);

OAI21x1_ASAP7_75t_L g11013 ( 
.A1(n_10742),
.A2(n_651),
.B(n_652),
.Y(n_11013)
);

OAI21x1_ASAP7_75t_L g11014 ( 
.A1(n_10818),
.A2(n_652),
.B(n_653),
.Y(n_11014)
);

BUFx6f_ASAP7_75t_L g11015 ( 
.A(n_10644),
.Y(n_11015)
);

INVx1_ASAP7_75t_L g11016 ( 
.A(n_10419),
.Y(n_11016)
);

INVx2_ASAP7_75t_L g11017 ( 
.A(n_10378),
.Y(n_11017)
);

OA21x2_ASAP7_75t_L g11018 ( 
.A1(n_10445),
.A2(n_653),
.B(n_654),
.Y(n_11018)
);

INVx4_ASAP7_75t_L g11019 ( 
.A(n_10644),
.Y(n_11019)
);

BUFx12f_ASAP7_75t_L g11020 ( 
.A(n_10775),
.Y(n_11020)
);

NOR2xp33_ASAP7_75t_L g11021 ( 
.A(n_10661),
.B(n_1447),
.Y(n_11021)
);

OAI21x1_ASAP7_75t_SL g11022 ( 
.A1(n_10700),
.A2(n_653),
.B(n_654),
.Y(n_11022)
);

AO21x2_ASAP7_75t_L g11023 ( 
.A1(n_10551),
.A2(n_654),
.B(n_655),
.Y(n_11023)
);

NOR2xp33_ASAP7_75t_L g11024 ( 
.A(n_10769),
.B(n_1447),
.Y(n_11024)
);

HB1xp67_ASAP7_75t_L g11025 ( 
.A(n_10455),
.Y(n_11025)
);

INVx1_ASAP7_75t_L g11026 ( 
.A(n_10468),
.Y(n_11026)
);

OAI21x1_ASAP7_75t_L g11027 ( 
.A1(n_10827),
.A2(n_655),
.B(n_656),
.Y(n_11027)
);

NAND2xp5_ASAP7_75t_L g11028 ( 
.A(n_10579),
.B(n_1448),
.Y(n_11028)
);

INVx1_ASAP7_75t_L g11029 ( 
.A(n_10541),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_10555),
.Y(n_11030)
);

INVx1_ASAP7_75t_L g11031 ( 
.A(n_10544),
.Y(n_11031)
);

NAND2xp5_ASAP7_75t_L g11032 ( 
.A(n_10565),
.B(n_1448),
.Y(n_11032)
);

INVx1_ASAP7_75t_L g11033 ( 
.A(n_10476),
.Y(n_11033)
);

INVx3_ASAP7_75t_L g11034 ( 
.A(n_10614),
.Y(n_11034)
);

OAI21x1_ASAP7_75t_L g11035 ( 
.A1(n_10628),
.A2(n_655),
.B(n_656),
.Y(n_11035)
);

NAND2x1p5_ASAP7_75t_L g11036 ( 
.A(n_10790),
.B(n_1449),
.Y(n_11036)
);

INVx2_ASAP7_75t_L g11037 ( 
.A(n_10446),
.Y(n_11037)
);

INVx2_ASAP7_75t_SL g11038 ( 
.A(n_10684),
.Y(n_11038)
);

AOI21x1_ASAP7_75t_L g11039 ( 
.A1(n_10732),
.A2(n_656),
.B(n_657),
.Y(n_11039)
);

OAI21x1_ASAP7_75t_L g11040 ( 
.A1(n_10819),
.A2(n_657),
.B(n_658),
.Y(n_11040)
);

AND2x4_ASAP7_75t_L g11041 ( 
.A(n_10704),
.B(n_1449),
.Y(n_11041)
);

AND2x2_ASAP7_75t_L g11042 ( 
.A(n_10697),
.B(n_658),
.Y(n_11042)
);

OR2x2_ASAP7_75t_L g11043 ( 
.A(n_10422),
.B(n_658),
.Y(n_11043)
);

OAI22xp5_ASAP7_75t_L g11044 ( 
.A1(n_10387),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_11044)
);

INVx2_ASAP7_75t_L g11045 ( 
.A(n_10521),
.Y(n_11045)
);

INVxp67_ASAP7_75t_SL g11046 ( 
.A(n_10479),
.Y(n_11046)
);

OAI21x1_ASAP7_75t_L g11047 ( 
.A1(n_10498),
.A2(n_659),
.B(n_660),
.Y(n_11047)
);

INVx2_ASAP7_75t_L g11048 ( 
.A(n_10557),
.Y(n_11048)
);

AOI21xp5_ASAP7_75t_L g11049 ( 
.A1(n_10516),
.A2(n_659),
.B(n_660),
.Y(n_11049)
);

OAI21x1_ASAP7_75t_L g11050 ( 
.A1(n_10518),
.A2(n_661),
.B(n_662),
.Y(n_11050)
);

BUFx2_ASAP7_75t_L g11051 ( 
.A(n_10817),
.Y(n_11051)
);

AOI21x1_ASAP7_75t_L g11052 ( 
.A1(n_10412),
.A2(n_10711),
.B(n_10542),
.Y(n_11052)
);

BUFx6f_ASAP7_75t_L g11053 ( 
.A(n_10684),
.Y(n_11053)
);

AND2x4_ASAP7_75t_SL g11054 ( 
.A(n_10778),
.B(n_1450),
.Y(n_11054)
);

CKINVDCx11_ASAP7_75t_R g11055 ( 
.A(n_10770),
.Y(n_11055)
);

INVx3_ASAP7_75t_SL g11056 ( 
.A(n_10709),
.Y(n_11056)
);

OAI21x1_ASAP7_75t_L g11057 ( 
.A1(n_10523),
.A2(n_661),
.B(n_662),
.Y(n_11057)
);

AOI21xp33_ASAP7_75t_L g11058 ( 
.A1(n_10392),
.A2(n_10391),
.B(n_10405),
.Y(n_11058)
);

BUFx6f_ASAP7_75t_L g11059 ( 
.A(n_10770),
.Y(n_11059)
);

AO21x2_ASAP7_75t_L g11060 ( 
.A1(n_10804),
.A2(n_663),
.B(n_664),
.Y(n_11060)
);

OAI21x1_ASAP7_75t_L g11061 ( 
.A1(n_10532),
.A2(n_663),
.B(n_664),
.Y(n_11061)
);

OA21x2_ASAP7_75t_L g11062 ( 
.A1(n_10442),
.A2(n_663),
.B(n_664),
.Y(n_11062)
);

NOR3xp33_ASAP7_75t_L g11063 ( 
.A(n_10731),
.B(n_1452),
.C(n_1451),
.Y(n_11063)
);

NOR2x1_ASAP7_75t_SL g11064 ( 
.A(n_10471),
.B(n_665),
.Y(n_11064)
);

BUFx2_ASAP7_75t_R g11065 ( 
.A(n_10553),
.Y(n_11065)
);

AO21x2_ASAP7_75t_L g11066 ( 
.A1(n_10472),
.A2(n_665),
.B(n_666),
.Y(n_11066)
);

INVx1_ASAP7_75t_L g11067 ( 
.A(n_10480),
.Y(n_11067)
);

INVx1_ASAP7_75t_L g11068 ( 
.A(n_10490),
.Y(n_11068)
);

INVxp67_ASAP7_75t_SL g11069 ( 
.A(n_10431),
.Y(n_11069)
);

BUFx3_ASAP7_75t_L g11070 ( 
.A(n_10461),
.Y(n_11070)
);

AO21x2_ASAP7_75t_L g11071 ( 
.A1(n_10701),
.A2(n_665),
.B(n_666),
.Y(n_11071)
);

OAI21x1_ASAP7_75t_L g11072 ( 
.A1(n_10543),
.A2(n_666),
.B(n_667),
.Y(n_11072)
);

BUFx12f_ASAP7_75t_L g11073 ( 
.A(n_10531),
.Y(n_11073)
);

INVx1_ASAP7_75t_L g11074 ( 
.A(n_10415),
.Y(n_11074)
);

INVx3_ASAP7_75t_L g11075 ( 
.A(n_10841),
.Y(n_11075)
);

OAI21x1_ASAP7_75t_L g11076 ( 
.A1(n_10546),
.A2(n_667),
.B(n_668),
.Y(n_11076)
);

INVx1_ASAP7_75t_L g11077 ( 
.A(n_10511),
.Y(n_11077)
);

NOR2xp33_ASAP7_75t_L g11078 ( 
.A(n_10682),
.B(n_1451),
.Y(n_11078)
);

AOI22x1_ASAP7_75t_L g11079 ( 
.A1(n_10478),
.A2(n_670),
.B1(n_668),
.B2(n_669),
.Y(n_11079)
);

OA21x2_ASAP7_75t_L g11080 ( 
.A1(n_10448),
.A2(n_669),
.B(n_671),
.Y(n_11080)
);

INVx2_ASAP7_75t_SL g11081 ( 
.A(n_10841),
.Y(n_11081)
);

OAI22xp5_ASAP7_75t_L g11082 ( 
.A1(n_10587),
.A2(n_672),
.B1(n_669),
.B2(n_671),
.Y(n_11082)
);

NAND2x1p5_ASAP7_75t_L g11083 ( 
.A(n_10833),
.B(n_1452),
.Y(n_11083)
);

AOI22xp33_ASAP7_75t_L g11084 ( 
.A1(n_10678),
.A2(n_10768),
.B1(n_10609),
.B2(n_10607),
.Y(n_11084)
);

AO21x2_ASAP7_75t_L g11085 ( 
.A1(n_10549),
.A2(n_672),
.B(n_673),
.Y(n_11085)
);

INVx2_ASAP7_75t_L g11086 ( 
.A(n_10447),
.Y(n_11086)
);

INVx2_ASAP7_75t_SL g11087 ( 
.A(n_10588),
.Y(n_11087)
);

INVx1_ASAP7_75t_L g11088 ( 
.A(n_10481),
.Y(n_11088)
);

A2O1A1Ixp33_ASAP7_75t_L g11089 ( 
.A1(n_10502),
.A2(n_1454),
.B(n_1455),
.C(n_1453),
.Y(n_11089)
);

NAND2xp5_ASAP7_75t_L g11090 ( 
.A(n_10545),
.B(n_1455),
.Y(n_11090)
);

AOI21x1_ASAP7_75t_L g11091 ( 
.A1(n_10608),
.A2(n_672),
.B(n_673),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10535),
.Y(n_11092)
);

BUFx8_ASAP7_75t_L g11093 ( 
.A(n_10823),
.Y(n_11093)
);

AO21x1_ASAP7_75t_L g11094 ( 
.A1(n_10377),
.A2(n_673),
.B(n_674),
.Y(n_11094)
);

CKINVDCx20_ASAP7_75t_R g11095 ( 
.A(n_10683),
.Y(n_11095)
);

OAI221xp5_ASAP7_75t_L g11096 ( 
.A1(n_10444),
.A2(n_676),
.B1(n_674),
.B2(n_675),
.C(n_677),
.Y(n_11096)
);

AO21x2_ASAP7_75t_L g11097 ( 
.A1(n_10508),
.A2(n_675),
.B(n_676),
.Y(n_11097)
);

NAND2xp5_ASAP7_75t_SL g11098 ( 
.A(n_10469),
.B(n_1456),
.Y(n_11098)
);

NAND3xp33_ASAP7_75t_L g11099 ( 
.A(n_10724),
.B(n_10577),
.C(n_10570),
.Y(n_11099)
);

BUFx6f_ASAP7_75t_L g11100 ( 
.A(n_10622),
.Y(n_11100)
);

AOI22xp5_ASAP7_75t_L g11101 ( 
.A1(n_10649),
.A2(n_1457),
.B1(n_1458),
.B2(n_1456),
.Y(n_11101)
);

INVx2_ASAP7_75t_L g11102 ( 
.A(n_10515),
.Y(n_11102)
);

INVx6_ASAP7_75t_L g11103 ( 
.A(n_10690),
.Y(n_11103)
);

OAI21x1_ASAP7_75t_SL g11104 ( 
.A1(n_10612),
.A2(n_675),
.B(n_677),
.Y(n_11104)
);

OAI21x1_ASAP7_75t_SL g11105 ( 
.A1(n_10394),
.A2(n_677),
.B(n_678),
.Y(n_11105)
);

OAI21x1_ASAP7_75t_L g11106 ( 
.A1(n_10558),
.A2(n_678),
.B(n_679),
.Y(n_11106)
);

INVx1_ASAP7_75t_L g11107 ( 
.A(n_10663),
.Y(n_11107)
);

OAI21x1_ASAP7_75t_L g11108 ( 
.A1(n_10562),
.A2(n_678),
.B(n_679),
.Y(n_11108)
);

OAI21x1_ASAP7_75t_L g11109 ( 
.A1(n_10578),
.A2(n_679),
.B(n_680),
.Y(n_11109)
);

OAI21xp5_ASAP7_75t_L g11110 ( 
.A1(n_10581),
.A2(n_1459),
.B(n_1457),
.Y(n_11110)
);

INVx1_ASAP7_75t_L g11111 ( 
.A(n_10740),
.Y(n_11111)
);

INVx1_ASAP7_75t_L g11112 ( 
.A(n_10519),
.Y(n_11112)
);

OAI21x1_ASAP7_75t_SL g11113 ( 
.A1(n_10382),
.A2(n_681),
.B(n_682),
.Y(n_11113)
);

OAI21x1_ASAP7_75t_L g11114 ( 
.A1(n_10596),
.A2(n_681),
.B(n_682),
.Y(n_11114)
);

NAND3xp33_ASAP7_75t_L g11115 ( 
.A(n_10586),
.B(n_1460),
.C(n_1459),
.Y(n_11115)
);

OAI21x1_ASAP7_75t_L g11116 ( 
.A1(n_10602),
.A2(n_683),
.B(n_684),
.Y(n_11116)
);

AND2x4_ASAP7_75t_L g11117 ( 
.A(n_10574),
.B(n_1460),
.Y(n_11117)
);

CKINVDCx11_ASAP7_75t_R g11118 ( 
.A(n_10826),
.Y(n_11118)
);

AO21x2_ASAP7_75t_L g11119 ( 
.A1(n_10537),
.A2(n_683),
.B(n_684),
.Y(n_11119)
);

CKINVDCx8_ASAP7_75t_R g11120 ( 
.A(n_10536),
.Y(n_11120)
);

NAND2xp33_ASAP7_75t_R g11121 ( 
.A(n_10552),
.B(n_685),
.Y(n_11121)
);

OAI21xp5_ASAP7_75t_L g11122 ( 
.A1(n_10413),
.A2(n_1462),
.B(n_1461),
.Y(n_11122)
);

BUFx12f_ASAP7_75t_L g11123 ( 
.A(n_10563),
.Y(n_11123)
);

NAND2xp5_ASAP7_75t_L g11124 ( 
.A(n_10843),
.B(n_1461),
.Y(n_11124)
);

AND2x2_ASAP7_75t_L g11125 ( 
.A(n_10556),
.B(n_685),
.Y(n_11125)
);

INVx1_ASAP7_75t_SL g11126 ( 
.A(n_10811),
.Y(n_11126)
);

AND2x4_ASAP7_75t_L g11127 ( 
.A(n_10735),
.B(n_1462),
.Y(n_11127)
);

CKINVDCx14_ASAP7_75t_R g11128 ( 
.A(n_10767),
.Y(n_11128)
);

AOI22x1_ASAP7_75t_L g11129 ( 
.A1(n_10803),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.Y(n_11129)
);

BUFx6f_ASAP7_75t_L g11130 ( 
.A(n_10720),
.Y(n_11130)
);

INVxp67_ASAP7_75t_SL g11131 ( 
.A(n_10832),
.Y(n_11131)
);

OR2x6_ASAP7_75t_L g11132 ( 
.A(n_10801),
.B(n_1463),
.Y(n_11132)
);

NOR2xp33_ASAP7_75t_L g11133 ( 
.A(n_10673),
.B(n_1463),
.Y(n_11133)
);

INVx8_ASAP7_75t_L g11134 ( 
.A(n_10699),
.Y(n_11134)
);

OAI21x1_ASAP7_75t_L g11135 ( 
.A1(n_10606),
.A2(n_686),
.B(n_687),
.Y(n_11135)
);

NOR2xp33_ASAP7_75t_SL g11136 ( 
.A(n_10715),
.B(n_1465),
.Y(n_11136)
);

OAI21x1_ASAP7_75t_L g11137 ( 
.A1(n_10621),
.A2(n_686),
.B(n_687),
.Y(n_11137)
);

NAND2x1p5_ASAP7_75t_L g11138 ( 
.A(n_10719),
.B(n_1465),
.Y(n_11138)
);

OAI21xp5_ASAP7_75t_L g11139 ( 
.A1(n_10443),
.A2(n_1467),
.B(n_1466),
.Y(n_11139)
);

AND2x4_ASAP7_75t_L g11140 ( 
.A(n_10820),
.B(n_10625),
.Y(n_11140)
);

OAI21x1_ASAP7_75t_L g11141 ( 
.A1(n_10631),
.A2(n_688),
.B(n_689),
.Y(n_11141)
);

HB1xp67_ASAP7_75t_L g11142 ( 
.A(n_10597),
.Y(n_11142)
);

HB1xp67_ASAP7_75t_L g11143 ( 
.A(n_10597),
.Y(n_11143)
);

OAI21xp5_ASAP7_75t_L g11144 ( 
.A1(n_10452),
.A2(n_1467),
.B(n_1466),
.Y(n_11144)
);

OR2x6_ASAP7_75t_L g11145 ( 
.A(n_10509),
.B(n_1468),
.Y(n_11145)
);

HB1xp67_ASAP7_75t_L g11146 ( 
.A(n_10575),
.Y(n_11146)
);

INVx4_ASAP7_75t_L g11147 ( 
.A(n_10634),
.Y(n_11147)
);

OAI22xp33_ASAP7_75t_L g11148 ( 
.A1(n_10675),
.A2(n_1469),
.B1(n_1470),
.B2(n_1468),
.Y(n_11148)
);

BUFx6f_ASAP7_75t_L g11149 ( 
.A(n_10798),
.Y(n_11149)
);

OAI21x1_ASAP7_75t_L g11150 ( 
.A1(n_10632),
.A2(n_688),
.B(n_689),
.Y(n_11150)
);

OAI21x1_ASAP7_75t_L g11151 ( 
.A1(n_10641),
.A2(n_689),
.B(n_690),
.Y(n_11151)
);

AOI22xp5_ASAP7_75t_L g11152 ( 
.A1(n_10441),
.A2(n_1471),
.B1(n_1472),
.B2(n_1470),
.Y(n_11152)
);

INVx1_ASAP7_75t_L g11153 ( 
.A(n_10575),
.Y(n_11153)
);

OA21x2_ASAP7_75t_L g11154 ( 
.A1(n_10794),
.A2(n_690),
.B(n_691),
.Y(n_11154)
);

INVx2_ASAP7_75t_L g11155 ( 
.A(n_10652),
.Y(n_11155)
);

NAND2xp33_ASAP7_75t_L g11156 ( 
.A(n_10603),
.B(n_10635),
.Y(n_11156)
);

OAI21x1_ASAP7_75t_L g11157 ( 
.A1(n_10655),
.A2(n_690),
.B(n_691),
.Y(n_11157)
);

INVx1_ASAP7_75t_L g11158 ( 
.A(n_10438),
.Y(n_11158)
);

AO21x2_ASAP7_75t_L g11159 ( 
.A1(n_10459),
.A2(n_691),
.B(n_692),
.Y(n_11159)
);

INVxp67_ASAP7_75t_SL g11160 ( 
.A(n_10759),
.Y(n_11160)
);

OR2x2_ASAP7_75t_L g11161 ( 
.A(n_10653),
.B(n_692),
.Y(n_11161)
);

NAND2x1p5_ASAP7_75t_L g11162 ( 
.A(n_10659),
.B(n_1471),
.Y(n_11162)
);

CKINVDCx20_ASAP7_75t_R g11163 ( 
.A(n_10687),
.Y(n_11163)
);

OAI21x1_ASAP7_75t_L g11164 ( 
.A1(n_10664),
.A2(n_692),
.B(n_693),
.Y(n_11164)
);

AOI22x1_ASAP7_75t_L g11165 ( 
.A1(n_10611),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.Y(n_11165)
);

OAI21xp5_ASAP7_75t_L g11166 ( 
.A1(n_10464),
.A2(n_10638),
.B(n_10629),
.Y(n_11166)
);

BUFx3_ASAP7_75t_L g11167 ( 
.A(n_10836),
.Y(n_11167)
);

AO21x2_ASAP7_75t_L g11168 ( 
.A1(n_10491),
.A2(n_693),
.B(n_694),
.Y(n_11168)
);

AO21x2_ASAP7_75t_L g11169 ( 
.A1(n_10693),
.A2(n_694),
.B(n_695),
.Y(n_11169)
);

INVx2_ASAP7_75t_L g11170 ( 
.A(n_10688),
.Y(n_11170)
);

OAI21x1_ASAP7_75t_L g11171 ( 
.A1(n_10698),
.A2(n_695),
.B(n_696),
.Y(n_11171)
);

INVx1_ASAP7_75t_L g11172 ( 
.A(n_10438),
.Y(n_11172)
);

BUFx5_ASAP7_75t_L g11173 ( 
.A(n_10812),
.Y(n_11173)
);

NAND2x1p5_ASAP7_75t_L g11174 ( 
.A(n_10620),
.B(n_1472),
.Y(n_11174)
);

OAI21x1_ASAP7_75t_L g11175 ( 
.A1(n_10840),
.A2(n_696),
.B(n_697),
.Y(n_11175)
);

HB1xp67_ASAP7_75t_L g11176 ( 
.A(n_10496),
.Y(n_11176)
);

AO21x1_ASAP7_75t_L g11177 ( 
.A1(n_10702),
.A2(n_10669),
.B(n_10830),
.Y(n_11177)
);

AOI21xp5_ASAP7_75t_L g11178 ( 
.A1(n_10493),
.A2(n_697),
.B(n_698),
.Y(n_11178)
);

OA21x2_ASAP7_75t_L g11179 ( 
.A1(n_10593),
.A2(n_697),
.B(n_698),
.Y(n_11179)
);

INVx1_ASAP7_75t_L g11180 ( 
.A(n_10496),
.Y(n_11180)
);

CKINVDCx20_ASAP7_75t_R g11181 ( 
.A(n_10667),
.Y(n_11181)
);

INVx1_ASAP7_75t_L g11182 ( 
.A(n_10527),
.Y(n_11182)
);

INVx4_ASAP7_75t_L g11183 ( 
.A(n_10488),
.Y(n_11183)
);

OAI21x1_ASAP7_75t_L g11184 ( 
.A1(n_10696),
.A2(n_698),
.B(n_699),
.Y(n_11184)
);

INVx1_ASAP7_75t_L g11185 ( 
.A(n_10695),
.Y(n_11185)
);

CKINVDCx20_ASAP7_75t_R g11186 ( 
.A(n_10677),
.Y(n_11186)
);

OAI21x1_ASAP7_75t_L g11187 ( 
.A1(n_10636),
.A2(n_699),
.B(n_700),
.Y(n_11187)
);

BUFx3_ASAP7_75t_L g11188 ( 
.A(n_10686),
.Y(n_11188)
);

OAI21x1_ASAP7_75t_L g11189 ( 
.A1(n_10681),
.A2(n_10692),
.B(n_10685),
.Y(n_11189)
);

AO21x2_ASAP7_75t_L g11190 ( 
.A1(n_10694),
.A2(n_10776),
.B(n_10741),
.Y(n_11190)
);

AO21x2_ASAP7_75t_L g11191 ( 
.A1(n_10751),
.A2(n_699),
.B(n_700),
.Y(n_11191)
);

OAI21x1_ASAP7_75t_L g11192 ( 
.A1(n_10651),
.A2(n_700),
.B(n_701),
.Y(n_11192)
);

INVx1_ASAP7_75t_L g11193 ( 
.A(n_10695),
.Y(n_11193)
);

BUFx6f_ASAP7_75t_L g11194 ( 
.A(n_10703),
.Y(n_11194)
);

INVx1_ASAP7_75t_L g11195 ( 
.A(n_10547),
.Y(n_11195)
);

OR2x2_ASAP7_75t_L g11196 ( 
.A(n_10646),
.B(n_702),
.Y(n_11196)
);

AO21x2_ASAP7_75t_L g11197 ( 
.A1(n_10762),
.A2(n_702),
.B(n_703),
.Y(n_11197)
);

INVx2_ASAP7_75t_L g11198 ( 
.A(n_10844),
.Y(n_11198)
);

OA21x2_ASAP7_75t_L g11199 ( 
.A1(n_10484),
.A2(n_702),
.B(n_703),
.Y(n_11199)
);

INVx2_ASAP7_75t_L g11200 ( 
.A(n_10705),
.Y(n_11200)
);

OAI21x1_ASAP7_75t_L g11201 ( 
.A1(n_10707),
.A2(n_10746),
.B(n_10737),
.Y(n_11201)
);

INVx1_ASAP7_75t_L g11202 ( 
.A(n_10640),
.Y(n_11202)
);

AO21x2_ASAP7_75t_L g11203 ( 
.A1(n_11160),
.A2(n_10400),
.B(n_10418),
.Y(n_11203)
);

INVx1_ASAP7_75t_L g11204 ( 
.A(n_10862),
.Y(n_11204)
);

INVx1_ASAP7_75t_L g11205 ( 
.A(n_10865),
.Y(n_11205)
);

NAND2xp5_ASAP7_75t_L g11206 ( 
.A(n_11046),
.B(n_10712),
.Y(n_11206)
);

OA21x2_ASAP7_75t_L g11207 ( 
.A1(n_10858),
.A2(n_10665),
.B(n_10744),
.Y(n_11207)
);

OAI21x1_ASAP7_75t_L g11208 ( 
.A1(n_10944),
.A2(n_10845),
.B(n_10748),
.Y(n_11208)
);

OA21x2_ASAP7_75t_L g11209 ( 
.A1(n_10955),
.A2(n_10757),
.B(n_10749),
.Y(n_11209)
);

NAND2x1p5_ASAP7_75t_L g11210 ( 
.A(n_10851),
.B(n_10590),
.Y(n_11210)
);

NOR2xp67_ASAP7_75t_L g11211 ( 
.A(n_11183),
.B(n_10758),
.Y(n_11211)
);

AOI21xp33_ASAP7_75t_SL g11212 ( 
.A1(n_10936),
.A2(n_11056),
.B(n_11138),
.Y(n_11212)
);

OAI21x1_ASAP7_75t_L g11213 ( 
.A1(n_10953),
.A2(n_10676),
.B(n_10589),
.Y(n_11213)
);

AOI21xp5_ASAP7_75t_L g11214 ( 
.A1(n_10915),
.A2(n_11166),
.B(n_11058),
.Y(n_11214)
);

AOI22xp33_ASAP7_75t_L g11215 ( 
.A1(n_11063),
.A2(n_11177),
.B1(n_11099),
.B2(n_10984),
.Y(n_11215)
);

OAI21x1_ASAP7_75t_SL g11216 ( 
.A1(n_10860),
.A2(n_10666),
.B(n_10728),
.Y(n_11216)
);

INVx1_ASAP7_75t_L g11217 ( 
.A(n_10886),
.Y(n_11217)
);

AND2x2_ASAP7_75t_L g11218 ( 
.A(n_10923),
.B(n_10771),
.Y(n_11218)
);

OAI21x1_ASAP7_75t_L g11219 ( 
.A1(n_10870),
.A2(n_11074),
.B(n_10938),
.Y(n_11219)
);

BUFx2_ASAP7_75t_L g11220 ( 
.A(n_10855),
.Y(n_11220)
);

OAI21xp5_ASAP7_75t_L g11221 ( 
.A1(n_10900),
.A2(n_10642),
.B(n_10385),
.Y(n_11221)
);

OAI21x1_ASAP7_75t_L g11222 ( 
.A1(n_11077),
.A2(n_10706),
.B(n_10524),
.Y(n_11222)
);

OR2x2_ASAP7_75t_L g11223 ( 
.A(n_10871),
.B(n_10772),
.Y(n_11223)
);

NAND2xp5_ASAP7_75t_L g11224 ( 
.A(n_10898),
.B(n_10777),
.Y(n_11224)
);

BUFx2_ASAP7_75t_L g11225 ( 
.A(n_10960),
.Y(n_11225)
);

OAI21x1_ASAP7_75t_L g11226 ( 
.A1(n_11092),
.A2(n_10795),
.B(n_10501),
.Y(n_11226)
);

INVx1_ASAP7_75t_SL g11227 ( 
.A(n_11055),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_10852),
.Y(n_11228)
);

OAI21xp33_ASAP7_75t_L g11229 ( 
.A1(n_11084),
.A2(n_10474),
.B(n_10618),
.Y(n_11229)
);

AND2x4_ASAP7_75t_L g11230 ( 
.A(n_11017),
.B(n_10828),
.Y(n_11230)
);

INVx1_ASAP7_75t_L g11231 ( 
.A(n_10854),
.Y(n_11231)
);

OA21x2_ASAP7_75t_L g11232 ( 
.A1(n_11107),
.A2(n_10781),
.B(n_10779),
.Y(n_11232)
);

OAI21x1_ASAP7_75t_L g11233 ( 
.A1(n_11111),
.A2(n_10393),
.B(n_10424),
.Y(n_11233)
);

OR2x2_ASAP7_75t_L g11234 ( 
.A(n_10889),
.B(n_10782),
.Y(n_11234)
);

BUFx4f_ASAP7_75t_SL g11235 ( 
.A(n_10908),
.Y(n_11235)
);

OAI21x1_ASAP7_75t_L g11236 ( 
.A1(n_11155),
.A2(n_10485),
.B(n_10477),
.Y(n_11236)
);

NAND2xp5_ASAP7_75t_L g11237 ( 
.A(n_10857),
.B(n_10784),
.Y(n_11237)
);

OA21x2_ASAP7_75t_L g11238 ( 
.A1(n_10903),
.A2(n_10797),
.B(n_10792),
.Y(n_11238)
);

OAI21x1_ASAP7_75t_L g11239 ( 
.A1(n_11170),
.A2(n_10499),
.B(n_10548),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_10872),
.B(n_10805),
.Y(n_11240)
);

OAI21x1_ASAP7_75t_L g11241 ( 
.A1(n_10937),
.A2(n_10591),
.B(n_10572),
.Y(n_11241)
);

AOI21x1_ASAP7_75t_L g11242 ( 
.A1(n_11025),
.A2(n_10814),
.B(n_10806),
.Y(n_11242)
);

OAI21x1_ASAP7_75t_L g11243 ( 
.A1(n_11153),
.A2(n_11172),
.B(n_11158),
.Y(n_11243)
);

BUFx2_ASAP7_75t_L g11244 ( 
.A(n_10921),
.Y(n_11244)
);

OAI21x1_ASAP7_75t_L g11245 ( 
.A1(n_11180),
.A2(n_10633),
.B(n_10554),
.Y(n_11245)
);

INVx2_ASAP7_75t_L g11246 ( 
.A(n_10856),
.Y(n_11246)
);

AO21x2_ASAP7_75t_L g11247 ( 
.A1(n_10849),
.A2(n_10671),
.B(n_10837),
.Y(n_11247)
);

OAI21x1_ASAP7_75t_L g11248 ( 
.A1(n_10917),
.A2(n_10595),
.B(n_10799),
.Y(n_11248)
);

INVx1_ASAP7_75t_L g11249 ( 
.A(n_10930),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_L g11250 ( 
.A(n_11069),
.B(n_10465),
.Y(n_11250)
);

OAI21x1_ASAP7_75t_L g11251 ( 
.A1(n_10884),
.A2(n_10717),
.B(n_10835),
.Y(n_11251)
);

NAND2x1p5_ASAP7_75t_L g11252 ( 
.A(n_10922),
.B(n_10787),
.Y(n_11252)
);

OA21x2_ASAP7_75t_L g11253 ( 
.A1(n_10873),
.A2(n_10807),
.B(n_10529),
.Y(n_11253)
);

INVx2_ASAP7_75t_L g11254 ( 
.A(n_10910),
.Y(n_11254)
);

INVx1_ASAP7_75t_L g11255 ( 
.A(n_10933),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_10913),
.Y(n_11256)
);

INVx1_ASAP7_75t_L g11257 ( 
.A(n_10919),
.Y(n_11257)
);

AO21x2_ASAP7_75t_L g11258 ( 
.A1(n_11142),
.A2(n_11146),
.B(n_11143),
.Y(n_11258)
);

AOI21xp5_ASAP7_75t_L g11259 ( 
.A1(n_10965),
.A2(n_11178),
.B(n_11148),
.Y(n_11259)
);

HB1xp67_ASAP7_75t_L g11260 ( 
.A(n_10973),
.Y(n_11260)
);

OR2x2_ASAP7_75t_L g11261 ( 
.A(n_10961),
.B(n_10828),
.Y(n_11261)
);

OAI21x1_ASAP7_75t_L g11262 ( 
.A1(n_11202),
.A2(n_10842),
.B(n_10791),
.Y(n_11262)
);

BUFx2_ASAP7_75t_L g11263 ( 
.A(n_10868),
.Y(n_11263)
);

INVx1_ASAP7_75t_L g11264 ( 
.A(n_10920),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_10934),
.Y(n_11265)
);

OAI21x1_ASAP7_75t_L g11266 ( 
.A1(n_11185),
.A2(n_10800),
.B(n_10789),
.Y(n_11266)
);

OAI21xp5_ASAP7_75t_L g11267 ( 
.A1(n_10859),
.A2(n_11049),
.B(n_11115),
.Y(n_11267)
);

OR2x2_ASAP7_75t_L g11268 ( 
.A(n_10876),
.B(n_10640),
.Y(n_11268)
);

AO31x2_ASAP7_75t_L g11269 ( 
.A1(n_11094),
.A2(n_11193),
.A3(n_10964),
.B(n_11182),
.Y(n_11269)
);

NAND2xp5_ASAP7_75t_L g11270 ( 
.A(n_10994),
.B(n_10689),
.Y(n_11270)
);

OAI21xp5_ASAP7_75t_L g11271 ( 
.A1(n_11156),
.A2(n_10672),
.B(n_10513),
.Y(n_11271)
);

INVx2_ASAP7_75t_L g11272 ( 
.A(n_10943),
.Y(n_11272)
);

AND2x4_ASAP7_75t_L g11273 ( 
.A(n_10893),
.B(n_10689),
.Y(n_11273)
);

BUFx2_ASAP7_75t_L g11274 ( 
.A(n_10866),
.Y(n_11274)
);

INVx2_ASAP7_75t_L g11275 ( 
.A(n_10945),
.Y(n_11275)
);

NAND3xp33_ASAP7_75t_L g11276 ( 
.A(n_10952),
.B(n_10755),
.C(n_10522),
.Y(n_11276)
);

OA21x2_ASAP7_75t_L g11277 ( 
.A1(n_10971),
.A2(n_10887),
.B(n_10948),
.Y(n_11277)
);

AOI21xp5_ASAP7_75t_L g11278 ( 
.A1(n_10980),
.A2(n_10512),
.B(n_10533),
.Y(n_11278)
);

OAI21x1_ASAP7_75t_L g11279 ( 
.A1(n_10881),
.A2(n_10567),
.B(n_10561),
.Y(n_11279)
);

HB1xp67_ASAP7_75t_L g11280 ( 
.A(n_10848),
.Y(n_11280)
);

AOI21xp5_ASAP7_75t_SL g11281 ( 
.A1(n_11064),
.A2(n_10786),
.B(n_10739),
.Y(n_11281)
);

OA21x2_ASAP7_75t_L g11282 ( 
.A1(n_11131),
.A2(n_10888),
.B(n_10853),
.Y(n_11282)
);

AOI22xp33_ASAP7_75t_L g11283 ( 
.A1(n_11190),
.A2(n_10713),
.B1(n_10437),
.B2(n_10389),
.Y(n_11283)
);

OAI21x1_ASAP7_75t_SL g11284 ( 
.A1(n_11052),
.A2(n_10978),
.B(n_10878),
.Y(n_11284)
);

INVx1_ASAP7_75t_L g11285 ( 
.A(n_10967),
.Y(n_11285)
);

HB1xp67_ASAP7_75t_L g11286 ( 
.A(n_11176),
.Y(n_11286)
);

AO31x2_ASAP7_75t_L g11287 ( 
.A1(n_11195),
.A2(n_10808),
.A3(n_10765),
.B(n_10747),
.Y(n_11287)
);

NAND2xp5_ASAP7_75t_L g11288 ( 
.A(n_11026),
.B(n_10788),
.Y(n_11288)
);

AO21x2_ASAP7_75t_L g11289 ( 
.A1(n_11016),
.A2(n_10838),
.B(n_10831),
.Y(n_11289)
);

OA21x2_ASAP7_75t_L g11290 ( 
.A1(n_10942),
.A2(n_10824),
.B(n_10723),
.Y(n_11290)
);

BUFx3_ASAP7_75t_L g11291 ( 
.A(n_10861),
.Y(n_11291)
);

NOR2xp33_ASAP7_75t_L g11292 ( 
.A(n_10883),
.B(n_10834),
.Y(n_11292)
);

AND2x4_ASAP7_75t_L g11293 ( 
.A(n_10885),
.B(n_10788),
.Y(n_11293)
);

BUFx6f_ASAP7_75t_L g11294 ( 
.A(n_10861),
.Y(n_11294)
);

INVx1_ASAP7_75t_L g11295 ( 
.A(n_10882),
.Y(n_11295)
);

AO21x2_ASAP7_75t_L g11296 ( 
.A1(n_11031),
.A2(n_10483),
.B(n_10463),
.Y(n_11296)
);

AO21x2_ASAP7_75t_L g11297 ( 
.A1(n_11033),
.A2(n_10390),
.B(n_10691),
.Y(n_11297)
);

NAND2x1p5_ASAP7_75t_L g11298 ( 
.A(n_10940),
.B(n_10829),
.Y(n_11298)
);

OAI21x1_ASAP7_75t_L g11299 ( 
.A1(n_10847),
.A2(n_10390),
.B(n_10829),
.Y(n_11299)
);

OR2x6_ASAP7_75t_L g11300 ( 
.A(n_10918),
.B(n_10559),
.Y(n_11300)
);

NAND2xp5_ASAP7_75t_L g11301 ( 
.A(n_11067),
.B(n_1473),
.Y(n_11301)
);

INVxp67_ASAP7_75t_L g11302 ( 
.A(n_11018),
.Y(n_11302)
);

AND2x4_ASAP7_75t_L g11303 ( 
.A(n_11045),
.B(n_1473),
.Y(n_11303)
);

AO21x2_ASAP7_75t_L g11304 ( 
.A1(n_11068),
.A2(n_10559),
.B(n_704),
.Y(n_11304)
);

BUFx10_ASAP7_75t_L g11305 ( 
.A(n_11054),
.Y(n_11305)
);

OAI21x1_ASAP7_75t_L g11306 ( 
.A1(n_10850),
.A2(n_704),
.B(n_705),
.Y(n_11306)
);

INVx1_ASAP7_75t_L g11307 ( 
.A(n_10951),
.Y(n_11307)
);

NAND2xp5_ASAP7_75t_SL g11308 ( 
.A(n_11002),
.B(n_1474),
.Y(n_11308)
);

INVx2_ASAP7_75t_L g11309 ( 
.A(n_10891),
.Y(n_11309)
);

CKINVDCx5p33_ASAP7_75t_R g11310 ( 
.A(n_10924),
.Y(n_11310)
);

AO21x2_ASAP7_75t_L g11311 ( 
.A1(n_11088),
.A2(n_704),
.B(n_705),
.Y(n_11311)
);

OAI21x1_ASAP7_75t_L g11312 ( 
.A1(n_10906),
.A2(n_705),
.B(n_706),
.Y(n_11312)
);

INVx2_ASAP7_75t_L g11313 ( 
.A(n_10926),
.Y(n_11313)
);

OAI21x1_ASAP7_75t_L g11314 ( 
.A1(n_10927),
.A2(n_10894),
.B(n_10925),
.Y(n_11314)
);

NAND2xp5_ASAP7_75t_L g11315 ( 
.A(n_11112),
.B(n_11102),
.Y(n_11315)
);

NAND2xp5_ASAP7_75t_L g11316 ( 
.A(n_11029),
.B(n_1474),
.Y(n_11316)
);

BUFx3_ASAP7_75t_L g11317 ( 
.A(n_10939),
.Y(n_11317)
);

AND2x4_ASAP7_75t_L g11318 ( 
.A(n_11048),
.B(n_1475),
.Y(n_11318)
);

OAI21x1_ASAP7_75t_L g11319 ( 
.A1(n_10959),
.A2(n_706),
.B(n_707),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_10992),
.Y(n_11320)
);

OR2x2_ASAP7_75t_L g11321 ( 
.A(n_10962),
.B(n_707),
.Y(n_11321)
);

NAND2xp5_ASAP7_75t_L g11322 ( 
.A(n_11030),
.B(n_1475),
.Y(n_11322)
);

OAI21x1_ASAP7_75t_SL g11323 ( 
.A1(n_11039),
.A2(n_708),
.B(n_709),
.Y(n_11323)
);

AOI22xp5_ASAP7_75t_L g11324 ( 
.A1(n_10969),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_11324)
);

NAND3xp33_ASAP7_75t_L g11325 ( 
.A(n_10911),
.B(n_708),
.C(n_709),
.Y(n_11325)
);

OAI21x1_ASAP7_75t_SL g11326 ( 
.A1(n_10993),
.A2(n_710),
.B(n_711),
.Y(n_11326)
);

OA21x2_ASAP7_75t_L g11327 ( 
.A1(n_10949),
.A2(n_710),
.B(n_712),
.Y(n_11327)
);

BUFx3_ASAP7_75t_L g11328 ( 
.A(n_10863),
.Y(n_11328)
);

NOR2xp33_ASAP7_75t_L g11329 ( 
.A(n_10931),
.B(n_1476),
.Y(n_11329)
);

NAND2xp5_ASAP7_75t_L g11330 ( 
.A(n_11198),
.B(n_1477),
.Y(n_11330)
);

BUFx6f_ASAP7_75t_L g11331 ( 
.A(n_10880),
.Y(n_11331)
);

AO21x2_ASAP7_75t_L g11332 ( 
.A1(n_10972),
.A2(n_10981),
.B(n_10974),
.Y(n_11332)
);

OAI21x1_ASAP7_75t_L g11333 ( 
.A1(n_10864),
.A2(n_712),
.B(n_713),
.Y(n_11333)
);

OAI21x1_ASAP7_75t_L g11334 ( 
.A1(n_10950),
.A2(n_712),
.B(n_713),
.Y(n_11334)
);

NAND2x1p5_ASAP7_75t_L g11335 ( 
.A(n_10941),
.B(n_1477),
.Y(n_11335)
);

OAI21xp5_ASAP7_75t_L g11336 ( 
.A1(n_11110),
.A2(n_11139),
.B(n_11122),
.Y(n_11336)
);

NAND2x1p5_ASAP7_75t_L g11337 ( 
.A(n_10957),
.B(n_1478),
.Y(n_11337)
);

NAND2x1p5_ASAP7_75t_L g11338 ( 
.A(n_10970),
.B(n_1478),
.Y(n_11338)
);

CKINVDCx5p33_ASAP7_75t_R g11339 ( 
.A(n_10905),
.Y(n_11339)
);

OR2x2_ASAP7_75t_L g11340 ( 
.A(n_11012),
.B(n_10989),
.Y(n_11340)
);

INVx2_ASAP7_75t_L g11341 ( 
.A(n_10954),
.Y(n_11341)
);

OA21x2_ASAP7_75t_L g11342 ( 
.A1(n_10995),
.A2(n_714),
.B(n_715),
.Y(n_11342)
);

OAI21x1_ASAP7_75t_L g11343 ( 
.A1(n_11189),
.A2(n_714),
.B(n_715),
.Y(n_11343)
);

OAI21x1_ASAP7_75t_L g11344 ( 
.A1(n_10867),
.A2(n_715),
.B(n_716),
.Y(n_11344)
);

BUFx3_ASAP7_75t_L g11345 ( 
.A(n_11051),
.Y(n_11345)
);

HB1xp67_ASAP7_75t_L g11346 ( 
.A(n_10928),
.Y(n_11346)
);

AOI21x1_ASAP7_75t_L g11347 ( 
.A1(n_11005),
.A2(n_716),
.B(n_717),
.Y(n_11347)
);

OAI21xp33_ASAP7_75t_SL g11348 ( 
.A1(n_11126),
.A2(n_716),
.B(n_718),
.Y(n_11348)
);

INVx2_ASAP7_75t_SL g11349 ( 
.A(n_10947),
.Y(n_11349)
);

OR2x2_ASAP7_75t_L g11350 ( 
.A(n_10998),
.B(n_718),
.Y(n_11350)
);

INVx1_ASAP7_75t_L g11351 ( 
.A(n_11000),
.Y(n_11351)
);

CKINVDCx20_ASAP7_75t_R g11352 ( 
.A(n_11095),
.Y(n_11352)
);

OAI21x1_ASAP7_75t_L g11353 ( 
.A1(n_11006),
.A2(n_719),
.B(n_720),
.Y(n_11353)
);

NAND2x1p5_ASAP7_75t_L g11354 ( 
.A(n_11034),
.B(n_1479),
.Y(n_11354)
);

NAND2x1p5_ASAP7_75t_L g11355 ( 
.A(n_11147),
.B(n_1479),
.Y(n_11355)
);

OA21x2_ASAP7_75t_L g11356 ( 
.A1(n_10899),
.A2(n_719),
.B(n_720),
.Y(n_11356)
);

BUFx2_ASAP7_75t_L g11357 ( 
.A(n_11173),
.Y(n_11357)
);

OAI21xp5_ASAP7_75t_L g11358 ( 
.A1(n_11144),
.A2(n_10890),
.B(n_11201),
.Y(n_11358)
);

NOR2xp33_ASAP7_75t_L g11359 ( 
.A(n_10911),
.B(n_1480),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_10907),
.Y(n_11360)
);

AOI21xp5_ASAP7_75t_L g11361 ( 
.A1(n_10979),
.A2(n_1481),
.B(n_1480),
.Y(n_11361)
);

AND2x2_ASAP7_75t_L g11362 ( 
.A(n_11037),
.B(n_719),
.Y(n_11362)
);

NAND2xp5_ASAP7_75t_L g11363 ( 
.A(n_11200),
.B(n_1482),
.Y(n_11363)
);

NOR2xp33_ASAP7_75t_L g11364 ( 
.A(n_11194),
.B(n_1482),
.Y(n_11364)
);

NAND2xp5_ASAP7_75t_L g11365 ( 
.A(n_10869),
.B(n_1483),
.Y(n_11365)
);

NOR2xp67_ASAP7_75t_L g11366 ( 
.A(n_10875),
.B(n_720),
.Y(n_11366)
);

INVx1_ASAP7_75t_SL g11367 ( 
.A(n_10902),
.Y(n_11367)
);

OAI21x1_ASAP7_75t_SL g11368 ( 
.A1(n_11022),
.A2(n_721),
.B(n_722),
.Y(n_11368)
);

AND2x2_ASAP7_75t_L g11369 ( 
.A(n_11086),
.B(n_721),
.Y(n_11369)
);

NAND2xp5_ASAP7_75t_L g11370 ( 
.A(n_10904),
.B(n_1484),
.Y(n_11370)
);

AO31x2_ASAP7_75t_L g11371 ( 
.A1(n_11024),
.A2(n_723),
.A3(n_721),
.B(n_722),
.Y(n_11371)
);

OAI21x1_ASAP7_75t_L g11372 ( 
.A1(n_10990),
.A2(n_722),
.B(n_723),
.Y(n_11372)
);

INVx1_ASAP7_75t_L g11373 ( 
.A(n_11140),
.Y(n_11373)
);

OAI21x1_ASAP7_75t_L g11374 ( 
.A1(n_10963),
.A2(n_723),
.B(n_724),
.Y(n_11374)
);

INVx2_ASAP7_75t_L g11375 ( 
.A(n_11173),
.Y(n_11375)
);

AOI21x1_ASAP7_75t_L g11376 ( 
.A1(n_10968),
.A2(n_724),
.B(n_725),
.Y(n_11376)
);

INVx1_ASAP7_75t_L g11377 ( 
.A(n_10877),
.Y(n_11377)
);

OAI21x1_ASAP7_75t_L g11378 ( 
.A1(n_10966),
.A2(n_724),
.B(n_725),
.Y(n_11378)
);

OAI21x1_ASAP7_75t_SL g11379 ( 
.A1(n_10987),
.A2(n_726),
.B(n_727),
.Y(n_11379)
);

NAND2xp5_ASAP7_75t_L g11380 ( 
.A(n_11188),
.B(n_1484),
.Y(n_11380)
);

NAND2xp5_ASAP7_75t_L g11381 ( 
.A(n_11194),
.B(n_1485),
.Y(n_11381)
);

AO31x2_ASAP7_75t_L g11382 ( 
.A1(n_10958),
.A2(n_728),
.A3(n_726),
.B(n_727),
.Y(n_11382)
);

INVx2_ASAP7_75t_L g11383 ( 
.A(n_11173),
.Y(n_11383)
);

OAI21x1_ASAP7_75t_L g11384 ( 
.A1(n_11014),
.A2(n_726),
.B(n_727),
.Y(n_11384)
);

NAND2x1p5_ASAP7_75t_L g11385 ( 
.A(n_10874),
.B(n_1486),
.Y(n_11385)
);

BUFx6f_ASAP7_75t_L g11386 ( 
.A(n_10880),
.Y(n_11386)
);

HB1xp67_ASAP7_75t_L g11387 ( 
.A(n_10946),
.Y(n_11387)
);

AOI21xp5_ASAP7_75t_L g11388 ( 
.A1(n_11089),
.A2(n_1487),
.B(n_1486),
.Y(n_11388)
);

NAND3xp33_ASAP7_75t_L g11389 ( 
.A(n_11165),
.B(n_10986),
.C(n_10879),
.Y(n_11389)
);

OAI21x1_ASAP7_75t_L g11390 ( 
.A1(n_11027),
.A2(n_728),
.B(n_729),
.Y(n_11390)
);

INVx1_ASAP7_75t_L g11391 ( 
.A(n_11062),
.Y(n_11391)
);

INVx2_ASAP7_75t_L g11392 ( 
.A(n_10929),
.Y(n_11392)
);

NAND2x1p5_ASAP7_75t_L g11393 ( 
.A(n_11149),
.B(n_1487),
.Y(n_11393)
);

NAND2xp5_ASAP7_75t_L g11394 ( 
.A(n_10897),
.B(n_1488),
.Y(n_11394)
);

BUFx2_ASAP7_75t_L g11395 ( 
.A(n_11123),
.Y(n_11395)
);

AO31x2_ASAP7_75t_L g11396 ( 
.A1(n_10985),
.A2(n_730),
.A3(n_728),
.B(n_729),
.Y(n_11396)
);

OAI21xp33_ASAP7_75t_SL g11397 ( 
.A1(n_10991),
.A2(n_729),
.B(n_730),
.Y(n_11397)
);

AO21x2_ASAP7_75t_L g11398 ( 
.A1(n_11066),
.A2(n_730),
.B(n_731),
.Y(n_11398)
);

NAND2x1p5_ASAP7_75t_L g11399 ( 
.A(n_11149),
.B(n_1488),
.Y(n_11399)
);

OAI21x1_ASAP7_75t_L g11400 ( 
.A1(n_11035),
.A2(n_731),
.B(n_732),
.Y(n_11400)
);

CKINVDCx5p33_ASAP7_75t_R g11401 ( 
.A(n_11118),
.Y(n_11401)
);

BUFx2_ASAP7_75t_L g11402 ( 
.A(n_11130),
.Y(n_11402)
);

INVx2_ASAP7_75t_L g11403 ( 
.A(n_10932),
.Y(n_11403)
);

INVx1_ASAP7_75t_L g11404 ( 
.A(n_11004),
.Y(n_11404)
);

BUFx6f_ASAP7_75t_L g11405 ( 
.A(n_10912),
.Y(n_11405)
);

INVx2_ASAP7_75t_SL g11406 ( 
.A(n_11134),
.Y(n_11406)
);

OAI21x1_ASAP7_75t_L g11407 ( 
.A1(n_11040),
.A2(n_731),
.B(n_732),
.Y(n_11407)
);

AOI21xp33_ASAP7_75t_SL g11408 ( 
.A1(n_11121),
.A2(n_732),
.B(n_733),
.Y(n_11408)
);

OAI21x1_ASAP7_75t_L g11409 ( 
.A1(n_10975),
.A2(n_733),
.B(n_734),
.Y(n_11409)
);

OAI21x1_ASAP7_75t_L g11410 ( 
.A1(n_10988),
.A2(n_734),
.B(n_735),
.Y(n_11410)
);

BUFx2_ASAP7_75t_L g11411 ( 
.A(n_11130),
.Y(n_11411)
);

AND2x4_ASAP7_75t_L g11412 ( 
.A(n_11075),
.B(n_1489),
.Y(n_11412)
);

NOR2xp33_ASAP7_75t_L g11413 ( 
.A(n_11120),
.B(n_11010),
.Y(n_11413)
);

AND2x4_ASAP7_75t_SL g11414 ( 
.A(n_10935),
.B(n_1490),
.Y(n_11414)
);

AO21x2_ASAP7_75t_L g11415 ( 
.A1(n_11104),
.A2(n_735),
.B(n_736),
.Y(n_11415)
);

OA21x2_ASAP7_75t_L g11416 ( 
.A1(n_10892),
.A2(n_735),
.B(n_736),
.Y(n_11416)
);

INVx1_ASAP7_75t_L g11417 ( 
.A(n_11080),
.Y(n_11417)
);

OAI21xp5_ASAP7_75t_L g11418 ( 
.A1(n_10916),
.A2(n_736),
.B(n_737),
.Y(n_11418)
);

BUFx6f_ASAP7_75t_L g11419 ( 
.A(n_10912),
.Y(n_11419)
);

OAI21xp5_ASAP7_75t_L g11420 ( 
.A1(n_11133),
.A2(n_737),
.B(n_738),
.Y(n_11420)
);

BUFx2_ASAP7_75t_L g11421 ( 
.A(n_11167),
.Y(n_11421)
);

OAI21x1_ASAP7_75t_L g11422 ( 
.A1(n_11047),
.A2(n_738),
.B(n_739),
.Y(n_11422)
);

OA21x2_ASAP7_75t_L g11423 ( 
.A1(n_10956),
.A2(n_738),
.B(n_739),
.Y(n_11423)
);

AO21x2_ASAP7_75t_L g11424 ( 
.A1(n_11001),
.A2(n_739),
.B(n_740),
.Y(n_11424)
);

INVx1_ASAP7_75t_L g11425 ( 
.A(n_11085),
.Y(n_11425)
);

NOR2xp33_ASAP7_75t_L g11426 ( 
.A(n_11028),
.B(n_1490),
.Y(n_11426)
);

INVx2_ASAP7_75t_L g11427 ( 
.A(n_11038),
.Y(n_11427)
);

OAI21x1_ASAP7_75t_L g11428 ( 
.A1(n_11050),
.A2(n_11061),
.B(n_11057),
.Y(n_11428)
);

INVx1_ASAP7_75t_L g11429 ( 
.A(n_11097),
.Y(n_11429)
);

NAND2xp5_ASAP7_75t_L g11430 ( 
.A(n_11119),
.B(n_1491),
.Y(n_11430)
);

INVx2_ASAP7_75t_L g11431 ( 
.A(n_11081),
.Y(n_11431)
);

OA21x2_ASAP7_75t_L g11432 ( 
.A1(n_11090),
.A2(n_11007),
.B(n_11072),
.Y(n_11432)
);

AOI21xp33_ASAP7_75t_SL g11433 ( 
.A1(n_11132),
.A2(n_740),
.B(n_741),
.Y(n_11433)
);

NOR2x1_ASAP7_75t_SL g11434 ( 
.A(n_11020),
.B(n_741),
.Y(n_11434)
);

OAI21x1_ASAP7_75t_L g11435 ( 
.A1(n_11076),
.A2(n_741),
.B(n_742),
.Y(n_11435)
);

OAI21xp5_ASAP7_75t_L g11436 ( 
.A1(n_11032),
.A2(n_742),
.B(n_743),
.Y(n_11436)
);

OR2x2_ASAP7_75t_L g11437 ( 
.A(n_11043),
.B(n_742),
.Y(n_11437)
);

OA21x2_ASAP7_75t_L g11438 ( 
.A1(n_11106),
.A2(n_743),
.B(n_744),
.Y(n_11438)
);

CKINVDCx6p67_ASAP7_75t_R g11439 ( 
.A(n_11145),
.Y(n_11439)
);

INVx1_ASAP7_75t_L g11440 ( 
.A(n_11003),
.Y(n_11440)
);

OAI21x1_ASAP7_75t_L g11441 ( 
.A1(n_11108),
.A2(n_743),
.B(n_744),
.Y(n_11441)
);

OR2x2_ASAP7_75t_L g11442 ( 
.A(n_11161),
.B(n_744),
.Y(n_11442)
);

AOI21x1_ASAP7_75t_L g11443 ( 
.A1(n_11098),
.A2(n_745),
.B(n_746),
.Y(n_11443)
);

AOI22xp33_ASAP7_75t_L g11444 ( 
.A1(n_11159),
.A2(n_1492),
.B1(n_1493),
.B2(n_1491),
.Y(n_11444)
);

AO21x2_ASAP7_75t_L g11445 ( 
.A1(n_11124),
.A2(n_745),
.B(n_746),
.Y(n_11445)
);

OR2x6_ASAP7_75t_L g11446 ( 
.A(n_11134),
.B(n_1492),
.Y(n_11446)
);

NAND2xp5_ASAP7_75t_L g11447 ( 
.A(n_10997),
.B(n_1493),
.Y(n_11447)
);

NAND2xp5_ASAP7_75t_L g11448 ( 
.A(n_11021),
.B(n_1496),
.Y(n_11448)
);

OAI21x1_ASAP7_75t_L g11449 ( 
.A1(n_11109),
.A2(n_746),
.B(n_747),
.Y(n_11449)
);

INVx1_ASAP7_75t_L g11450 ( 
.A(n_11008),
.Y(n_11450)
);

OAI21x1_ASAP7_75t_L g11451 ( 
.A1(n_11114),
.A2(n_747),
.B(n_748),
.Y(n_11451)
);

INVx2_ASAP7_75t_L g11452 ( 
.A(n_11087),
.Y(n_11452)
);

BUFx2_ASAP7_75t_L g11453 ( 
.A(n_11073),
.Y(n_11453)
);

OAI21x1_ASAP7_75t_L g11454 ( 
.A1(n_11116),
.A2(n_748),
.B(n_749),
.Y(n_11454)
);

INVx3_ASAP7_75t_L g11455 ( 
.A(n_11019),
.Y(n_11455)
);

OAI21x1_ASAP7_75t_SL g11456 ( 
.A1(n_11091),
.A2(n_748),
.B(n_749),
.Y(n_11456)
);

OAI21x1_ASAP7_75t_L g11457 ( 
.A1(n_11135),
.A2(n_749),
.B(n_750),
.Y(n_11457)
);

AO21x2_ASAP7_75t_L g11458 ( 
.A1(n_10999),
.A2(n_750),
.B(n_751),
.Y(n_11458)
);

NAND2x1p5_ASAP7_75t_L g11459 ( 
.A(n_11070),
.B(n_1496),
.Y(n_11459)
);

OA21x2_ASAP7_75t_L g11460 ( 
.A1(n_11137),
.A2(n_750),
.B(n_751),
.Y(n_11460)
);

OAI21x1_ASAP7_75t_L g11461 ( 
.A1(n_11141),
.A2(n_751),
.B(n_752),
.Y(n_11461)
);

A2O1A1Ixp33_ASAP7_75t_L g11462 ( 
.A1(n_10977),
.A2(n_754),
.B(n_752),
.C(n_753),
.Y(n_11462)
);

INVx1_ASAP7_75t_L g11463 ( 
.A(n_11011),
.Y(n_11463)
);

OAI21x1_ASAP7_75t_SL g11464 ( 
.A1(n_11105),
.A2(n_753),
.B(n_754),
.Y(n_11464)
);

OAI21x1_ASAP7_75t_L g11465 ( 
.A1(n_11150),
.A2(n_753),
.B(n_754),
.Y(n_11465)
);

OA21x2_ASAP7_75t_L g11466 ( 
.A1(n_11151),
.A2(n_11164),
.B(n_11157),
.Y(n_11466)
);

OA21x2_ASAP7_75t_L g11467 ( 
.A1(n_11171),
.A2(n_755),
.B(n_756),
.Y(n_11467)
);

OAI21x1_ASAP7_75t_L g11468 ( 
.A1(n_11013),
.A2(n_755),
.B(n_756),
.Y(n_11468)
);

AO21x2_ASAP7_75t_L g11469 ( 
.A1(n_11113),
.A2(n_755),
.B(n_757),
.Y(n_11469)
);

AND2x2_ASAP7_75t_L g11470 ( 
.A(n_11128),
.B(n_757),
.Y(n_11470)
);

OAI21x1_ASAP7_75t_L g11471 ( 
.A1(n_11184),
.A2(n_11175),
.B(n_11187),
.Y(n_11471)
);

OA21x2_ASAP7_75t_L g11472 ( 
.A1(n_10901),
.A2(n_757),
.B(n_758),
.Y(n_11472)
);

AO21x2_ASAP7_75t_L g11473 ( 
.A1(n_11168),
.A2(n_758),
.B(n_759),
.Y(n_11473)
);

AND2x2_ASAP7_75t_L g11474 ( 
.A(n_11100),
.B(n_759),
.Y(n_11474)
);

INVx2_ASAP7_75t_L g11475 ( 
.A(n_11100),
.Y(n_11475)
);

OR2x2_ASAP7_75t_L g11476 ( 
.A(n_11196),
.B(n_760),
.Y(n_11476)
);

AOI22xp33_ASAP7_75t_L g11477 ( 
.A1(n_11096),
.A2(n_11197),
.B1(n_11199),
.B2(n_11169),
.Y(n_11477)
);

INVx3_ASAP7_75t_L g11478 ( 
.A(n_11015),
.Y(n_11478)
);

INVx3_ASAP7_75t_L g11479 ( 
.A(n_11015),
.Y(n_11479)
);

NOR2x1_ASAP7_75t_SL g11480 ( 
.A(n_11053),
.B(n_760),
.Y(n_11480)
);

NAND2xp5_ASAP7_75t_L g11481 ( 
.A(n_11078),
.B(n_1497),
.Y(n_11481)
);

AND2x4_ASAP7_75t_L g11482 ( 
.A(n_11053),
.B(n_1497),
.Y(n_11482)
);

OAI21x1_ASAP7_75t_L g11483 ( 
.A1(n_11162),
.A2(n_761),
.B(n_762),
.Y(n_11483)
);

AOI21xp5_ASAP7_75t_L g11484 ( 
.A1(n_11044),
.A2(n_1499),
.B(n_1498),
.Y(n_11484)
);

AND3x2_ASAP7_75t_L g11485 ( 
.A(n_11136),
.B(n_761),
.C(n_762),
.Y(n_11485)
);

A2O1A1Ixp33_ASAP7_75t_L g11486 ( 
.A1(n_10996),
.A2(n_763),
.B(n_761),
.C(n_762),
.Y(n_11486)
);

INVx2_ASAP7_75t_L g11487 ( 
.A(n_11059),
.Y(n_11487)
);

INVx1_ASAP7_75t_L g11488 ( 
.A(n_11154),
.Y(n_11488)
);

AND2x2_ASAP7_75t_L g11489 ( 
.A(n_11059),
.B(n_763),
.Y(n_11489)
);

INVx1_ASAP7_75t_L g11490 ( 
.A(n_10976),
.Y(n_11490)
);

OAI21x1_ASAP7_75t_L g11491 ( 
.A1(n_11174),
.A2(n_764),
.B(n_765),
.Y(n_11491)
);

AO21x2_ASAP7_75t_L g11492 ( 
.A1(n_11042),
.A2(n_764),
.B(n_765),
.Y(n_11492)
);

INVx2_ASAP7_75t_L g11493 ( 
.A(n_11103),
.Y(n_11493)
);

AO31x2_ASAP7_75t_L g11494 ( 
.A1(n_11082),
.A2(n_767),
.A3(n_765),
.B(n_766),
.Y(n_11494)
);

OAI21x1_ASAP7_75t_L g11495 ( 
.A1(n_10914),
.A2(n_766),
.B(n_767),
.Y(n_11495)
);

OAI21x1_ASAP7_75t_L g11496 ( 
.A1(n_11192),
.A2(n_766),
.B(n_767),
.Y(n_11496)
);

AND2x2_ASAP7_75t_L g11497 ( 
.A(n_11125),
.B(n_768),
.Y(n_11497)
);

OA21x2_ASAP7_75t_L g11498 ( 
.A1(n_10895),
.A2(n_10982),
.B(n_11117),
.Y(n_11498)
);

OAI21x1_ASAP7_75t_L g11499 ( 
.A1(n_10909),
.A2(n_768),
.B(n_769),
.Y(n_11499)
);

AND2x4_ASAP7_75t_L g11500 ( 
.A(n_11041),
.B(n_1498),
.Y(n_11500)
);

AOI21x1_ASAP7_75t_L g11501 ( 
.A1(n_11179),
.A2(n_768),
.B(n_769),
.Y(n_11501)
);

INVx1_ASAP7_75t_L g11502 ( 
.A(n_11009),
.Y(n_11502)
);

INVxp67_ASAP7_75t_SL g11503 ( 
.A(n_11093),
.Y(n_11503)
);

AOI21xp5_ASAP7_75t_L g11504 ( 
.A1(n_10896),
.A2(n_1500),
.B(n_1499),
.Y(n_11504)
);

INVx1_ASAP7_75t_L g11505 ( 
.A(n_11023),
.Y(n_11505)
);

AO21x2_ASAP7_75t_L g11506 ( 
.A1(n_11060),
.A2(n_11191),
.B(n_11071),
.Y(n_11506)
);

OAI21x1_ASAP7_75t_L g11507 ( 
.A1(n_11036),
.A2(n_769),
.B(n_770),
.Y(n_11507)
);

OAI21x1_ASAP7_75t_SL g11508 ( 
.A1(n_10983),
.A2(n_770),
.B(n_771),
.Y(n_11508)
);

INVx3_ASAP7_75t_L g11509 ( 
.A(n_11127),
.Y(n_11509)
);

OAI21x1_ASAP7_75t_L g11510 ( 
.A1(n_11083),
.A2(n_770),
.B(n_771),
.Y(n_11510)
);

AO21x2_ASAP7_75t_L g11511 ( 
.A1(n_11101),
.A2(n_11152),
.B(n_11065),
.Y(n_11511)
);

NAND2xp5_ASAP7_75t_L g11512 ( 
.A(n_11186),
.B(n_1500),
.Y(n_11512)
);

OA21x2_ASAP7_75t_L g11513 ( 
.A1(n_11129),
.A2(n_771),
.B(n_772),
.Y(n_11513)
);

INVx3_ASAP7_75t_L g11514 ( 
.A(n_11163),
.Y(n_11514)
);

OAI21x1_ASAP7_75t_L g11515 ( 
.A1(n_11079),
.A2(n_772),
.B(n_773),
.Y(n_11515)
);

OA21x2_ASAP7_75t_L g11516 ( 
.A1(n_11181),
.A2(n_772),
.B(n_773),
.Y(n_11516)
);

OA21x2_ASAP7_75t_L g11517 ( 
.A1(n_10858),
.A2(n_773),
.B(n_774),
.Y(n_11517)
);

INVx1_ASAP7_75t_L g11518 ( 
.A(n_10862),
.Y(n_11518)
);

OAI21x1_ASAP7_75t_L g11519 ( 
.A1(n_10944),
.A2(n_774),
.B(n_775),
.Y(n_11519)
);

AND2x2_ASAP7_75t_L g11520 ( 
.A(n_10923),
.B(n_774),
.Y(n_11520)
);

BUFx12f_ASAP7_75t_L g11521 ( 
.A(n_10861),
.Y(n_11521)
);

NAND2x1p5_ASAP7_75t_L g11522 ( 
.A(n_10851),
.B(n_1501),
.Y(n_11522)
);

INVx2_ASAP7_75t_L g11523 ( 
.A(n_10851),
.Y(n_11523)
);

OR2x6_ASAP7_75t_L g11524 ( 
.A(n_10861),
.B(n_1502),
.Y(n_11524)
);

AOI21xp33_ASAP7_75t_SL g11525 ( 
.A1(n_10936),
.A2(n_775),
.B(n_776),
.Y(n_11525)
);

NAND2x1_ASAP7_75t_L g11526 ( 
.A(n_10851),
.B(n_775),
.Y(n_11526)
);

CKINVDCx11_ASAP7_75t_R g11527 ( 
.A(n_10861),
.Y(n_11527)
);

AOI21xp5_ASAP7_75t_L g11528 ( 
.A1(n_11160),
.A2(n_1503),
.B(n_1502),
.Y(n_11528)
);

INVx3_ASAP7_75t_L g11529 ( 
.A(n_10960),
.Y(n_11529)
);

INVx1_ASAP7_75t_L g11530 ( 
.A(n_11256),
.Y(n_11530)
);

OAI22xp5_ASAP7_75t_L g11531 ( 
.A1(n_11215),
.A2(n_778),
.B1(n_776),
.B2(n_777),
.Y(n_11531)
);

HB1xp67_ASAP7_75t_L g11532 ( 
.A(n_11260),
.Y(n_11532)
);

O2A1O1Ixp5_ASAP7_75t_L g11533 ( 
.A1(n_11214),
.A2(n_778),
.B(n_776),
.C(n_777),
.Y(n_11533)
);

INVx1_ASAP7_75t_L g11534 ( 
.A(n_11257),
.Y(n_11534)
);

AND2x2_ASAP7_75t_L g11535 ( 
.A(n_11244),
.B(n_777),
.Y(n_11535)
);

AOI21x1_ASAP7_75t_SL g11536 ( 
.A1(n_11237),
.A2(n_11365),
.B(n_11270),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_11209),
.B(n_1503),
.Y(n_11537)
);

INVx2_ASAP7_75t_L g11538 ( 
.A(n_11277),
.Y(n_11538)
);

AND2x2_ASAP7_75t_L g11539 ( 
.A(n_11220),
.B(n_778),
.Y(n_11539)
);

O2A1O1Ixp33_ASAP7_75t_L g11540 ( 
.A1(n_11397),
.A2(n_781),
.B(n_779),
.C(n_780),
.Y(n_11540)
);

OA21x2_ASAP7_75t_L g11541 ( 
.A1(n_11302),
.A2(n_779),
.B(n_780),
.Y(n_11541)
);

O2A1O1Ixp5_ASAP7_75t_L g11542 ( 
.A1(n_11267),
.A2(n_11358),
.B(n_11221),
.C(n_11271),
.Y(n_11542)
);

NAND2xp5_ASAP7_75t_L g11543 ( 
.A(n_11238),
.B(n_1504),
.Y(n_11543)
);

NAND2xp5_ASAP7_75t_L g11544 ( 
.A(n_11232),
.B(n_1504),
.Y(n_11544)
);

BUFx2_ASAP7_75t_L g11545 ( 
.A(n_11345),
.Y(n_11545)
);

BUFx2_ASAP7_75t_L g11546 ( 
.A(n_11225),
.Y(n_11546)
);

OAI22xp5_ASAP7_75t_L g11547 ( 
.A1(n_11300),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_11547)
);

OR2x2_ASAP7_75t_L g11548 ( 
.A(n_11240),
.B(n_782),
.Y(n_11548)
);

BUFx12f_ASAP7_75t_L g11549 ( 
.A(n_11527),
.Y(n_11549)
);

OR2x2_ASAP7_75t_L g11550 ( 
.A(n_11360),
.B(n_782),
.Y(n_11550)
);

OR2x6_ASAP7_75t_L g11551 ( 
.A(n_11522),
.B(n_1505),
.Y(n_11551)
);

OR2x2_ASAP7_75t_L g11552 ( 
.A(n_11295),
.B(n_782),
.Y(n_11552)
);

AO21x1_ASAP7_75t_L g11553 ( 
.A1(n_11391),
.A2(n_783),
.B(n_784),
.Y(n_11553)
);

INVx2_ASAP7_75t_L g11554 ( 
.A(n_11314),
.Y(n_11554)
);

O2A1O1Ixp33_ASAP7_75t_L g11555 ( 
.A1(n_11408),
.A2(n_785),
.B(n_783),
.C(n_784),
.Y(n_11555)
);

INVx1_ASAP7_75t_SL g11556 ( 
.A(n_11352),
.Y(n_11556)
);

AOI21xp5_ASAP7_75t_L g11557 ( 
.A1(n_11336),
.A2(n_783),
.B(n_784),
.Y(n_11557)
);

NAND2xp5_ASAP7_75t_L g11558 ( 
.A(n_11332),
.B(n_1508),
.Y(n_11558)
);

O2A1O1Ixp5_ASAP7_75t_L g11559 ( 
.A1(n_11526),
.A2(n_787),
.B(n_785),
.C(n_786),
.Y(n_11559)
);

O2A1O1Ixp33_ASAP7_75t_L g11560 ( 
.A1(n_11525),
.A2(n_787),
.B(n_785),
.C(n_786),
.Y(n_11560)
);

NAND2xp5_ASAP7_75t_L g11561 ( 
.A(n_11432),
.B(n_1508),
.Y(n_11561)
);

NAND2xp5_ASAP7_75t_L g11562 ( 
.A(n_11404),
.B(n_1509),
.Y(n_11562)
);

INVx2_ASAP7_75t_L g11563 ( 
.A(n_11243),
.Y(n_11563)
);

BUFx12f_ASAP7_75t_L g11564 ( 
.A(n_11521),
.Y(n_11564)
);

INVx4_ASAP7_75t_SL g11565 ( 
.A(n_11294),
.Y(n_11565)
);

AND2x2_ASAP7_75t_SL g11566 ( 
.A(n_11498),
.B(n_786),
.Y(n_11566)
);

O2A1O1Ixp33_ASAP7_75t_L g11567 ( 
.A1(n_11216),
.A2(n_789),
.B(n_787),
.C(n_788),
.Y(n_11567)
);

AND2x2_ASAP7_75t_L g11568 ( 
.A(n_11263),
.B(n_788),
.Y(n_11568)
);

AND2x2_ASAP7_75t_L g11569 ( 
.A(n_11274),
.B(n_788),
.Y(n_11569)
);

NOR2xp67_ASAP7_75t_L g11570 ( 
.A(n_11212),
.B(n_789),
.Y(n_11570)
);

INVx1_ASAP7_75t_L g11571 ( 
.A(n_11264),
.Y(n_11571)
);

AOI21x1_ASAP7_75t_SL g11572 ( 
.A1(n_11394),
.A2(n_789),
.B(n_790),
.Y(n_11572)
);

HB1xp67_ASAP7_75t_L g11573 ( 
.A(n_11286),
.Y(n_11573)
);

AND2x2_ASAP7_75t_L g11574 ( 
.A(n_11402),
.B(n_790),
.Y(n_11574)
);

AND2x2_ASAP7_75t_L g11575 ( 
.A(n_11411),
.B(n_11523),
.Y(n_11575)
);

OAI22xp5_ASAP7_75t_L g11576 ( 
.A1(n_11477),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.Y(n_11576)
);

NAND2xp5_ASAP7_75t_L g11577 ( 
.A(n_11304),
.B(n_1509),
.Y(n_11577)
);

INVx2_ASAP7_75t_L g11578 ( 
.A(n_11375),
.Y(n_11578)
);

O2A1O1Ixp5_ASAP7_75t_L g11579 ( 
.A1(n_11308),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_11579)
);

CKINVDCx20_ASAP7_75t_R g11580 ( 
.A(n_11235),
.Y(n_11580)
);

AND2x2_ASAP7_75t_L g11581 ( 
.A(n_11392),
.B(n_791),
.Y(n_11581)
);

OR2x2_ASAP7_75t_L g11582 ( 
.A(n_11268),
.B(n_11321),
.Y(n_11582)
);

OA21x2_ASAP7_75t_L g11583 ( 
.A1(n_11219),
.A2(n_792),
.B(n_793),
.Y(n_11583)
);

AOI21x1_ASAP7_75t_SL g11584 ( 
.A1(n_11288),
.A2(n_794),
.B(n_795),
.Y(n_11584)
);

OR2x2_ASAP7_75t_L g11585 ( 
.A(n_11223),
.B(n_794),
.Y(n_11585)
);

AOI21x1_ASAP7_75t_SL g11586 ( 
.A1(n_11387),
.A2(n_794),
.B(n_795),
.Y(n_11586)
);

INVx2_ASAP7_75t_SL g11587 ( 
.A(n_11291),
.Y(n_11587)
);

NAND2xp5_ASAP7_75t_L g11588 ( 
.A(n_11230),
.B(n_1511),
.Y(n_11588)
);

O2A1O1Ixp5_ASAP7_75t_L g11589 ( 
.A1(n_11502),
.A2(n_797),
.B(n_795),
.C(n_796),
.Y(n_11589)
);

A2O1A1Ixp33_ASAP7_75t_L g11590 ( 
.A1(n_11229),
.A2(n_798),
.B(n_796),
.C(n_797),
.Y(n_11590)
);

NAND2xp5_ASAP7_75t_L g11591 ( 
.A(n_11425),
.B(n_11429),
.Y(n_11591)
);

AND2x2_ASAP7_75t_L g11592 ( 
.A(n_11421),
.B(n_796),
.Y(n_11592)
);

AOI21xp5_ASAP7_75t_L g11593 ( 
.A1(n_11259),
.A2(n_797),
.B(n_798),
.Y(n_11593)
);

OAI22xp5_ASAP7_75t_L g11594 ( 
.A1(n_11276),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.Y(n_11594)
);

AOI21xp5_ASAP7_75t_L g11595 ( 
.A1(n_11278),
.A2(n_799),
.B(n_800),
.Y(n_11595)
);

AND2x2_ASAP7_75t_L g11596 ( 
.A(n_11218),
.B(n_800),
.Y(n_11596)
);

AND2x4_ASAP7_75t_L g11597 ( 
.A(n_11529),
.B(n_801),
.Y(n_11597)
);

AND2x2_ASAP7_75t_L g11598 ( 
.A(n_11403),
.B(n_801),
.Y(n_11598)
);

CKINVDCx14_ASAP7_75t_R g11599 ( 
.A(n_11439),
.Y(n_11599)
);

O2A1O1Ixp33_ASAP7_75t_L g11600 ( 
.A1(n_11284),
.A2(n_803),
.B(n_801),
.C(n_802),
.Y(n_11600)
);

AOI21xp5_ASAP7_75t_L g11601 ( 
.A1(n_11361),
.A2(n_11281),
.B(n_11504),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_11265),
.Y(n_11602)
);

NAND2xp5_ASAP7_75t_L g11603 ( 
.A(n_11247),
.B(n_1511),
.Y(n_11603)
);

AND2x2_ASAP7_75t_L g11604 ( 
.A(n_11452),
.B(n_11373),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_L g11605 ( 
.A(n_11252),
.B(n_1512),
.Y(n_11605)
);

AND2x2_ASAP7_75t_L g11606 ( 
.A(n_11427),
.B(n_803),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_11204),
.Y(n_11607)
);

AND2x2_ASAP7_75t_L g11608 ( 
.A(n_11431),
.B(n_803),
.Y(n_11608)
);

OAI22xp5_ASAP7_75t_L g11609 ( 
.A1(n_11283),
.A2(n_806),
.B1(n_804),
.B2(n_805),
.Y(n_11609)
);

OR2x2_ASAP7_75t_L g11610 ( 
.A(n_11206),
.B(n_804),
.Y(n_11610)
);

OR2x2_ASAP7_75t_L g11611 ( 
.A(n_11224),
.B(n_804),
.Y(n_11611)
);

AND2x2_ASAP7_75t_L g11612 ( 
.A(n_11383),
.B(n_805),
.Y(n_11612)
);

AND2x2_ASAP7_75t_L g11613 ( 
.A(n_11377),
.B(n_806),
.Y(n_11613)
);

NAND2xp5_ASAP7_75t_L g11614 ( 
.A(n_11440),
.B(n_1512),
.Y(n_11614)
);

INVx2_ASAP7_75t_L g11615 ( 
.A(n_11340),
.Y(n_11615)
);

NAND2xp5_ASAP7_75t_L g11616 ( 
.A(n_11450),
.B(n_1513),
.Y(n_11616)
);

INVx2_ASAP7_75t_L g11617 ( 
.A(n_11357),
.Y(n_11617)
);

AND2x2_ASAP7_75t_L g11618 ( 
.A(n_11475),
.B(n_806),
.Y(n_11618)
);

AOI21xp5_ASAP7_75t_L g11619 ( 
.A1(n_11389),
.A2(n_807),
.B(n_808),
.Y(n_11619)
);

AOI21xp5_ASAP7_75t_L g11620 ( 
.A1(n_11203),
.A2(n_11511),
.B(n_11528),
.Y(n_11620)
);

NAND2xp5_ASAP7_75t_L g11621 ( 
.A(n_11463),
.B(n_1513),
.Y(n_11621)
);

A2O1A1Ixp33_ASAP7_75t_L g11622 ( 
.A1(n_11325),
.A2(n_11348),
.B(n_11324),
.C(n_11359),
.Y(n_11622)
);

CKINVDCx20_ASAP7_75t_R g11623 ( 
.A(n_11310),
.Y(n_11623)
);

O2A1O1Ixp33_ASAP7_75t_L g11624 ( 
.A1(n_11433),
.A2(n_809),
.B(n_807),
.C(n_808),
.Y(n_11624)
);

AND2x4_ASAP7_75t_L g11625 ( 
.A(n_11455),
.B(n_807),
.Y(n_11625)
);

AOI221x1_ASAP7_75t_SL g11626 ( 
.A1(n_11250),
.A2(n_811),
.B1(n_809),
.B2(n_810),
.C(n_812),
.Y(n_11626)
);

NAND2xp5_ASAP7_75t_L g11627 ( 
.A(n_11242),
.B(n_1514),
.Y(n_11627)
);

BUFx3_ASAP7_75t_L g11628 ( 
.A(n_11294),
.Y(n_11628)
);

AND2x4_ASAP7_75t_L g11629 ( 
.A(n_11406),
.B(n_810),
.Y(n_11629)
);

AND2x2_ASAP7_75t_L g11630 ( 
.A(n_11273),
.B(n_810),
.Y(n_11630)
);

O2A1O1Ixp33_ASAP7_75t_L g11631 ( 
.A1(n_11462),
.A2(n_814),
.B(n_811),
.C(n_813),
.Y(n_11631)
);

AND2x4_ASAP7_75t_L g11632 ( 
.A(n_11349),
.B(n_811),
.Y(n_11632)
);

HB1xp67_ASAP7_75t_L g11633 ( 
.A(n_11258),
.Y(n_11633)
);

INVx1_ASAP7_75t_SL g11634 ( 
.A(n_11367),
.Y(n_11634)
);

BUFx6f_ASAP7_75t_SL g11635 ( 
.A(n_11524),
.Y(n_11635)
);

A2O1A1Ixp33_ASAP7_75t_L g11636 ( 
.A1(n_11418),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_11636)
);

CKINVDCx5p33_ASAP7_75t_R g11637 ( 
.A(n_11339),
.Y(n_11637)
);

INVx1_ASAP7_75t_L g11638 ( 
.A(n_11205),
.Y(n_11638)
);

AOI21xp5_ASAP7_75t_SL g11639 ( 
.A1(n_11480),
.A2(n_813),
.B(n_814),
.Y(n_11639)
);

OAI22xp5_ASAP7_75t_L g11640 ( 
.A1(n_11210),
.A2(n_817),
.B1(n_815),
.B2(n_816),
.Y(n_11640)
);

A2O1A1Ixp33_ASAP7_75t_L g11641 ( 
.A1(n_11388),
.A2(n_817),
.B(n_815),
.C(n_816),
.Y(n_11641)
);

A2O1A1Ixp33_ASAP7_75t_L g11642 ( 
.A1(n_11420),
.A2(n_818),
.B(n_816),
.C(n_817),
.Y(n_11642)
);

INVx1_ASAP7_75t_L g11643 ( 
.A(n_11249),
.Y(n_11643)
);

OA21x2_ASAP7_75t_L g11644 ( 
.A1(n_11346),
.A2(n_818),
.B(n_819),
.Y(n_11644)
);

NOR2x1_ASAP7_75t_SL g11645 ( 
.A(n_11446),
.B(n_818),
.Y(n_11645)
);

NAND2xp5_ASAP7_75t_L g11646 ( 
.A(n_11315),
.B(n_1514),
.Y(n_11646)
);

NAND2x1p5_ASAP7_75t_L g11647 ( 
.A(n_11514),
.B(n_819),
.Y(n_11647)
);

AND2x2_ASAP7_75t_L g11648 ( 
.A(n_11487),
.B(n_819),
.Y(n_11648)
);

OAI22xp5_ASAP7_75t_L g11649 ( 
.A1(n_11211),
.A2(n_822),
.B1(n_820),
.B2(n_821),
.Y(n_11649)
);

AOI21xp5_ASAP7_75t_L g11650 ( 
.A1(n_11241),
.A2(n_820),
.B(n_822),
.Y(n_11650)
);

OAI22xp5_ASAP7_75t_L g11651 ( 
.A1(n_11207),
.A2(n_824),
.B1(n_820),
.B2(n_823),
.Y(n_11651)
);

O2A1O1Ixp33_ASAP7_75t_L g11652 ( 
.A1(n_11486),
.A2(n_825),
.B(n_823),
.C(n_824),
.Y(n_11652)
);

AND2x2_ASAP7_75t_L g11653 ( 
.A(n_11493),
.B(n_823),
.Y(n_11653)
);

OR2x2_ASAP7_75t_L g11654 ( 
.A(n_11234),
.B(n_825),
.Y(n_11654)
);

HB1xp67_ASAP7_75t_L g11655 ( 
.A(n_11466),
.Y(n_11655)
);

AOI21xp5_ASAP7_75t_SL g11656 ( 
.A1(n_11434),
.A2(n_11398),
.B(n_11416),
.Y(n_11656)
);

AND2x2_ASAP7_75t_L g11657 ( 
.A(n_11293),
.B(n_826),
.Y(n_11657)
);

AND2x2_ASAP7_75t_L g11658 ( 
.A(n_11490),
.B(n_826),
.Y(n_11658)
);

HB1xp67_ASAP7_75t_L g11659 ( 
.A(n_11488),
.Y(n_11659)
);

OA21x2_ASAP7_75t_L g11660 ( 
.A1(n_11417),
.A2(n_826),
.B(n_827),
.Y(n_11660)
);

OA21x2_ASAP7_75t_L g11661 ( 
.A1(n_11280),
.A2(n_827),
.B(n_828),
.Y(n_11661)
);

AND2x2_ASAP7_75t_L g11662 ( 
.A(n_11478),
.B(n_11479),
.Y(n_11662)
);

OAI22xp5_ASAP7_75t_L g11663 ( 
.A1(n_11290),
.A2(n_829),
.B1(n_827),
.B2(n_828),
.Y(n_11663)
);

INVx2_ASAP7_75t_SL g11664 ( 
.A(n_11305),
.Y(n_11664)
);

NAND2xp5_ASAP7_75t_L g11665 ( 
.A(n_11517),
.B(n_1515),
.Y(n_11665)
);

AOI21xp5_ASAP7_75t_SL g11666 ( 
.A1(n_11516),
.A2(n_828),
.B(n_829),
.Y(n_11666)
);

OR2x2_ASAP7_75t_L g11667 ( 
.A(n_11261),
.B(n_829),
.Y(n_11667)
);

NAND2xp5_ASAP7_75t_L g11668 ( 
.A(n_11505),
.B(n_1516),
.Y(n_11668)
);

AND2x4_ASAP7_75t_L g11669 ( 
.A(n_11395),
.B(n_830),
.Y(n_11669)
);

NOR2xp67_ASAP7_75t_L g11670 ( 
.A(n_11366),
.B(n_11401),
.Y(n_11670)
);

INVx2_ASAP7_75t_L g11671 ( 
.A(n_11341),
.Y(n_11671)
);

INVx2_ASAP7_75t_L g11672 ( 
.A(n_11309),
.Y(n_11672)
);

INVxp33_ASAP7_75t_L g11673 ( 
.A(n_11413),
.Y(n_11673)
);

O2A1O1Ixp33_ASAP7_75t_L g11674 ( 
.A1(n_11430),
.A2(n_832),
.B(n_830),
.C(n_831),
.Y(n_11674)
);

NAND2xp5_ASAP7_75t_L g11675 ( 
.A(n_11356),
.B(n_1516),
.Y(n_11675)
);

A2O1A1Ixp33_ASAP7_75t_SL g11676 ( 
.A1(n_11292),
.A2(n_833),
.B(n_830),
.C(n_832),
.Y(n_11676)
);

AND2x2_ASAP7_75t_L g11677 ( 
.A(n_11282),
.B(n_832),
.Y(n_11677)
);

O2A1O1Ixp5_ASAP7_75t_L g11678 ( 
.A1(n_11436),
.A2(n_835),
.B(n_833),
.C(n_834),
.Y(n_11678)
);

AOI21xp5_ASAP7_75t_L g11679 ( 
.A1(n_11253),
.A2(n_833),
.B(n_834),
.Y(n_11679)
);

NOR2xp67_ASAP7_75t_L g11680 ( 
.A(n_11217),
.B(n_834),
.Y(n_11680)
);

HB1xp67_ASAP7_75t_L g11681 ( 
.A(n_11269),
.Y(n_11681)
);

INVx1_ASAP7_75t_SL g11682 ( 
.A(n_11227),
.Y(n_11682)
);

AND2x4_ASAP7_75t_L g11683 ( 
.A(n_11453),
.B(n_835),
.Y(n_11683)
);

INVx1_ASAP7_75t_L g11684 ( 
.A(n_11255),
.Y(n_11684)
);

INVx1_ASAP7_75t_L g11685 ( 
.A(n_11518),
.Y(n_11685)
);

INVxp67_ASAP7_75t_L g11686 ( 
.A(n_11445),
.Y(n_11686)
);

NAND2xp5_ASAP7_75t_L g11687 ( 
.A(n_11269),
.B(n_1517),
.Y(n_11687)
);

O2A1O1Ixp33_ASAP7_75t_L g11688 ( 
.A1(n_11464),
.A2(n_837),
.B(n_835),
.C(n_836),
.Y(n_11688)
);

CKINVDCx5p33_ASAP7_75t_R g11689 ( 
.A(n_11317),
.Y(n_11689)
);

OAI22xp5_ASAP7_75t_L g11690 ( 
.A1(n_11298),
.A2(n_838),
.B1(n_836),
.B2(n_837),
.Y(n_11690)
);

AND2x2_ASAP7_75t_L g11691 ( 
.A(n_11313),
.B(n_838),
.Y(n_11691)
);

INVx2_ASAP7_75t_L g11692 ( 
.A(n_11246),
.Y(n_11692)
);

A2O1A1Ixp33_ASAP7_75t_L g11693 ( 
.A1(n_11279),
.A2(n_841),
.B(n_839),
.C(n_840),
.Y(n_11693)
);

OA21x2_ASAP7_75t_L g11694 ( 
.A1(n_11208),
.A2(n_839),
.B(n_840),
.Y(n_11694)
);

AOI21xp5_ASAP7_75t_L g11695 ( 
.A1(n_11506),
.A2(n_839),
.B(n_840),
.Y(n_11695)
);

OR2x2_ASAP7_75t_SL g11696 ( 
.A(n_11472),
.B(n_841),
.Y(n_11696)
);

OAI22xp5_ASAP7_75t_L g11697 ( 
.A1(n_11444),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_11697)
);

OA21x2_ASAP7_75t_L g11698 ( 
.A1(n_11299),
.A2(n_842),
.B(n_843),
.Y(n_11698)
);

INVx2_ASAP7_75t_L g11699 ( 
.A(n_11254),
.Y(n_11699)
);

NAND2xp5_ASAP7_75t_L g11700 ( 
.A(n_11330),
.B(n_1517),
.Y(n_11700)
);

NAND2xp5_ASAP7_75t_L g11701 ( 
.A(n_11363),
.B(n_1518),
.Y(n_11701)
);

AND2x2_ASAP7_75t_L g11702 ( 
.A(n_11509),
.B(n_843),
.Y(n_11702)
);

OR2x2_ASAP7_75t_L g11703 ( 
.A(n_11307),
.B(n_844),
.Y(n_11703)
);

A2O1A1Ixp33_ASAP7_75t_L g11704 ( 
.A1(n_11233),
.A2(n_846),
.B(n_844),
.C(n_845),
.Y(n_11704)
);

BUFx4f_ASAP7_75t_L g11705 ( 
.A(n_11459),
.Y(n_11705)
);

INVx2_ASAP7_75t_SL g11706 ( 
.A(n_11328),
.Y(n_11706)
);

HB1xp67_ASAP7_75t_L g11707 ( 
.A(n_11428),
.Y(n_11707)
);

OAI22xp5_ASAP7_75t_L g11708 ( 
.A1(n_11423),
.A2(n_846),
.B1(n_844),
.B2(n_845),
.Y(n_11708)
);

INVx2_ASAP7_75t_L g11709 ( 
.A(n_11272),
.Y(n_11709)
);

AND2x2_ASAP7_75t_L g11710 ( 
.A(n_11285),
.B(n_845),
.Y(n_11710)
);

AND2x2_ASAP7_75t_L g11711 ( 
.A(n_11275),
.B(n_847),
.Y(n_11711)
);

NOR2xp67_ASAP7_75t_L g11712 ( 
.A(n_11470),
.B(n_847),
.Y(n_11712)
);

O2A1O1Ixp33_ASAP7_75t_L g11713 ( 
.A1(n_11508),
.A2(n_849),
.B(n_847),
.C(n_848),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_11228),
.B(n_848),
.Y(n_11714)
);

AND2x4_ASAP7_75t_L g11715 ( 
.A(n_11503),
.B(n_849),
.Y(n_11715)
);

OAI22xp5_ASAP7_75t_SL g11716 ( 
.A1(n_11335),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_11301),
.B(n_1519),
.Y(n_11717)
);

A2O1A1Ixp33_ASAP7_75t_L g11718 ( 
.A1(n_11262),
.A2(n_852),
.B(n_850),
.C(n_851),
.Y(n_11718)
);

HB1xp67_ASAP7_75t_L g11719 ( 
.A(n_11471),
.Y(n_11719)
);

A2O1A1Ixp33_ASAP7_75t_L g11720 ( 
.A1(n_11266),
.A2(n_853),
.B(n_851),
.C(n_852),
.Y(n_11720)
);

NAND2xp5_ASAP7_75t_L g11721 ( 
.A(n_11316),
.B(n_1519),
.Y(n_11721)
);

AND2x2_ASAP7_75t_L g11722 ( 
.A(n_11231),
.B(n_853),
.Y(n_11722)
);

HB1xp67_ASAP7_75t_L g11723 ( 
.A(n_11327),
.Y(n_11723)
);

OA21x2_ASAP7_75t_L g11724 ( 
.A1(n_11248),
.A2(n_854),
.B(n_855),
.Y(n_11724)
);

INVx2_ASAP7_75t_L g11725 ( 
.A(n_11320),
.Y(n_11725)
);

OAI22xp5_ASAP7_75t_L g11726 ( 
.A1(n_11501),
.A2(n_856),
.B1(n_854),
.B2(n_855),
.Y(n_11726)
);

AOI21xp5_ASAP7_75t_L g11727 ( 
.A1(n_11296),
.A2(n_854),
.B(n_855),
.Y(n_11727)
);

AOI21xp5_ASAP7_75t_L g11728 ( 
.A1(n_11226),
.A2(n_856),
.B(n_857),
.Y(n_11728)
);

INVx1_ASAP7_75t_L g11729 ( 
.A(n_11351),
.Y(n_11729)
);

AOI21xp5_ASAP7_75t_L g11730 ( 
.A1(n_11236),
.A2(n_856),
.B(n_857),
.Y(n_11730)
);

NAND2xp5_ASAP7_75t_L g11731 ( 
.A(n_11297),
.B(n_1520),
.Y(n_11731)
);

A2O1A1Ixp33_ASAP7_75t_L g11732 ( 
.A1(n_11484),
.A2(n_859),
.B(n_857),
.C(n_858),
.Y(n_11732)
);

AND2x4_ASAP7_75t_L g11733 ( 
.A(n_11520),
.B(n_11331),
.Y(n_11733)
);

CKINVDCx5p33_ASAP7_75t_R g11734 ( 
.A(n_11414),
.Y(n_11734)
);

INVx3_ASAP7_75t_L g11735 ( 
.A(n_11331),
.Y(n_11735)
);

OAI22xp5_ASAP7_75t_L g11736 ( 
.A1(n_11385),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_11736)
);

AND2x2_ASAP7_75t_L g11737 ( 
.A(n_11386),
.B(n_858),
.Y(n_11737)
);

OAI22xp5_ASAP7_75t_L g11738 ( 
.A1(n_11342),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.Y(n_11738)
);

AND2x4_ASAP7_75t_L g11739 ( 
.A(n_11386),
.B(n_860),
.Y(n_11739)
);

O2A1O1Ixp33_ASAP7_75t_L g11740 ( 
.A1(n_11326),
.A2(n_863),
.B(n_861),
.C(n_862),
.Y(n_11740)
);

AND2x4_ASAP7_75t_L g11741 ( 
.A(n_11405),
.B(n_861),
.Y(n_11741)
);

AND2x2_ASAP7_75t_L g11742 ( 
.A(n_11405),
.B(n_862),
.Y(n_11742)
);

HB1xp67_ASAP7_75t_L g11743 ( 
.A(n_11312),
.Y(n_11743)
);

OR2x2_ASAP7_75t_L g11744 ( 
.A(n_11350),
.B(n_862),
.Y(n_11744)
);

AND2x4_ASAP7_75t_L g11745 ( 
.A(n_11419),
.B(n_863),
.Y(n_11745)
);

AND2x2_ASAP7_75t_L g11746 ( 
.A(n_11419),
.B(n_863),
.Y(n_11746)
);

INVx2_ASAP7_75t_L g11747 ( 
.A(n_11306),
.Y(n_11747)
);

O2A1O1Ixp33_ASAP7_75t_L g11748 ( 
.A1(n_11368),
.A2(n_866),
.B(n_864),
.C(n_865),
.Y(n_11748)
);

INVx1_ASAP7_75t_L g11749 ( 
.A(n_11519),
.Y(n_11749)
);

OAI22xp5_ASAP7_75t_L g11750 ( 
.A1(n_11513),
.A2(n_866),
.B1(n_864),
.B2(n_865),
.Y(n_11750)
);

O2A1O1Ixp5_ASAP7_75t_L g11751 ( 
.A1(n_11376),
.A2(n_869),
.B(n_867),
.C(n_868),
.Y(n_11751)
);

AND2x2_ASAP7_75t_L g11752 ( 
.A(n_11369),
.B(n_867),
.Y(n_11752)
);

AOI21xp33_ASAP7_75t_L g11753 ( 
.A1(n_11289),
.A2(n_867),
.B(n_868),
.Y(n_11753)
);

INVx1_ASAP7_75t_L g11754 ( 
.A(n_11343),
.Y(n_11754)
);

AOI21xp5_ASAP7_75t_L g11755 ( 
.A1(n_11239),
.A2(n_11222),
.B(n_11473),
.Y(n_11755)
);

OAI22xp5_ASAP7_75t_L g11756 ( 
.A1(n_11322),
.A2(n_870),
.B1(n_868),
.B2(n_869),
.Y(n_11756)
);

NAND2xp5_ASAP7_75t_L g11757 ( 
.A(n_11424),
.B(n_1520),
.Y(n_11757)
);

O2A1O1Ixp33_ASAP7_75t_L g11758 ( 
.A1(n_11456),
.A2(n_870),
.B(n_1522),
.C(n_1521),
.Y(n_11758)
);

OAI22xp5_ASAP7_75t_L g11759 ( 
.A1(n_11355),
.A2(n_1523),
.B1(n_1521),
.B2(n_1522),
.Y(n_11759)
);

O2A1O1Ixp5_ASAP7_75t_L g11760 ( 
.A1(n_11347),
.A2(n_1525),
.B(n_1523),
.C(n_1524),
.Y(n_11760)
);

A2O1A1Ixp33_ASAP7_75t_L g11761 ( 
.A1(n_11495),
.A2(n_1526),
.B(n_1524),
.C(n_1525),
.Y(n_11761)
);

AND2x2_ASAP7_75t_L g11762 ( 
.A(n_11362),
.B(n_1526),
.Y(n_11762)
);

A2O1A1Ixp33_ASAP7_75t_L g11763 ( 
.A1(n_11344),
.A2(n_1529),
.B(n_1527),
.C(n_1528),
.Y(n_11763)
);

AND2x2_ASAP7_75t_L g11764 ( 
.A(n_11303),
.B(n_1527),
.Y(n_11764)
);

OAI22xp5_ASAP7_75t_L g11765 ( 
.A1(n_11337),
.A2(n_1531),
.B1(n_1528),
.B2(n_1530),
.Y(n_11765)
);

O2A1O1Ixp33_ASAP7_75t_L g11766 ( 
.A1(n_11323),
.A2(n_1533),
.B(n_1531),
.C(n_1532),
.Y(n_11766)
);

O2A1O1Ixp33_ASAP7_75t_L g11767 ( 
.A1(n_11492),
.A2(n_1534),
.B(n_1532),
.C(n_1533),
.Y(n_11767)
);

NAND2xp5_ASAP7_75t_L g11768 ( 
.A(n_11380),
.B(n_11458),
.Y(n_11768)
);

OAI22xp5_ASAP7_75t_SL g11769 ( 
.A1(n_11512),
.A2(n_1537),
.B1(n_1535),
.B2(n_1536),
.Y(n_11769)
);

INVx2_ASAP7_75t_L g11770 ( 
.A(n_11333),
.Y(n_11770)
);

NAND2xp5_ASAP7_75t_L g11771 ( 
.A(n_11370),
.B(n_11371),
.Y(n_11771)
);

AOI21xp5_ASAP7_75t_SL g11772 ( 
.A1(n_11438),
.A2(n_1535),
.B(n_1536),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_11460),
.Y(n_11773)
);

HB1xp67_ASAP7_75t_L g11774 ( 
.A(n_11467),
.Y(n_11774)
);

O2A1O1Ixp33_ASAP7_75t_L g11775 ( 
.A1(n_11379),
.A2(n_1539),
.B(n_1537),
.C(n_1538),
.Y(n_11775)
);

BUFx6f_ASAP7_75t_L g11776 ( 
.A(n_11412),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_11311),
.Y(n_11777)
);

OAI22xp5_ASAP7_75t_L g11778 ( 
.A1(n_11338),
.A2(n_1542),
.B1(n_1540),
.B2(n_1541),
.Y(n_11778)
);

INVx1_ASAP7_75t_SL g11779 ( 
.A(n_11476),
.Y(n_11779)
);

INVx2_ASAP7_75t_L g11780 ( 
.A(n_11318),
.Y(n_11780)
);

AND2x2_ASAP7_75t_L g11781 ( 
.A(n_11474),
.B(n_1541),
.Y(n_11781)
);

OAI22xp5_ASAP7_75t_L g11782 ( 
.A1(n_11354),
.A2(n_1545),
.B1(n_1543),
.B2(n_1544),
.Y(n_11782)
);

O2A1O1Ixp5_ASAP7_75t_L g11783 ( 
.A1(n_11443),
.A2(n_1545),
.B(n_1543),
.C(n_1544),
.Y(n_11783)
);

AOI21xp5_ASAP7_75t_L g11784 ( 
.A1(n_11213),
.A2(n_1546),
.B(n_1547),
.Y(n_11784)
);

CKINVDCx14_ASAP7_75t_R g11785 ( 
.A(n_11329),
.Y(n_11785)
);

AOI21x1_ASAP7_75t_SL g11786 ( 
.A1(n_11381),
.A2(n_1546),
.B(n_1547),
.Y(n_11786)
);

BUFx3_ASAP7_75t_L g11787 ( 
.A(n_11489),
.Y(n_11787)
);

OR2x2_ASAP7_75t_L g11788 ( 
.A(n_11287),
.B(n_1548),
.Y(n_11788)
);

O2A1O1Ixp33_ASAP7_75t_L g11789 ( 
.A1(n_11448),
.A2(n_1550),
.B(n_1548),
.C(n_1549),
.Y(n_11789)
);

AOI21xp5_ASAP7_75t_L g11790 ( 
.A1(n_11481),
.A2(n_1550),
.B(n_1551),
.Y(n_11790)
);

NAND2xp5_ASAP7_75t_L g11791 ( 
.A(n_11371),
.B(n_1552),
.Y(n_11791)
);

OA21x2_ASAP7_75t_L g11792 ( 
.A1(n_11251),
.A2(n_1553),
.B(n_1555),
.Y(n_11792)
);

NAND2xp5_ASAP7_75t_L g11793 ( 
.A(n_11287),
.B(n_1555),
.Y(n_11793)
);

OR2x2_ASAP7_75t_L g11794 ( 
.A(n_11245),
.B(n_1556),
.Y(n_11794)
);

OAI22xp5_ASAP7_75t_L g11795 ( 
.A1(n_11393),
.A2(n_11399),
.B1(n_11447),
.B2(n_11426),
.Y(n_11795)
);

AND2x2_ASAP7_75t_L g11796 ( 
.A(n_11364),
.B(n_1556),
.Y(n_11796)
);

AOI21x1_ASAP7_75t_SL g11797 ( 
.A1(n_11482),
.A2(n_1557),
.B(n_1558),
.Y(n_11797)
);

HB1xp67_ASAP7_75t_L g11798 ( 
.A(n_11319),
.Y(n_11798)
);

BUFx3_ASAP7_75t_L g11799 ( 
.A(n_11500),
.Y(n_11799)
);

OAI22xp5_ASAP7_75t_L g11800 ( 
.A1(n_11437),
.A2(n_1560),
.B1(n_1558),
.B2(n_1559),
.Y(n_11800)
);

A2O1A1Ixp33_ASAP7_75t_L g11801 ( 
.A1(n_11499),
.A2(n_1562),
.B(n_1560),
.C(n_1561),
.Y(n_11801)
);

OA21x2_ASAP7_75t_L g11802 ( 
.A1(n_11334),
.A2(n_1562),
.B(n_1563),
.Y(n_11802)
);

O2A1O1Ixp33_ASAP7_75t_L g11803 ( 
.A1(n_11415),
.A2(n_1565),
.B(n_1563),
.C(n_1564),
.Y(n_11803)
);

INVx2_ASAP7_75t_L g11804 ( 
.A(n_11372),
.Y(n_11804)
);

INVx2_ASAP7_75t_L g11805 ( 
.A(n_11374),
.Y(n_11805)
);

BUFx4f_ASAP7_75t_SL g11806 ( 
.A(n_11497),
.Y(n_11806)
);

OAI22xp5_ASAP7_75t_L g11807 ( 
.A1(n_11442),
.A2(n_1567),
.B1(n_1565),
.B2(n_1566),
.Y(n_11807)
);

AND2x2_ASAP7_75t_L g11808 ( 
.A(n_11483),
.B(n_1567),
.Y(n_11808)
);

AND2x2_ASAP7_75t_L g11809 ( 
.A(n_11491),
.B(n_1568),
.Y(n_11809)
);

HB1xp67_ASAP7_75t_L g11810 ( 
.A(n_11382),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_11378),
.Y(n_11811)
);

NAND2xp5_ASAP7_75t_SL g11812 ( 
.A(n_11507),
.B(n_1568),
.Y(n_11812)
);

INVx1_ASAP7_75t_L g11813 ( 
.A(n_11384),
.Y(n_11813)
);

O2A1O1Ixp5_ASAP7_75t_L g11814 ( 
.A1(n_11485),
.A2(n_1571),
.B(n_1569),
.C(n_1570),
.Y(n_11814)
);

O2A1O1Ixp33_ASAP7_75t_L g11815 ( 
.A1(n_11469),
.A2(n_1573),
.B(n_1571),
.C(n_1572),
.Y(n_11815)
);

CKINVDCx5p33_ASAP7_75t_R g11816 ( 
.A(n_11382),
.Y(n_11816)
);

INVx1_ASAP7_75t_L g11817 ( 
.A(n_11390),
.Y(n_11817)
);

INVx2_ASAP7_75t_L g11818 ( 
.A(n_11400),
.Y(n_11818)
);

OA21x2_ASAP7_75t_L g11819 ( 
.A1(n_11353),
.A2(n_1572),
.B(n_1574),
.Y(n_11819)
);

INVx2_ASAP7_75t_L g11820 ( 
.A(n_11409),
.Y(n_11820)
);

AND2x4_ASAP7_75t_L g11821 ( 
.A(n_11496),
.B(n_1574),
.Y(n_11821)
);

OA21x2_ASAP7_75t_L g11822 ( 
.A1(n_11407),
.A2(n_1575),
.B(n_1576),
.Y(n_11822)
);

AND2x2_ASAP7_75t_L g11823 ( 
.A(n_11396),
.B(n_1577),
.Y(n_11823)
);

OR2x2_ASAP7_75t_L g11824 ( 
.A(n_11396),
.B(n_1577),
.Y(n_11824)
);

O2A1O1Ixp33_ASAP7_75t_L g11825 ( 
.A1(n_11494),
.A2(n_1580),
.B(n_1578),
.C(n_1579),
.Y(n_11825)
);

OA21x2_ASAP7_75t_L g11826 ( 
.A1(n_11410),
.A2(n_1578),
.B(n_1580),
.Y(n_11826)
);

AOI21xp5_ASAP7_75t_SL g11827 ( 
.A1(n_11510),
.A2(n_1581),
.B(n_1582),
.Y(n_11827)
);

AOI21xp5_ASAP7_75t_SL g11828 ( 
.A1(n_11494),
.A2(n_1582),
.B(n_1583),
.Y(n_11828)
);

NAND2xp5_ASAP7_75t_L g11829 ( 
.A(n_11422),
.B(n_1584),
.Y(n_11829)
);

O2A1O1Ixp33_ASAP7_75t_L g11830 ( 
.A1(n_11515),
.A2(n_1587),
.B(n_1584),
.C(n_1586),
.Y(n_11830)
);

OR2x2_ASAP7_75t_L g11831 ( 
.A(n_11435),
.B(n_1586),
.Y(n_11831)
);

INVx1_ASAP7_75t_SL g11832 ( 
.A(n_11441),
.Y(n_11832)
);

AOI21xp5_ASAP7_75t_L g11833 ( 
.A1(n_11449),
.A2(n_1587),
.B(n_1588),
.Y(n_11833)
);

O2A1O1Ixp5_ASAP7_75t_L g11834 ( 
.A1(n_11451),
.A2(n_1590),
.B(n_1588),
.C(n_1589),
.Y(n_11834)
);

AND2x2_ASAP7_75t_L g11835 ( 
.A(n_11454),
.B(n_1589),
.Y(n_11835)
);

OAI22xp5_ASAP7_75t_L g11836 ( 
.A1(n_11457),
.A2(n_1592),
.B1(n_1590),
.B2(n_1591),
.Y(n_11836)
);

AND2x2_ASAP7_75t_L g11837 ( 
.A(n_11461),
.B(n_1591),
.Y(n_11837)
);

NOR2xp67_ASAP7_75t_L g11838 ( 
.A(n_11465),
.B(n_1592),
.Y(n_11838)
);

INVx1_ASAP7_75t_L g11839 ( 
.A(n_11468),
.Y(n_11839)
);

O2A1O1Ixp33_ASAP7_75t_L g11840 ( 
.A1(n_11397),
.A2(n_1595),
.B(n_1593),
.C(n_1594),
.Y(n_11840)
);

NAND2xp5_ASAP7_75t_L g11841 ( 
.A(n_11209),
.B(n_1593),
.Y(n_11841)
);

HB1xp67_ASAP7_75t_L g11842 ( 
.A(n_11260),
.Y(n_11842)
);

AOI21xp5_ASAP7_75t_SL g11843 ( 
.A1(n_11304),
.A2(n_1595),
.B(n_1596),
.Y(n_11843)
);

AND2x2_ASAP7_75t_L g11844 ( 
.A(n_11244),
.B(n_1596),
.Y(n_11844)
);

AND2x4_ASAP7_75t_L g11845 ( 
.A(n_11529),
.B(n_1597),
.Y(n_11845)
);

OA22x2_ASAP7_75t_L g11846 ( 
.A1(n_11271),
.A2(n_1599),
.B1(n_1597),
.B2(n_1598),
.Y(n_11846)
);

BUFx2_ASAP7_75t_SL g11847 ( 
.A(n_11366),
.Y(n_11847)
);

NAND2xp5_ASAP7_75t_L g11848 ( 
.A(n_11209),
.B(n_1598),
.Y(n_11848)
);

INVx2_ASAP7_75t_L g11849 ( 
.A(n_11277),
.Y(n_11849)
);

O2A1O1Ixp5_ASAP7_75t_L g11850 ( 
.A1(n_11214),
.A2(n_1602),
.B(n_1600),
.C(n_1601),
.Y(n_11850)
);

AOI21xp33_ASAP7_75t_L g11851 ( 
.A1(n_11215),
.A2(n_1601),
.B(n_1602),
.Y(n_11851)
);

AND2x2_ASAP7_75t_L g11852 ( 
.A(n_11244),
.B(n_1603),
.Y(n_11852)
);

AND2x2_ASAP7_75t_L g11853 ( 
.A(n_11244),
.B(n_1603),
.Y(n_11853)
);

NAND2xp5_ASAP7_75t_L g11854 ( 
.A(n_11209),
.B(n_1604),
.Y(n_11854)
);

OR2x2_ASAP7_75t_L g11855 ( 
.A(n_11240),
.B(n_1604),
.Y(n_11855)
);

OAI22xp5_ASAP7_75t_L g11856 ( 
.A1(n_11215),
.A2(n_1608),
.B1(n_1606),
.B2(n_1607),
.Y(n_11856)
);

CKINVDCx6p67_ASAP7_75t_R g11857 ( 
.A(n_11527),
.Y(n_11857)
);

AOI21x1_ASAP7_75t_SL g11858 ( 
.A1(n_11237),
.A2(n_1606),
.B(n_1607),
.Y(n_11858)
);

AND2x2_ASAP7_75t_L g11859 ( 
.A(n_11244),
.B(n_1608),
.Y(n_11859)
);

AOI22xp5_ASAP7_75t_L g11860 ( 
.A1(n_11566),
.A2(n_1611),
.B1(n_1609),
.B2(n_1610),
.Y(n_11860)
);

INVxp67_ASAP7_75t_L g11861 ( 
.A(n_11545),
.Y(n_11861)
);

INVx3_ASAP7_75t_L g11862 ( 
.A(n_11549),
.Y(n_11862)
);

INVx1_ASAP7_75t_L g11863 ( 
.A(n_11659),
.Y(n_11863)
);

HB1xp67_ASAP7_75t_L g11864 ( 
.A(n_11532),
.Y(n_11864)
);

NAND2xp5_ASAP7_75t_L g11865 ( 
.A(n_11727),
.B(n_1609),
.Y(n_11865)
);

OR2x2_ASAP7_75t_L g11866 ( 
.A(n_11582),
.B(n_1610),
.Y(n_11866)
);

BUFx2_ASAP7_75t_L g11867 ( 
.A(n_11599),
.Y(n_11867)
);

OAI21x1_ASAP7_75t_SL g11868 ( 
.A1(n_11620),
.A2(n_1611),
.B(n_1612),
.Y(n_11868)
);

BUFx2_ASAP7_75t_L g11869 ( 
.A(n_11546),
.Y(n_11869)
);

AND2x2_ASAP7_75t_L g11870 ( 
.A(n_11575),
.B(n_1613),
.Y(n_11870)
);

INVx1_ASAP7_75t_L g11871 ( 
.A(n_11530),
.Y(n_11871)
);

HB1xp67_ASAP7_75t_L g11872 ( 
.A(n_11842),
.Y(n_11872)
);

INVx1_ASAP7_75t_L g11873 ( 
.A(n_11534),
.Y(n_11873)
);

AND2x2_ASAP7_75t_L g11874 ( 
.A(n_11604),
.B(n_1613),
.Y(n_11874)
);

INVx1_ASAP7_75t_L g11875 ( 
.A(n_11571),
.Y(n_11875)
);

HB1xp67_ASAP7_75t_L g11876 ( 
.A(n_11723),
.Y(n_11876)
);

INVx1_ASAP7_75t_L g11877 ( 
.A(n_11602),
.Y(n_11877)
);

OR2x2_ASAP7_75t_L g11878 ( 
.A(n_11771),
.B(n_1614),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11607),
.Y(n_11879)
);

INVx2_ASAP7_75t_L g11880 ( 
.A(n_11664),
.Y(n_11880)
);

INVx2_ASAP7_75t_L g11881 ( 
.A(n_11662),
.Y(n_11881)
);

HB1xp67_ASAP7_75t_L g11882 ( 
.A(n_11573),
.Y(n_11882)
);

INVx1_ASAP7_75t_L g11883 ( 
.A(n_11638),
.Y(n_11883)
);

INVx2_ASAP7_75t_L g11884 ( 
.A(n_11787),
.Y(n_11884)
);

AO21x2_ASAP7_75t_L g11885 ( 
.A1(n_11681),
.A2(n_1615),
.B(n_1616),
.Y(n_11885)
);

INVx2_ASAP7_75t_L g11886 ( 
.A(n_11587),
.Y(n_11886)
);

HB1xp67_ASAP7_75t_L g11887 ( 
.A(n_11644),
.Y(n_11887)
);

BUFx3_ASAP7_75t_L g11888 ( 
.A(n_11564),
.Y(n_11888)
);

INVx2_ASAP7_75t_L g11889 ( 
.A(n_11706),
.Y(n_11889)
);

HB1xp67_ASAP7_75t_L g11890 ( 
.A(n_11644),
.Y(n_11890)
);

INVxp67_ASAP7_75t_L g11891 ( 
.A(n_11847),
.Y(n_11891)
);

INVx2_ASAP7_75t_L g11892 ( 
.A(n_11735),
.Y(n_11892)
);

BUFx3_ASAP7_75t_L g11893 ( 
.A(n_11857),
.Y(n_11893)
);

CKINVDCx5p33_ASAP7_75t_R g11894 ( 
.A(n_11580),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_11643),
.Y(n_11895)
);

NAND2xp5_ASAP7_75t_L g11896 ( 
.A(n_11679),
.B(n_1615),
.Y(n_11896)
);

INVx2_ASAP7_75t_L g11897 ( 
.A(n_11682),
.Y(n_11897)
);

INVx1_ASAP7_75t_L g11898 ( 
.A(n_11684),
.Y(n_11898)
);

AND2x2_ASAP7_75t_L g11899 ( 
.A(n_11779),
.B(n_1616),
.Y(n_11899)
);

OA21x2_ASAP7_75t_L g11900 ( 
.A1(n_11542),
.A2(n_1617),
.B(n_1618),
.Y(n_11900)
);

BUFx6f_ASAP7_75t_L g11901 ( 
.A(n_11715),
.Y(n_11901)
);

INVx2_ASAP7_75t_L g11902 ( 
.A(n_11628),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_11685),
.Y(n_11903)
);

NAND2xp33_ASAP7_75t_R g11904 ( 
.A(n_11661),
.B(n_1617),
.Y(n_11904)
);

INVx2_ASAP7_75t_L g11905 ( 
.A(n_11565),
.Y(n_11905)
);

INVx1_ASAP7_75t_L g11906 ( 
.A(n_11729),
.Y(n_11906)
);

INVx2_ASAP7_75t_L g11907 ( 
.A(n_11565),
.Y(n_11907)
);

INVx1_ASAP7_75t_L g11908 ( 
.A(n_11725),
.Y(n_11908)
);

INVx1_ASAP7_75t_L g11909 ( 
.A(n_11660),
.Y(n_11909)
);

AND2x2_ASAP7_75t_L g11910 ( 
.A(n_11634),
.B(n_11615),
.Y(n_11910)
);

INVx1_ASAP7_75t_L g11911 ( 
.A(n_11660),
.Y(n_11911)
);

BUFx3_ASAP7_75t_L g11912 ( 
.A(n_11623),
.Y(n_11912)
);

INVx1_ASAP7_75t_L g11913 ( 
.A(n_11661),
.Y(n_11913)
);

INVx1_ASAP7_75t_L g11914 ( 
.A(n_11810),
.Y(n_11914)
);

INVx2_ASAP7_75t_SL g11915 ( 
.A(n_11776),
.Y(n_11915)
);

INVx3_ASAP7_75t_L g11916 ( 
.A(n_11776),
.Y(n_11916)
);

INVx2_ASAP7_75t_L g11917 ( 
.A(n_11733),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_11699),
.Y(n_11918)
);

AND2x2_ASAP7_75t_L g11919 ( 
.A(n_11617),
.B(n_1619),
.Y(n_11919)
);

BUFx3_ASAP7_75t_L g11920 ( 
.A(n_11734),
.Y(n_11920)
);

INVx3_ASAP7_75t_L g11921 ( 
.A(n_11799),
.Y(n_11921)
);

BUFx2_ASAP7_75t_SL g11922 ( 
.A(n_11635),
.Y(n_11922)
);

INVx3_ASAP7_75t_L g11923 ( 
.A(n_11625),
.Y(n_11923)
);

INVx1_ASAP7_75t_L g11924 ( 
.A(n_11709),
.Y(n_11924)
);

OA21x2_ASAP7_75t_L g11925 ( 
.A1(n_11538),
.A2(n_1619),
.B(n_1620),
.Y(n_11925)
);

BUFx6f_ASAP7_75t_L g11926 ( 
.A(n_11683),
.Y(n_11926)
);

INVx2_ASAP7_75t_L g11927 ( 
.A(n_11563),
.Y(n_11927)
);

INVx1_ASAP7_75t_L g11928 ( 
.A(n_11774),
.Y(n_11928)
);

INVx3_ASAP7_75t_L g11929 ( 
.A(n_11669),
.Y(n_11929)
);

INVx5_ASAP7_75t_L g11930 ( 
.A(n_11677),
.Y(n_11930)
);

INVx1_ASAP7_75t_L g11931 ( 
.A(n_11541),
.Y(n_11931)
);

INVx2_ASAP7_75t_L g11932 ( 
.A(n_11578),
.Y(n_11932)
);

INVx2_ASAP7_75t_L g11933 ( 
.A(n_11671),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11541),
.Y(n_11934)
);

INVx2_ASAP7_75t_L g11935 ( 
.A(n_11672),
.Y(n_11935)
);

BUFx3_ASAP7_75t_L g11936 ( 
.A(n_11597),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11703),
.Y(n_11937)
);

INVx1_ASAP7_75t_L g11938 ( 
.A(n_11691),
.Y(n_11938)
);

INVx1_ASAP7_75t_L g11939 ( 
.A(n_11667),
.Y(n_11939)
);

HB1xp67_ASAP7_75t_L g11940 ( 
.A(n_11698),
.Y(n_11940)
);

INVx1_ASAP7_75t_L g11941 ( 
.A(n_11698),
.Y(n_11941)
);

AOI21x1_ASAP7_75t_L g11942 ( 
.A1(n_11633),
.A2(n_1620),
.B(n_1621),
.Y(n_11942)
);

INVx6_ASAP7_75t_L g11943 ( 
.A(n_11632),
.Y(n_11943)
);

INVx1_ASAP7_75t_L g11944 ( 
.A(n_11692),
.Y(n_11944)
);

INVx1_ASAP7_75t_L g11945 ( 
.A(n_11819),
.Y(n_11945)
);

INVx5_ASAP7_75t_L g11946 ( 
.A(n_11551),
.Y(n_11946)
);

NOR2xp33_ASAP7_75t_L g11947 ( 
.A(n_11673),
.B(n_1622),
.Y(n_11947)
);

AND2x2_ASAP7_75t_L g11948 ( 
.A(n_11780),
.B(n_1622),
.Y(n_11948)
);

BUFx2_ASAP7_75t_L g11949 ( 
.A(n_11696),
.Y(n_11949)
);

INVx3_ASAP7_75t_L g11950 ( 
.A(n_11705),
.Y(n_11950)
);

AND2x2_ASAP7_75t_L g11951 ( 
.A(n_11539),
.B(n_1623),
.Y(n_11951)
);

AO31x2_ASAP7_75t_L g11952 ( 
.A1(n_11651),
.A2(n_1627),
.A3(n_1625),
.B(n_1626),
.Y(n_11952)
);

INVx3_ASAP7_75t_L g11953 ( 
.A(n_11629),
.Y(n_11953)
);

INVx1_ASAP7_75t_L g11954 ( 
.A(n_11819),
.Y(n_11954)
);

INVx2_ASAP7_75t_L g11955 ( 
.A(n_11630),
.Y(n_11955)
);

INVx1_ASAP7_75t_L g11956 ( 
.A(n_11773),
.Y(n_11956)
);

BUFx3_ASAP7_75t_L g11957 ( 
.A(n_11739),
.Y(n_11957)
);

INVx1_ASAP7_75t_L g11958 ( 
.A(n_11552),
.Y(n_11958)
);

INVx1_ASAP7_75t_L g11959 ( 
.A(n_11550),
.Y(n_11959)
);

INVx2_ASAP7_75t_SL g11960 ( 
.A(n_11574),
.Y(n_11960)
);

BUFx6f_ASAP7_75t_L g11961 ( 
.A(n_11741),
.Y(n_11961)
);

INVx1_ASAP7_75t_L g11962 ( 
.A(n_11711),
.Y(n_11962)
);

INVx1_ASAP7_75t_SL g11963 ( 
.A(n_11806),
.Y(n_11963)
);

INVx1_ASAP7_75t_L g11964 ( 
.A(n_11591),
.Y(n_11964)
);

INVx2_ASAP7_75t_L g11965 ( 
.A(n_11657),
.Y(n_11965)
);

INVx2_ASAP7_75t_L g11966 ( 
.A(n_11694),
.Y(n_11966)
);

INVx2_ASAP7_75t_L g11967 ( 
.A(n_11694),
.Y(n_11967)
);

AND2x2_ASAP7_75t_L g11968 ( 
.A(n_11596),
.B(n_11569),
.Y(n_11968)
);

BUFx2_ASAP7_75t_L g11969 ( 
.A(n_11551),
.Y(n_11969)
);

INVx1_ASAP7_75t_L g11970 ( 
.A(n_11822),
.Y(n_11970)
);

AOI21x1_ASAP7_75t_L g11971 ( 
.A1(n_11680),
.A2(n_1626),
.B(n_1627),
.Y(n_11971)
);

INVx1_ASAP7_75t_L g11972 ( 
.A(n_11822),
.Y(n_11972)
);

OA21x2_ASAP7_75t_L g11973 ( 
.A1(n_11849),
.A2(n_11686),
.B(n_11755),
.Y(n_11973)
);

INVx1_ASAP7_75t_L g11974 ( 
.A(n_11826),
.Y(n_11974)
);

INVx2_ASAP7_75t_L g11975 ( 
.A(n_11747),
.Y(n_11975)
);

BUFx6f_ASAP7_75t_L g11976 ( 
.A(n_11745),
.Y(n_11976)
);

AO21x2_ASAP7_75t_L g11977 ( 
.A1(n_11603),
.A2(n_1628),
.B(n_1629),
.Y(n_11977)
);

AND2x2_ASAP7_75t_L g11978 ( 
.A(n_11568),
.B(n_1630),
.Y(n_11978)
);

INVx2_ASAP7_75t_L g11979 ( 
.A(n_11804),
.Y(n_11979)
);

INVx3_ASAP7_75t_L g11980 ( 
.A(n_11845),
.Y(n_11980)
);

INVx2_ASAP7_75t_L g11981 ( 
.A(n_11805),
.Y(n_11981)
);

INVx5_ASAP7_75t_SL g11982 ( 
.A(n_11821),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_11826),
.Y(n_11983)
);

BUFx3_ASAP7_75t_L g11984 ( 
.A(n_11689),
.Y(n_11984)
);

INVx2_ASAP7_75t_L g11985 ( 
.A(n_11818),
.Y(n_11985)
);

INVx2_ASAP7_75t_L g11986 ( 
.A(n_11820),
.Y(n_11986)
);

INVx1_ASAP7_75t_L g11987 ( 
.A(n_11710),
.Y(n_11987)
);

CKINVDCx5p33_ASAP7_75t_R g11988 ( 
.A(n_11637),
.Y(n_11988)
);

AOI22xp33_ASAP7_75t_L g11989 ( 
.A1(n_11601),
.A2(n_1632),
.B1(n_1630),
.B2(n_1631),
.Y(n_11989)
);

HB1xp67_ASAP7_75t_L g11990 ( 
.A(n_11583),
.Y(n_11990)
);

INVx1_ASAP7_75t_L g11991 ( 
.A(n_11731),
.Y(n_11991)
);

INVx2_ASAP7_75t_L g11992 ( 
.A(n_11554),
.Y(n_11992)
);

INVx1_ASAP7_75t_L g11993 ( 
.A(n_11714),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_11722),
.Y(n_11994)
);

INVx2_ASAP7_75t_L g11995 ( 
.A(n_11583),
.Y(n_11995)
);

INVx1_ASAP7_75t_L g11996 ( 
.A(n_11811),
.Y(n_11996)
);

INVx2_ASAP7_75t_L g11997 ( 
.A(n_11612),
.Y(n_11997)
);

INVx1_ASAP7_75t_L g11998 ( 
.A(n_11813),
.Y(n_11998)
);

BUFx3_ASAP7_75t_L g11999 ( 
.A(n_11737),
.Y(n_11999)
);

AND2x4_ASAP7_75t_SL g12000 ( 
.A(n_11535),
.B(n_1631),
.Y(n_12000)
);

OR2x2_ASAP7_75t_L g12001 ( 
.A(n_11768),
.B(n_1633),
.Y(n_12001)
);

OA21x2_ASAP7_75t_L g12002 ( 
.A1(n_11687),
.A2(n_1633),
.B(n_1634),
.Y(n_12002)
);

AO21x2_ASAP7_75t_L g12003 ( 
.A1(n_11558),
.A2(n_1634),
.B(n_1635),
.Y(n_12003)
);

INVx1_ASAP7_75t_L g12004 ( 
.A(n_11817),
.Y(n_12004)
);

AND2x2_ASAP7_75t_L g12005 ( 
.A(n_11770),
.B(n_1635),
.Y(n_12005)
);

INVx2_ASAP7_75t_L g12006 ( 
.A(n_11749),
.Y(n_12006)
);

INVx1_ASAP7_75t_L g12007 ( 
.A(n_11839),
.Y(n_12007)
);

INVx1_ASAP7_75t_L g12008 ( 
.A(n_11788),
.Y(n_12008)
);

INVx2_ASAP7_75t_L g12009 ( 
.A(n_11754),
.Y(n_12009)
);

AND2x2_ASAP7_75t_L g12010 ( 
.A(n_11832),
.B(n_1636),
.Y(n_12010)
);

INVx1_ASAP7_75t_L g12011 ( 
.A(n_11798),
.Y(n_12011)
);

INVx2_ASAP7_75t_L g12012 ( 
.A(n_11654),
.Y(n_12012)
);

INVx1_ASAP7_75t_L g12013 ( 
.A(n_11724),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_11585),
.Y(n_12014)
);

INVx4_ASAP7_75t_SL g12015 ( 
.A(n_11592),
.Y(n_12015)
);

INVx1_ASAP7_75t_L g12016 ( 
.A(n_11724),
.Y(n_12016)
);

INVx1_ASAP7_75t_L g12017 ( 
.A(n_11544),
.Y(n_12017)
);

INVxp67_ASAP7_75t_L g12018 ( 
.A(n_11645),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_11777),
.Y(n_12019)
);

INVx1_ASAP7_75t_L g12020 ( 
.A(n_11537),
.Y(n_12020)
);

INVx2_ASAP7_75t_L g12021 ( 
.A(n_11606),
.Y(n_12021)
);

INVx2_ASAP7_75t_L g12022 ( 
.A(n_11608),
.Y(n_12022)
);

INVx2_ASAP7_75t_L g12023 ( 
.A(n_11702),
.Y(n_12023)
);

INVx1_ASAP7_75t_L g12024 ( 
.A(n_11841),
.Y(n_12024)
);

AND2x2_ASAP7_75t_L g12025 ( 
.A(n_11613),
.B(n_1636),
.Y(n_12025)
);

INVx1_ASAP7_75t_L g12026 ( 
.A(n_11848),
.Y(n_12026)
);

INVx2_ASAP7_75t_L g12027 ( 
.A(n_11581),
.Y(n_12027)
);

BUFx2_ASAP7_75t_L g12028 ( 
.A(n_11816),
.Y(n_12028)
);

INVx1_ASAP7_75t_L g12029 ( 
.A(n_11854),
.Y(n_12029)
);

INVx2_ASAP7_75t_L g12030 ( 
.A(n_11598),
.Y(n_12030)
);

INVx2_ASAP7_75t_L g12031 ( 
.A(n_11618),
.Y(n_12031)
);

OR2x2_ASAP7_75t_L g12032 ( 
.A(n_11548),
.B(n_1637),
.Y(n_12032)
);

AND2x2_ASAP7_75t_L g12033 ( 
.A(n_11658),
.B(n_1638),
.Y(n_12033)
);

INVx1_ASAP7_75t_L g12034 ( 
.A(n_11794),
.Y(n_12034)
);

INVx1_ASAP7_75t_L g12035 ( 
.A(n_11792),
.Y(n_12035)
);

OAI21xp5_ASAP7_75t_L g12036 ( 
.A1(n_11557),
.A2(n_1638),
.B(n_1639),
.Y(n_12036)
);

AND2x4_ASAP7_75t_L g12037 ( 
.A(n_11570),
.B(n_1639),
.Y(n_12037)
);

AO21x1_ASAP7_75t_SL g12038 ( 
.A1(n_11543),
.A2(n_1640),
.B(n_1642),
.Y(n_12038)
);

AO31x2_ASAP7_75t_L g12039 ( 
.A1(n_11553),
.A2(n_1643),
.A3(n_1640),
.B(n_1642),
.Y(n_12039)
);

BUFx6f_ASAP7_75t_L g12040 ( 
.A(n_11742),
.Y(n_12040)
);

INVx3_ASAP7_75t_L g12041 ( 
.A(n_11556),
.Y(n_12041)
);

BUFx2_ASAP7_75t_L g12042 ( 
.A(n_11743),
.Y(n_12042)
);

OAI22xp33_ASAP7_75t_L g12043 ( 
.A1(n_11663),
.A2(n_1645),
.B1(n_1643),
.B2(n_1644),
.Y(n_12043)
);

AND2x2_ASAP7_75t_L g12044 ( 
.A(n_11844),
.B(n_1645),
.Y(n_12044)
);

HB1xp67_ASAP7_75t_L g12045 ( 
.A(n_11655),
.Y(n_12045)
);

INVx2_ASAP7_75t_L g12046 ( 
.A(n_11648),
.Y(n_12046)
);

AND2x2_ASAP7_75t_L g12047 ( 
.A(n_11852),
.B(n_1646),
.Y(n_12047)
);

OR2x2_ASAP7_75t_L g12048 ( 
.A(n_11855),
.B(n_1646),
.Y(n_12048)
);

BUFx6f_ASAP7_75t_L g12049 ( 
.A(n_11746),
.Y(n_12049)
);

INVx3_ASAP7_75t_L g12050 ( 
.A(n_11653),
.Y(n_12050)
);

INVx2_ASAP7_75t_L g12051 ( 
.A(n_11831),
.Y(n_12051)
);

INVx2_ASAP7_75t_L g12052 ( 
.A(n_11611),
.Y(n_12052)
);

INVx1_ASAP7_75t_L g12053 ( 
.A(n_11792),
.Y(n_12053)
);

INVx1_ASAP7_75t_L g12054 ( 
.A(n_11561),
.Y(n_12054)
);

AND2x2_ASAP7_75t_L g12055 ( 
.A(n_11853),
.B(n_1647),
.Y(n_12055)
);

INVx1_ASAP7_75t_L g12056 ( 
.A(n_11668),
.Y(n_12056)
);

NOR2xp33_ASAP7_75t_L g12057 ( 
.A(n_11785),
.B(n_1647),
.Y(n_12057)
);

INVx1_ASAP7_75t_L g12058 ( 
.A(n_11793),
.Y(n_12058)
);

HB1xp67_ASAP7_75t_L g12059 ( 
.A(n_11838),
.Y(n_12059)
);

BUFx2_ASAP7_75t_L g12060 ( 
.A(n_11647),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11824),
.Y(n_12061)
);

AO21x2_ASAP7_75t_L g12062 ( 
.A1(n_11627),
.A2(n_1648),
.B(n_1649),
.Y(n_12062)
);

INVx4_ASAP7_75t_SL g12063 ( 
.A(n_11716),
.Y(n_12063)
);

AND2x2_ASAP7_75t_L g12064 ( 
.A(n_11859),
.B(n_1648),
.Y(n_12064)
);

BUFx2_ASAP7_75t_L g12065 ( 
.A(n_11588),
.Y(n_12065)
);

AND2x4_ASAP7_75t_L g12066 ( 
.A(n_11670),
.B(n_1650),
.Y(n_12066)
);

INVx2_ASAP7_75t_L g12067 ( 
.A(n_11610),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_11802),
.Y(n_12068)
);

BUFx2_ASAP7_75t_L g12069 ( 
.A(n_11802),
.Y(n_12069)
);

INVx1_ASAP7_75t_L g12070 ( 
.A(n_11665),
.Y(n_12070)
);

AND2x4_ASAP7_75t_SL g12071 ( 
.A(n_11781),
.B(n_1650),
.Y(n_12071)
);

INVx2_ASAP7_75t_L g12072 ( 
.A(n_11744),
.Y(n_12072)
);

BUFx6f_ASAP7_75t_L g12073 ( 
.A(n_11764),
.Y(n_12073)
);

INVx1_ASAP7_75t_L g12074 ( 
.A(n_11675),
.Y(n_12074)
);

OA21x2_ASAP7_75t_L g12075 ( 
.A1(n_11695),
.A2(n_1651),
.B(n_1652),
.Y(n_12075)
);

AND2x2_ASAP7_75t_L g12076 ( 
.A(n_11719),
.B(n_1651),
.Y(n_12076)
);

OAI21x1_ASAP7_75t_L g12077 ( 
.A1(n_11536),
.A2(n_1652),
.B(n_1653),
.Y(n_12077)
);

INVx2_ASAP7_75t_L g12078 ( 
.A(n_11707),
.Y(n_12078)
);

AND2x4_ASAP7_75t_L g12079 ( 
.A(n_11712),
.B(n_1653),
.Y(n_12079)
);

OR2x2_ASAP7_75t_L g12080 ( 
.A(n_11614),
.B(n_1654),
.Y(n_12080)
);

INVx1_ASAP7_75t_L g12081 ( 
.A(n_11616),
.Y(n_12081)
);

INVx1_ASAP7_75t_L g12082 ( 
.A(n_11621),
.Y(n_12082)
);

AND2x4_ASAP7_75t_L g12083 ( 
.A(n_11808),
.B(n_1654),
.Y(n_12083)
);

INVx2_ASAP7_75t_L g12084 ( 
.A(n_11605),
.Y(n_12084)
);

INVx2_ASAP7_75t_L g12085 ( 
.A(n_11835),
.Y(n_12085)
);

INVx1_ASAP7_75t_L g12086 ( 
.A(n_11791),
.Y(n_12086)
);

AND2x2_ASAP7_75t_L g12087 ( 
.A(n_11752),
.B(n_1655),
.Y(n_12087)
);

HB1xp67_ASAP7_75t_L g12088 ( 
.A(n_11547),
.Y(n_12088)
);

INVx1_ASAP7_75t_L g12089 ( 
.A(n_11562),
.Y(n_12089)
);

AOI21xp5_ASAP7_75t_SL g12090 ( 
.A1(n_11567),
.A2(n_11718),
.B(n_11720),
.Y(n_12090)
);

OAI21x1_ASAP7_75t_L g12091 ( 
.A1(n_11656),
.A2(n_11730),
.B(n_11650),
.Y(n_12091)
);

INVx2_ASAP7_75t_SL g12092 ( 
.A(n_11762),
.Y(n_12092)
);

AND2x2_ASAP7_75t_L g12093 ( 
.A(n_11796),
.B(n_1656),
.Y(n_12093)
);

NAND2x1p5_ASAP7_75t_L g12094 ( 
.A(n_11812),
.B(n_1656),
.Y(n_12094)
);

INVx2_ASAP7_75t_SL g12095 ( 
.A(n_11846),
.Y(n_12095)
);

INVx2_ASAP7_75t_L g12096 ( 
.A(n_11837),
.Y(n_12096)
);

INVx3_ASAP7_75t_L g12097 ( 
.A(n_11809),
.Y(n_12097)
);

AND2x4_ASAP7_75t_L g12098 ( 
.A(n_11693),
.B(n_1657),
.Y(n_12098)
);

AND2x2_ASAP7_75t_L g12099 ( 
.A(n_11728),
.B(n_11646),
.Y(n_12099)
);

OR2x2_ASAP7_75t_L g12100 ( 
.A(n_11784),
.B(n_1657),
.Y(n_12100)
);

AND2x2_ASAP7_75t_L g12101 ( 
.A(n_11823),
.B(n_1658),
.Y(n_12101)
);

NAND2xp5_ASAP7_75t_L g12102 ( 
.A(n_11704),
.B(n_1658),
.Y(n_12102)
);

NAND2x1p5_ASAP7_75t_L g12103 ( 
.A(n_11577),
.B(n_1659),
.Y(n_12103)
);

HB1xp67_ASAP7_75t_L g12104 ( 
.A(n_11690),
.Y(n_12104)
);

OAI21x1_ASAP7_75t_L g12105 ( 
.A1(n_11843),
.A2(n_1659),
.B(n_1660),
.Y(n_12105)
);

INVx2_ASAP7_75t_L g12106 ( 
.A(n_11757),
.Y(n_12106)
);

BUFx4f_ASAP7_75t_SL g12107 ( 
.A(n_11639),
.Y(n_12107)
);

BUFx3_ASAP7_75t_L g12108 ( 
.A(n_11700),
.Y(n_12108)
);

INVx3_ASAP7_75t_L g12109 ( 
.A(n_11701),
.Y(n_12109)
);

INVx1_ASAP7_75t_L g12110 ( 
.A(n_11829),
.Y(n_12110)
);

INVx1_ASAP7_75t_L g12111 ( 
.A(n_11738),
.Y(n_12111)
);

INVx1_ASAP7_75t_L g12112 ( 
.A(n_11589),
.Y(n_12112)
);

AOI21x1_ASAP7_75t_L g12113 ( 
.A1(n_11640),
.A2(n_1660),
.B(n_1661),
.Y(n_12113)
);

INVx2_ASAP7_75t_SL g12114 ( 
.A(n_11795),
.Y(n_12114)
);

AND2x2_ASAP7_75t_L g12115 ( 
.A(n_11622),
.B(n_1662),
.Y(n_12115)
);

AO21x2_ASAP7_75t_L g12116 ( 
.A1(n_11753),
.A2(n_1662),
.B(n_1663),
.Y(n_12116)
);

INVx2_ASAP7_75t_L g12117 ( 
.A(n_11666),
.Y(n_12117)
);

AND2x2_ASAP7_75t_L g12118 ( 
.A(n_11717),
.B(n_1664),
.Y(n_12118)
);

OA21x2_ASAP7_75t_L g12119 ( 
.A1(n_11619),
.A2(n_1664),
.B(n_1665),
.Y(n_12119)
);

INVx1_ASAP7_75t_L g12120 ( 
.A(n_11750),
.Y(n_12120)
);

INVx1_ASAP7_75t_L g12121 ( 
.A(n_11708),
.Y(n_12121)
);

INVx1_ASAP7_75t_L g12122 ( 
.A(n_11751),
.Y(n_12122)
);

INVx1_ASAP7_75t_L g12123 ( 
.A(n_11726),
.Y(n_12123)
);

AND2x2_ASAP7_75t_L g12124 ( 
.A(n_11721),
.B(n_1666),
.Y(n_12124)
);

INVx3_ASAP7_75t_L g12125 ( 
.A(n_11827),
.Y(n_12125)
);

OAI21x1_ASAP7_75t_L g12126 ( 
.A1(n_11584),
.A2(n_1667),
.B(n_1668),
.Y(n_12126)
);

AND2x2_ASAP7_75t_L g12127 ( 
.A(n_11790),
.B(n_1669),
.Y(n_12127)
);

OR2x2_ASAP7_75t_L g12128 ( 
.A(n_11576),
.B(n_1669),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11834),
.Y(n_12129)
);

INVx2_ASAP7_75t_L g12130 ( 
.A(n_11559),
.Y(n_12130)
);

INVx2_ASAP7_75t_L g12131 ( 
.A(n_11772),
.Y(n_12131)
);

OAI21x1_ASAP7_75t_L g12132 ( 
.A1(n_11586),
.A2(n_1670),
.B(n_1672),
.Y(n_12132)
);

AO21x2_ASAP7_75t_L g12133 ( 
.A1(n_11851),
.A2(n_1673),
.B(n_1674),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_11760),
.Y(n_12134)
);

AND2x2_ASAP7_75t_L g12135 ( 
.A(n_11595),
.B(n_1673),
.Y(n_12135)
);

INVx3_ASAP7_75t_L g12136 ( 
.A(n_11572),
.Y(n_12136)
);

INVx1_ASAP7_75t_L g12137 ( 
.A(n_11533),
.Y(n_12137)
);

AO21x1_ASAP7_75t_SL g12138 ( 
.A1(n_11858),
.A2(n_1674),
.B(n_1675),
.Y(n_12138)
);

AND2x4_ASAP7_75t_L g12139 ( 
.A(n_11763),
.B(n_1675),
.Y(n_12139)
);

HB1xp67_ASAP7_75t_L g12140 ( 
.A(n_11649),
.Y(n_12140)
);

AND2x2_ASAP7_75t_L g12141 ( 
.A(n_11593),
.B(n_11833),
.Y(n_12141)
);

INVx2_ASAP7_75t_L g12142 ( 
.A(n_11850),
.Y(n_12142)
);

INVx1_ASAP7_75t_L g12143 ( 
.A(n_11825),
.Y(n_12143)
);

NAND2xp5_ASAP7_75t_L g12144 ( 
.A(n_11626),
.B(n_1676),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_11828),
.B(n_1676),
.Y(n_12145)
);

BUFx2_ASAP7_75t_L g12146 ( 
.A(n_11801),
.Y(n_12146)
);

INVx1_ASAP7_75t_L g12147 ( 
.A(n_11783),
.Y(n_12147)
);

HB1xp67_ASAP7_75t_L g12148 ( 
.A(n_11836),
.Y(n_12148)
);

OAI21x1_ASAP7_75t_L g12149 ( 
.A1(n_11600),
.A2(n_1677),
.B(n_1679),
.Y(n_12149)
);

INVx3_ASAP7_75t_L g12150 ( 
.A(n_11797),
.Y(n_12150)
);

AOI22xp33_ASAP7_75t_L g12151 ( 
.A1(n_11531),
.A2(n_1680),
.B1(n_1677),
.B2(n_1679),
.Y(n_12151)
);

INVx1_ASAP7_75t_L g12152 ( 
.A(n_11674),
.Y(n_12152)
);

INVx1_ASAP7_75t_L g12153 ( 
.A(n_11767),
.Y(n_12153)
);

AND2x2_ASAP7_75t_L g12154 ( 
.A(n_11756),
.B(n_1680),
.Y(n_12154)
);

AO21x2_ASAP7_75t_L g12155 ( 
.A1(n_11676),
.A2(n_1681),
.B(n_1682),
.Y(n_12155)
);

HB1xp67_ASAP7_75t_L g12156 ( 
.A(n_11736),
.Y(n_12156)
);

INVx2_ASAP7_75t_L g12157 ( 
.A(n_11814),
.Y(n_12157)
);

OA21x2_ASAP7_75t_L g12158 ( 
.A1(n_11678),
.A2(n_1682),
.B(n_1683),
.Y(n_12158)
);

INVx2_ASAP7_75t_L g12159 ( 
.A(n_11579),
.Y(n_12159)
);

INVx1_ASAP7_75t_L g12160 ( 
.A(n_11758),
.Y(n_12160)
);

OAI21xp5_ASAP7_75t_L g12161 ( 
.A1(n_11540),
.A2(n_11840),
.B(n_11856),
.Y(n_12161)
);

OAI21x1_ASAP7_75t_L g12162 ( 
.A1(n_11786),
.A2(n_1684),
.B(n_1685),
.Y(n_12162)
);

INVx2_ASAP7_75t_L g12163 ( 
.A(n_11769),
.Y(n_12163)
);

OAI22xp33_ASAP7_75t_L g12164 ( 
.A1(n_11609),
.A2(n_1687),
.B1(n_1685),
.B2(n_1686),
.Y(n_12164)
);

HB1xp67_ASAP7_75t_L g12165 ( 
.A(n_11800),
.Y(n_12165)
);

AND2x2_ASAP7_75t_L g12166 ( 
.A(n_11761),
.B(n_1687),
.Y(n_12166)
);

INVx2_ASAP7_75t_L g12167 ( 
.A(n_11807),
.Y(n_12167)
);

INVx2_ASAP7_75t_L g12168 ( 
.A(n_11594),
.Y(n_12168)
);

INVx1_ASAP7_75t_L g12169 ( 
.A(n_11815),
.Y(n_12169)
);

BUFx3_ASAP7_75t_L g12170 ( 
.A(n_11765),
.Y(n_12170)
);

INVx2_ASAP7_75t_L g12171 ( 
.A(n_11778),
.Y(n_12171)
);

BUFx6f_ASAP7_75t_L g12172 ( 
.A(n_11782),
.Y(n_12172)
);

AND2x2_ASAP7_75t_L g12173 ( 
.A(n_11590),
.B(n_11688),
.Y(n_12173)
);

AO21x2_ASAP7_75t_L g12174 ( 
.A1(n_11789),
.A2(n_1688),
.B(n_1689),
.Y(n_12174)
);

HB1xp67_ASAP7_75t_L g12175 ( 
.A(n_11759),
.Y(n_12175)
);

INVx2_ASAP7_75t_L g12176 ( 
.A(n_11697),
.Y(n_12176)
);

CKINVDCx5p33_ASAP7_75t_R g12177 ( 
.A(n_11555),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_11803),
.Y(n_12178)
);

INVx3_ASAP7_75t_L g12179 ( 
.A(n_11740),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11748),
.Y(n_12180)
);

OR2x2_ASAP7_75t_L g12181 ( 
.A(n_11642),
.B(n_1688),
.Y(n_12181)
);

INVx2_ASAP7_75t_L g12182 ( 
.A(n_11713),
.Y(n_12182)
);

OAI21x1_ASAP7_75t_L g12183 ( 
.A1(n_11766),
.A2(n_1689),
.B(n_1690),
.Y(n_12183)
);

INVx1_ASAP7_75t_L g12184 ( 
.A(n_11775),
.Y(n_12184)
);

AND2x2_ASAP7_75t_L g12185 ( 
.A(n_11732),
.B(n_1690),
.Y(n_12185)
);

OAI21xp5_ASAP7_75t_L g12186 ( 
.A1(n_11636),
.A2(n_1691),
.B(n_1692),
.Y(n_12186)
);

INVx3_ASAP7_75t_L g12187 ( 
.A(n_11560),
.Y(n_12187)
);

AO21x2_ASAP7_75t_L g12188 ( 
.A1(n_11641),
.A2(n_1692),
.B(n_1694),
.Y(n_12188)
);

INVx2_ASAP7_75t_L g12189 ( 
.A(n_11830),
.Y(n_12189)
);

BUFx3_ASAP7_75t_L g12190 ( 
.A(n_11624),
.Y(n_12190)
);

BUFx2_ASAP7_75t_L g12191 ( 
.A(n_11631),
.Y(n_12191)
);

AND2x2_ASAP7_75t_L g12192 ( 
.A(n_11652),
.B(n_1694),
.Y(n_12192)
);

INVx5_ASAP7_75t_SL g12193 ( 
.A(n_11857),
.Y(n_12193)
);

INVx1_ASAP7_75t_L g12194 ( 
.A(n_11659),
.Y(n_12194)
);

INVx1_ASAP7_75t_L g12195 ( 
.A(n_11659),
.Y(n_12195)
);

INVx1_ASAP7_75t_L g12196 ( 
.A(n_11659),
.Y(n_12196)
);

INVx3_ASAP7_75t_L g12197 ( 
.A(n_11549),
.Y(n_12197)
);

OAI21xp5_ASAP7_75t_L g12198 ( 
.A1(n_12091),
.A2(n_1695),
.B(n_1696),
.Y(n_12198)
);

AND2x4_ASAP7_75t_L g12199 ( 
.A(n_11862),
.B(n_1696),
.Y(n_12199)
);

AND2x2_ASAP7_75t_L g12200 ( 
.A(n_11867),
.B(n_1697),
.Y(n_12200)
);

NAND2xp5_ASAP7_75t_L g12201 ( 
.A(n_12095),
.B(n_1698),
.Y(n_12201)
);

AOI22xp5_ASAP7_75t_L g12202 ( 
.A1(n_12146),
.A2(n_1702),
.B1(n_1699),
.B2(n_1700),
.Y(n_12202)
);

INVx2_ASAP7_75t_L g12203 ( 
.A(n_11901),
.Y(n_12203)
);

INVx5_ASAP7_75t_L g12204 ( 
.A(n_12193),
.Y(n_12204)
);

AND2x2_ASAP7_75t_L g12205 ( 
.A(n_12015),
.B(n_1699),
.Y(n_12205)
);

OR2x2_ASAP7_75t_L g12206 ( 
.A(n_12072),
.B(n_1700),
.Y(n_12206)
);

INVx4_ASAP7_75t_L g12207 ( 
.A(n_11894),
.Y(n_12207)
);

A2O1A1Ixp33_ASAP7_75t_L g12208 ( 
.A1(n_12191),
.A2(n_1704),
.B(n_1702),
.C(n_1703),
.Y(n_12208)
);

OAI21xp5_ASAP7_75t_L g12209 ( 
.A1(n_12161),
.A2(n_12090),
.B(n_12125),
.Y(n_12209)
);

INVx2_ASAP7_75t_L g12210 ( 
.A(n_11901),
.Y(n_12210)
);

OR2x2_ASAP7_75t_L g12211 ( 
.A(n_12034),
.B(n_1703),
.Y(n_12211)
);

BUFx6f_ASAP7_75t_L g12212 ( 
.A(n_11893),
.Y(n_12212)
);

OAI21x1_ASAP7_75t_L g12213 ( 
.A1(n_11928),
.A2(n_12078),
.B(n_11876),
.Y(n_12213)
);

O2A1O1Ixp33_ASAP7_75t_L g12214 ( 
.A1(n_11887),
.A2(n_1707),
.B(n_1705),
.C(n_1706),
.Y(n_12214)
);

OR2x2_ASAP7_75t_L g12215 ( 
.A(n_11949),
.B(n_1705),
.Y(n_12215)
);

OR2x2_ASAP7_75t_L g12216 ( 
.A(n_12014),
.B(n_1706),
.Y(n_12216)
);

OR2x2_ASAP7_75t_L g12217 ( 
.A(n_12008),
.B(n_1707),
.Y(n_12217)
);

NAND2xp5_ASAP7_75t_L g12218 ( 
.A(n_11930),
.B(n_1708),
.Y(n_12218)
);

OAI21xp5_ASAP7_75t_L g12219 ( 
.A1(n_12112),
.A2(n_1709),
.B(n_1710),
.Y(n_12219)
);

O2A1O1Ixp33_ASAP7_75t_SL g12220 ( 
.A1(n_11890),
.A2(n_1712),
.B(n_1709),
.C(n_1711),
.Y(n_12220)
);

BUFx2_ASAP7_75t_L g12221 ( 
.A(n_11869),
.Y(n_12221)
);

AND2x2_ASAP7_75t_L g12222 ( 
.A(n_11922),
.B(n_1711),
.Y(n_12222)
);

OAI21xp5_ASAP7_75t_L g12223 ( 
.A1(n_12173),
.A2(n_1712),
.B(n_1713),
.Y(n_12223)
);

AND2x2_ASAP7_75t_L g12224 ( 
.A(n_11891),
.B(n_1713),
.Y(n_12224)
);

OR2x2_ASAP7_75t_L g12225 ( 
.A(n_12012),
.B(n_1714),
.Y(n_12225)
);

BUFx3_ASAP7_75t_L g12226 ( 
.A(n_12197),
.Y(n_12226)
);

BUFx2_ASAP7_75t_L g12227 ( 
.A(n_11969),
.Y(n_12227)
);

AND2x2_ASAP7_75t_L g12228 ( 
.A(n_11916),
.B(n_1714),
.Y(n_12228)
);

NOR2xp33_ASAP7_75t_L g12229 ( 
.A(n_11888),
.B(n_1715),
.Y(n_12229)
);

AND2x2_ASAP7_75t_L g12230 ( 
.A(n_11921),
.B(n_1715),
.Y(n_12230)
);

AND2x2_ASAP7_75t_L g12231 ( 
.A(n_11950),
.B(n_1716),
.Y(n_12231)
);

A2O1A1Ixp33_ASAP7_75t_L g12232 ( 
.A1(n_12190),
.A2(n_12179),
.B(n_12157),
.C(n_12117),
.Y(n_12232)
);

INVx1_ASAP7_75t_L g12233 ( 
.A(n_11864),
.Y(n_12233)
);

AND2x2_ASAP7_75t_L g12234 ( 
.A(n_11915),
.B(n_1716),
.Y(n_12234)
);

AND2x2_ASAP7_75t_L g12235 ( 
.A(n_11897),
.B(n_1717),
.Y(n_12235)
);

OR2x2_ASAP7_75t_L g12236 ( 
.A(n_12061),
.B(n_1718),
.Y(n_12236)
);

AND2x2_ASAP7_75t_L g12237 ( 
.A(n_11880),
.B(n_11889),
.Y(n_12237)
);

A2O1A1Ixp33_ASAP7_75t_L g12238 ( 
.A1(n_12187),
.A2(n_1720),
.B(n_1718),
.C(n_1719),
.Y(n_12238)
);

AO32x1_ASAP7_75t_L g12239 ( 
.A1(n_12129),
.A2(n_1722),
.A3(n_1719),
.B1(n_1721),
.B2(n_1723),
.Y(n_12239)
);

OA21x2_ASAP7_75t_L g12240 ( 
.A1(n_11913),
.A2(n_11911),
.B(n_11909),
.Y(n_12240)
);

HB1xp67_ASAP7_75t_L g12241 ( 
.A(n_12059),
.Y(n_12241)
);

AOI211xp5_ASAP7_75t_L g12242 ( 
.A1(n_12186),
.A2(n_1726),
.B(n_1721),
.C(n_1724),
.Y(n_12242)
);

O2A1O1Ixp33_ASAP7_75t_L g12243 ( 
.A1(n_11868),
.A2(n_1727),
.B(n_1724),
.C(n_1726),
.Y(n_12243)
);

OR2x2_ASAP7_75t_L g12244 ( 
.A(n_12051),
.B(n_1728),
.Y(n_12244)
);

INVx1_ASAP7_75t_L g12245 ( 
.A(n_11872),
.Y(n_12245)
);

O2A1O1Ixp33_ASAP7_75t_L g12246 ( 
.A1(n_12142),
.A2(n_1731),
.B(n_1729),
.C(n_1730),
.Y(n_12246)
);

HB1xp67_ASAP7_75t_L g12247 ( 
.A(n_11882),
.Y(n_12247)
);

OAI22xp5_ASAP7_75t_L g12248 ( 
.A1(n_12177),
.A2(n_12107),
.B1(n_12148),
.B2(n_11930),
.Y(n_12248)
);

NAND3xp33_ASAP7_75t_L g12249 ( 
.A(n_11904),
.B(n_1729),
.C(n_1730),
.Y(n_12249)
);

A2O1A1Ixp33_ASAP7_75t_L g12250 ( 
.A1(n_12131),
.A2(n_1734),
.B(n_1731),
.C(n_1733),
.Y(n_12250)
);

OR2x2_ASAP7_75t_L g12251 ( 
.A(n_11861),
.B(n_1733),
.Y(n_12251)
);

AND2x2_ASAP7_75t_L g12252 ( 
.A(n_11886),
.B(n_1734),
.Y(n_12252)
);

OA21x2_ASAP7_75t_L g12253 ( 
.A1(n_12018),
.A2(n_1735),
.B(n_1736),
.Y(n_12253)
);

NAND2xp5_ASAP7_75t_L g12254 ( 
.A(n_12130),
.B(n_1736),
.Y(n_12254)
);

INVx1_ASAP7_75t_L g12255 ( 
.A(n_11962),
.Y(n_12255)
);

A2O1A1Ixp33_ASAP7_75t_L g12256 ( 
.A1(n_12152),
.A2(n_1739),
.B(n_1737),
.C(n_1738),
.Y(n_12256)
);

AO32x2_ASAP7_75t_L g12257 ( 
.A1(n_11960),
.A2(n_1739),
.A3(n_1737),
.B1(n_1738),
.B2(n_1741),
.Y(n_12257)
);

HB1xp67_ASAP7_75t_L g12258 ( 
.A(n_12045),
.Y(n_12258)
);

NAND2xp5_ASAP7_75t_L g12259 ( 
.A(n_12159),
.B(n_1741),
.Y(n_12259)
);

INVx2_ASAP7_75t_L g12260 ( 
.A(n_11926),
.Y(n_12260)
);

O2A1O1Ixp33_ASAP7_75t_SL g12261 ( 
.A1(n_12144),
.A2(n_1744),
.B(n_1742),
.C(n_1743),
.Y(n_12261)
);

OAI22xp5_ASAP7_75t_L g12262 ( 
.A1(n_12120),
.A2(n_1744),
.B1(n_1742),
.B2(n_1743),
.Y(n_12262)
);

AOI21xp5_ASAP7_75t_L g12263 ( 
.A1(n_12137),
.A2(n_1745),
.B(n_1746),
.Y(n_12263)
);

BUFx6f_ASAP7_75t_L g12264 ( 
.A(n_11920),
.Y(n_12264)
);

AO21x2_ASAP7_75t_L g12265 ( 
.A1(n_11990),
.A2(n_1745),
.B(n_1747),
.Y(n_12265)
);

INVx2_ASAP7_75t_L g12266 ( 
.A(n_11926),
.Y(n_12266)
);

HB1xp67_ASAP7_75t_L g12267 ( 
.A(n_12042),
.Y(n_12267)
);

OAI21xp5_ASAP7_75t_L g12268 ( 
.A1(n_12143),
.A2(n_1748),
.B(n_1749),
.Y(n_12268)
);

OAI211xp5_ASAP7_75t_L g12269 ( 
.A1(n_11989),
.A2(n_1751),
.B(n_1749),
.C(n_1750),
.Y(n_12269)
);

AND2x2_ASAP7_75t_L g12270 ( 
.A(n_11917),
.B(n_1750),
.Y(n_12270)
);

AND2x2_ASAP7_75t_L g12271 ( 
.A(n_12060),
.B(n_1751),
.Y(n_12271)
);

AND2x2_ASAP7_75t_L g12272 ( 
.A(n_11902),
.B(n_1752),
.Y(n_12272)
);

OAI22xp5_ASAP7_75t_L g12273 ( 
.A1(n_12111),
.A2(n_1754),
.B1(n_1752),
.B2(n_1753),
.Y(n_12273)
);

AND2x2_ASAP7_75t_L g12274 ( 
.A(n_11884),
.B(n_1753),
.Y(n_12274)
);

NAND2x1p5_ASAP7_75t_L g12275 ( 
.A(n_11946),
.B(n_1755),
.Y(n_12275)
);

INVx3_ASAP7_75t_L g12276 ( 
.A(n_11961),
.Y(n_12276)
);

OAI21x1_ASAP7_75t_L g12277 ( 
.A1(n_11914),
.A2(n_1755),
.B(n_1756),
.Y(n_12277)
);

AND2x2_ASAP7_75t_L g12278 ( 
.A(n_12050),
.B(n_1756),
.Y(n_12278)
);

A2O1A1Ixp33_ASAP7_75t_L g12279 ( 
.A1(n_12150),
.A2(n_1759),
.B(n_1757),
.C(n_1758),
.Y(n_12279)
);

AOI221xp5_ASAP7_75t_L g12280 ( 
.A1(n_12134),
.A2(n_1760),
.B1(n_1758),
.B2(n_1759),
.C(n_1761),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_11956),
.Y(n_12281)
);

OAI22xp5_ASAP7_75t_SL g12282 ( 
.A1(n_11946),
.A2(n_1763),
.B1(n_1760),
.B2(n_1761),
.Y(n_12282)
);

INVx1_ASAP7_75t_L g12283 ( 
.A(n_11938),
.Y(n_12283)
);

NOR2x1_ASAP7_75t_SL g12284 ( 
.A(n_12138),
.B(n_1763),
.Y(n_12284)
);

AND2x2_ASAP7_75t_L g12285 ( 
.A(n_11910),
.B(n_1764),
.Y(n_12285)
);

OAI22xp5_ASAP7_75t_L g12286 ( 
.A1(n_12121),
.A2(n_1767),
.B1(n_1765),
.B2(n_1766),
.Y(n_12286)
);

AOI22xp33_ASAP7_75t_L g12287 ( 
.A1(n_12189),
.A2(n_1771),
.B1(n_1766),
.B2(n_1769),
.Y(n_12287)
);

AND2x4_ASAP7_75t_L g12288 ( 
.A(n_11905),
.B(n_1769),
.Y(n_12288)
);

AND2x2_ASAP7_75t_L g12289 ( 
.A(n_11955),
.B(n_1771),
.Y(n_12289)
);

INVx2_ASAP7_75t_L g12290 ( 
.A(n_11907),
.Y(n_12290)
);

OR2x2_ASAP7_75t_L g12291 ( 
.A(n_12052),
.B(n_1772),
.Y(n_12291)
);

AND2x4_ASAP7_75t_L g12292 ( 
.A(n_11963),
.B(n_1773),
.Y(n_12292)
);

INVx1_ASAP7_75t_L g12293 ( 
.A(n_11987),
.Y(n_12293)
);

OAI21xp5_ASAP7_75t_L g12294 ( 
.A1(n_12147),
.A2(n_1773),
.B(n_1774),
.Y(n_12294)
);

AND2x2_ASAP7_75t_L g12295 ( 
.A(n_11965),
.B(n_1774),
.Y(n_12295)
);

OR2x6_ASAP7_75t_L g12296 ( 
.A(n_12066),
.B(n_1775),
.Y(n_12296)
);

OR2x2_ASAP7_75t_L g12297 ( 
.A(n_12067),
.B(n_11939),
.Y(n_12297)
);

AND2x4_ASAP7_75t_L g12298 ( 
.A(n_11929),
.B(n_1776),
.Y(n_12298)
);

AO21x2_ASAP7_75t_L g12299 ( 
.A1(n_12013),
.A2(n_1776),
.B(n_1777),
.Y(n_12299)
);

AND2x2_ASAP7_75t_L g12300 ( 
.A(n_11892),
.B(n_1777),
.Y(n_12300)
);

OAI22xp5_ASAP7_75t_L g12301 ( 
.A1(n_12123),
.A2(n_1780),
.B1(n_1778),
.B2(n_1779),
.Y(n_12301)
);

AOI21xp5_ASAP7_75t_L g12302 ( 
.A1(n_12122),
.A2(n_1778),
.B(n_1780),
.Y(n_12302)
);

AND2x2_ASAP7_75t_L g12303 ( 
.A(n_12097),
.B(n_1781),
.Y(n_12303)
);

AND2x4_ASAP7_75t_SL g12304 ( 
.A(n_12041),
.B(n_1781),
.Y(n_12304)
);

OR2x2_ASAP7_75t_L g12305 ( 
.A(n_11958),
.B(n_1782),
.Y(n_12305)
);

INVx1_ASAP7_75t_L g12306 ( 
.A(n_11993),
.Y(n_12306)
);

OAI21x1_ASAP7_75t_L g12307 ( 
.A1(n_11863),
.A2(n_1782),
.B(n_1783),
.Y(n_12307)
);

AOI21xp5_ASAP7_75t_L g12308 ( 
.A1(n_12169),
.A2(n_1783),
.B(n_1784),
.Y(n_12308)
);

AND2x2_ASAP7_75t_L g12309 ( 
.A(n_11999),
.B(n_1784),
.Y(n_12309)
);

AND2x4_ASAP7_75t_L g12310 ( 
.A(n_11936),
.B(n_1785),
.Y(n_12310)
);

AND2x4_ASAP7_75t_L g12311 ( 
.A(n_11980),
.B(n_1785),
.Y(n_12311)
);

OA21x2_ASAP7_75t_L g12312 ( 
.A1(n_12069),
.A2(n_12016),
.B(n_11941),
.Y(n_12312)
);

OA21x2_ASAP7_75t_L g12313 ( 
.A1(n_11931),
.A2(n_1786),
.B(n_1787),
.Y(n_12313)
);

AND2x2_ASAP7_75t_L g12314 ( 
.A(n_11997),
.B(n_1786),
.Y(n_12314)
);

NAND2xp5_ASAP7_75t_L g12315 ( 
.A(n_12184),
.B(n_12182),
.Y(n_12315)
);

OAI21xp5_ASAP7_75t_L g12316 ( 
.A1(n_11860),
.A2(n_1787),
.B(n_1788),
.Y(n_12316)
);

NAND4xp25_ASAP7_75t_L g12317 ( 
.A(n_12028),
.B(n_1791),
.C(n_1789),
.D(n_1790),
.Y(n_12317)
);

INVx1_ASAP7_75t_L g12318 ( 
.A(n_11994),
.Y(n_12318)
);

OAI21xp5_ASAP7_75t_L g12319 ( 
.A1(n_12115),
.A2(n_1789),
.B(n_1790),
.Y(n_12319)
);

NAND2xp5_ASAP7_75t_L g12320 ( 
.A(n_12180),
.B(n_1791),
.Y(n_12320)
);

AOI22xp5_ASAP7_75t_L g12321 ( 
.A1(n_12178),
.A2(n_12153),
.B1(n_12160),
.B2(n_12088),
.Y(n_12321)
);

OAI21xp5_ASAP7_75t_L g12322 ( 
.A1(n_12036),
.A2(n_1792),
.B(n_1793),
.Y(n_12322)
);

INVx3_ASAP7_75t_L g12323 ( 
.A(n_11961),
.Y(n_12323)
);

INVx1_ASAP7_75t_L g12324 ( 
.A(n_11871),
.Y(n_12324)
);

INVxp67_ASAP7_75t_L g12325 ( 
.A(n_12038),
.Y(n_12325)
);

OR2x6_ASAP7_75t_L g12326 ( 
.A(n_12040),
.B(n_1792),
.Y(n_12326)
);

OAI21xp5_ASAP7_75t_L g12327 ( 
.A1(n_12105),
.A2(n_1794),
.B(n_1795),
.Y(n_12327)
);

AND2x2_ASAP7_75t_SL g12328 ( 
.A(n_12141),
.B(n_1794),
.Y(n_12328)
);

INVx1_ASAP7_75t_L g12329 ( 
.A(n_11873),
.Y(n_12329)
);

OAI22xp5_ASAP7_75t_L g12330 ( 
.A1(n_12165),
.A2(n_1797),
.B1(n_1795),
.B2(n_1796),
.Y(n_12330)
);

AOI21xp5_ASAP7_75t_L g12331 ( 
.A1(n_11865),
.A2(n_12140),
.B(n_11896),
.Y(n_12331)
);

CKINVDCx5p33_ASAP7_75t_R g12332 ( 
.A(n_11988),
.Y(n_12332)
);

OAI21xp33_ASAP7_75t_SL g12333 ( 
.A1(n_11940),
.A2(n_1797),
.B(n_1798),
.Y(n_12333)
);

O2A1O1Ixp33_ASAP7_75t_L g12334 ( 
.A1(n_12102),
.A2(n_1800),
.B(n_1798),
.C(n_1799),
.Y(n_12334)
);

AND2x2_ASAP7_75t_L g12335 ( 
.A(n_11968),
.B(n_12021),
.Y(n_12335)
);

OAI22xp5_ASAP7_75t_L g12336 ( 
.A1(n_12114),
.A2(n_1802),
.B1(n_1800),
.B2(n_1801),
.Y(n_12336)
);

OR2x6_ASAP7_75t_L g12337 ( 
.A(n_12040),
.B(n_1801),
.Y(n_12337)
);

AO21x2_ASAP7_75t_L g12338 ( 
.A1(n_11934),
.A2(n_1802),
.B(n_1803),
.Y(n_12338)
);

OA21x2_ASAP7_75t_L g12339 ( 
.A1(n_12035),
.A2(n_1803),
.B(n_1804),
.Y(n_12339)
);

INVx2_ASAP7_75t_L g12340 ( 
.A(n_12049),
.Y(n_12340)
);

AND2x2_ASAP7_75t_L g12341 ( 
.A(n_12022),
.B(n_1805),
.Y(n_12341)
);

AO32x2_ASAP7_75t_L g12342 ( 
.A1(n_12092),
.A2(n_1808),
.A3(n_1806),
.B1(n_1807),
.B2(n_1809),
.Y(n_12342)
);

AOI22xp5_ASAP7_75t_L g12343 ( 
.A1(n_12063),
.A2(n_1809),
.B1(n_1807),
.B2(n_1808),
.Y(n_12343)
);

NAND2xp5_ASAP7_75t_L g12344 ( 
.A(n_12136),
.B(n_1810),
.Y(n_12344)
);

INVx1_ASAP7_75t_L g12345 ( 
.A(n_11875),
.Y(n_12345)
);

INVx2_ASAP7_75t_L g12346 ( 
.A(n_12049),
.Y(n_12346)
);

O2A1O1Ixp33_ASAP7_75t_L g12347 ( 
.A1(n_12163),
.A2(n_1812),
.B(n_1810),
.C(n_1811),
.Y(n_12347)
);

AND2x2_ASAP7_75t_L g12348 ( 
.A(n_12085),
.B(n_1811),
.Y(n_12348)
);

OAI21xp5_ASAP7_75t_L g12349 ( 
.A1(n_12077),
.A2(n_1813),
.B(n_1814),
.Y(n_12349)
);

NAND4xp25_ASAP7_75t_L g12350 ( 
.A(n_12170),
.B(n_1816),
.C(n_1813),
.D(n_1815),
.Y(n_12350)
);

NAND2xp5_ASAP7_75t_L g12351 ( 
.A(n_12099),
.B(n_1815),
.Y(n_12351)
);

INVx1_ASAP7_75t_L g12352 ( 
.A(n_11877),
.Y(n_12352)
);

OR2x2_ASAP7_75t_L g12353 ( 
.A(n_11959),
.B(n_1817),
.Y(n_12353)
);

A2O1A1Ixp33_ASAP7_75t_L g12354 ( 
.A1(n_12139),
.A2(n_1819),
.B(n_1817),
.C(n_1818),
.Y(n_12354)
);

AND2x2_ASAP7_75t_L g12355 ( 
.A(n_12096),
.B(n_1818),
.Y(n_12355)
);

BUFx3_ASAP7_75t_L g12356 ( 
.A(n_11912),
.Y(n_12356)
);

NAND2xp5_ASAP7_75t_L g12357 ( 
.A(n_12031),
.B(n_1819),
.Y(n_12357)
);

AO32x2_ASAP7_75t_L g12358 ( 
.A1(n_11973),
.A2(n_1822),
.A3(n_1820),
.B1(n_1821),
.B2(n_1823),
.Y(n_12358)
);

A2O1A1Ixp33_ASAP7_75t_L g12359 ( 
.A1(n_12098),
.A2(n_12166),
.B(n_12181),
.C(n_12149),
.Y(n_12359)
);

OAI221xp5_ASAP7_75t_L g12360 ( 
.A1(n_12058),
.A2(n_1822),
.B1(n_1820),
.B2(n_1821),
.C(n_1823),
.Y(n_12360)
);

AND2x2_ASAP7_75t_L g12361 ( 
.A(n_12046),
.B(n_1824),
.Y(n_12361)
);

BUFx3_ASAP7_75t_L g12362 ( 
.A(n_11943),
.Y(n_12362)
);

OR2x2_ASAP7_75t_L g12363 ( 
.A(n_11937),
.B(n_12106),
.Y(n_12363)
);

AND2x2_ASAP7_75t_L g12364 ( 
.A(n_12023),
.B(n_1824),
.Y(n_12364)
);

NOR2x1_ASAP7_75t_SL g12365 ( 
.A(n_11885),
.B(n_1825),
.Y(n_12365)
);

AND2x2_ASAP7_75t_L g12366 ( 
.A(n_11881),
.B(n_1825),
.Y(n_12366)
);

AOI221xp5_ASAP7_75t_L g12367 ( 
.A1(n_12053),
.A2(n_1828),
.B1(n_1826),
.B2(n_1827),
.C(n_1829),
.Y(n_12367)
);

INVxp67_ASAP7_75t_L g12368 ( 
.A(n_12057),
.Y(n_12368)
);

OAI21xp5_ASAP7_75t_L g12369 ( 
.A1(n_12192),
.A2(n_1826),
.B(n_1827),
.Y(n_12369)
);

BUFx10_ASAP7_75t_L g12370 ( 
.A(n_12079),
.Y(n_12370)
);

AND2x4_ASAP7_75t_L g12371 ( 
.A(n_11923),
.B(n_11953),
.Y(n_12371)
);

A2O1A1Ixp33_ASAP7_75t_L g12372 ( 
.A1(n_12145),
.A2(n_1830),
.B(n_1828),
.C(n_1829),
.Y(n_12372)
);

HB1xp67_ASAP7_75t_L g12373 ( 
.A(n_11925),
.Y(n_12373)
);

AND2x2_ASAP7_75t_L g12374 ( 
.A(n_12027),
.B(n_1830),
.Y(n_12374)
);

A2O1A1Ixp33_ASAP7_75t_L g12375 ( 
.A1(n_12183),
.A2(n_1834),
.B(n_1831),
.C(n_1833),
.Y(n_12375)
);

AOI221xp5_ASAP7_75t_L g12376 ( 
.A1(n_11991),
.A2(n_1834),
.B1(n_1831),
.B2(n_1833),
.C(n_1835),
.Y(n_12376)
);

BUFx3_ASAP7_75t_L g12377 ( 
.A(n_11976),
.Y(n_12377)
);

AND2x6_ASAP7_75t_L g12378 ( 
.A(n_12037),
.B(n_1836),
.Y(n_12378)
);

INVx1_ASAP7_75t_L g12379 ( 
.A(n_11879),
.Y(n_12379)
);

OAI21xp5_ASAP7_75t_L g12380 ( 
.A1(n_11900),
.A2(n_1836),
.B(n_1837),
.Y(n_12380)
);

AO21x2_ASAP7_75t_L g12381 ( 
.A1(n_11995),
.A2(n_1837),
.B(n_1838),
.Y(n_12381)
);

AOI22xp33_ASAP7_75t_SL g12382 ( 
.A1(n_12175),
.A2(n_1840),
.B1(n_1838),
.B2(n_1839),
.Y(n_12382)
);

AND2x4_ASAP7_75t_L g12383 ( 
.A(n_11957),
.B(n_1839),
.Y(n_12383)
);

NAND2xp5_ASAP7_75t_L g12384 ( 
.A(n_12030),
.B(n_1840),
.Y(n_12384)
);

INVx1_ASAP7_75t_SL g12385 ( 
.A(n_12000),
.Y(n_12385)
);

A2O1A1Ixp33_ASAP7_75t_L g12386 ( 
.A1(n_12104),
.A2(n_1843),
.B(n_1841),
.C(n_1842),
.Y(n_12386)
);

AOI21xp5_ASAP7_75t_L g12387 ( 
.A1(n_12156),
.A2(n_1841),
.B(n_1843),
.Y(n_12387)
);

BUFx4f_ASAP7_75t_L g12388 ( 
.A(n_11976),
.Y(n_12388)
);

INVx3_ASAP7_75t_L g12389 ( 
.A(n_11984),
.Y(n_12389)
);

NAND4xp25_ASAP7_75t_L g12390 ( 
.A(n_12054),
.B(n_1846),
.C(n_1844),
.D(n_1845),
.Y(n_12390)
);

AND2x2_ASAP7_75t_L g12391 ( 
.A(n_12065),
.B(n_1845),
.Y(n_12391)
);

AND2x2_ASAP7_75t_L g12392 ( 
.A(n_12109),
.B(n_1847),
.Y(n_12392)
);

AND2x2_ASAP7_75t_L g12393 ( 
.A(n_12108),
.B(n_1847),
.Y(n_12393)
);

INVx1_ASAP7_75t_L g12394 ( 
.A(n_11883),
.Y(n_12394)
);

OAI22xp5_ASAP7_75t_L g12395 ( 
.A1(n_12167),
.A2(n_1850),
.B1(n_1848),
.B2(n_1849),
.Y(n_12395)
);

NOR2x1_ASAP7_75t_L g12396 ( 
.A(n_12003),
.B(n_1848),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_11895),
.Y(n_12397)
);

AND2x4_ASAP7_75t_L g12398 ( 
.A(n_12073),
.B(n_1849),
.Y(n_12398)
);

AND2x2_ASAP7_75t_L g12399 ( 
.A(n_11982),
.B(n_1851),
.Y(n_12399)
);

INVx1_ASAP7_75t_L g12400 ( 
.A(n_11898),
.Y(n_12400)
);

AND2x4_ASAP7_75t_SL g12401 ( 
.A(n_12073),
.B(n_1851),
.Y(n_12401)
);

AND2x2_ASAP7_75t_L g12402 ( 
.A(n_12084),
.B(n_1852),
.Y(n_12402)
);

OAI21xp5_ASAP7_75t_L g12403 ( 
.A1(n_12168),
.A2(n_1852),
.B(n_1853),
.Y(n_12403)
);

INVx1_ASAP7_75t_L g12404 ( 
.A(n_11903),
.Y(n_12404)
);

AOI22xp5_ASAP7_75t_L g12405 ( 
.A1(n_12174),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.Y(n_12405)
);

BUFx3_ASAP7_75t_L g12406 ( 
.A(n_12071),
.Y(n_12406)
);

INVx1_ASAP7_75t_L g12407 ( 
.A(n_11906),
.Y(n_12407)
);

AO21x1_ASAP7_75t_L g12408 ( 
.A1(n_11945),
.A2(n_1855),
.B(n_1856),
.Y(n_12408)
);

NOR2x1_ASAP7_75t_SL g12409 ( 
.A(n_11971),
.B(n_1857),
.Y(n_12409)
);

INVx1_ASAP7_75t_L g12410 ( 
.A(n_11908),
.Y(n_12410)
);

A2O1A1Ixp33_ASAP7_75t_L g12411 ( 
.A1(n_12132),
.A2(n_1861),
.B(n_1859),
.C(n_1860),
.Y(n_12411)
);

AND2x4_ASAP7_75t_L g12412 ( 
.A(n_11870),
.B(n_1859),
.Y(n_12412)
);

AND2x2_ASAP7_75t_L g12413 ( 
.A(n_12089),
.B(n_1860),
.Y(n_12413)
);

HB1xp67_ASAP7_75t_L g12414 ( 
.A(n_12194),
.Y(n_12414)
);

NOR2xp33_ASAP7_75t_L g12415 ( 
.A(n_12070),
.B(n_1861),
.Y(n_12415)
);

AND2x2_ASAP7_75t_L g12416 ( 
.A(n_12171),
.B(n_1862),
.Y(n_12416)
);

AND2x2_ASAP7_75t_L g12417 ( 
.A(n_12074),
.B(n_1862),
.Y(n_12417)
);

NAND2xp5_ASAP7_75t_L g12418 ( 
.A(n_12010),
.B(n_1863),
.Y(n_12418)
);

OR2x2_ASAP7_75t_L g12419 ( 
.A(n_12001),
.B(n_1863),
.Y(n_12419)
);

AND2x2_ASAP7_75t_L g12420 ( 
.A(n_12110),
.B(n_1864),
.Y(n_12420)
);

NOR2x1_ASAP7_75t_L g12421 ( 
.A(n_11977),
.B(n_1864),
.Y(n_12421)
);

NAND3xp33_ASAP7_75t_L g12422 ( 
.A(n_11954),
.B(n_1865),
.C(n_1866),
.Y(n_12422)
);

NAND2xp5_ASAP7_75t_SL g12423 ( 
.A(n_12172),
.B(n_1865),
.Y(n_12423)
);

OAI22xp5_ASAP7_75t_L g12424 ( 
.A1(n_12176),
.A2(n_1869),
.B1(n_1867),
.B2(n_1868),
.Y(n_12424)
);

OAI21xp5_ASAP7_75t_L g12425 ( 
.A1(n_12068),
.A2(n_1867),
.B(n_1868),
.Y(n_12425)
);

O2A1O1Ixp33_ASAP7_75t_SL g12426 ( 
.A1(n_12100),
.A2(n_1871),
.B(n_1869),
.C(n_1870),
.Y(n_12426)
);

NAND2xp5_ASAP7_75t_L g12427 ( 
.A(n_12062),
.B(n_1870),
.Y(n_12427)
);

AOI22xp5_ASAP7_75t_L g12428 ( 
.A1(n_12172),
.A2(n_1873),
.B1(n_1871),
.B2(n_1872),
.Y(n_12428)
);

AOI22xp5_ASAP7_75t_L g12429 ( 
.A1(n_12155),
.A2(n_1875),
.B1(n_1872),
.B2(n_1874),
.Y(n_12429)
);

NAND2xp5_ASAP7_75t_L g12430 ( 
.A(n_12002),
.B(n_1874),
.Y(n_12430)
);

INVx3_ASAP7_75t_L g12431 ( 
.A(n_12083),
.Y(n_12431)
);

NAND2xp5_ASAP7_75t_L g12432 ( 
.A(n_12020),
.B(n_1875),
.Y(n_12432)
);

HB1xp67_ASAP7_75t_L g12433 ( 
.A(n_12195),
.Y(n_12433)
);

OR2x2_ASAP7_75t_L g12434 ( 
.A(n_12024),
.B(n_1876),
.Y(n_12434)
);

AND2x2_ASAP7_75t_L g12435 ( 
.A(n_12081),
.B(n_1876),
.Y(n_12435)
);

OR2x2_ASAP7_75t_L g12436 ( 
.A(n_12026),
.B(n_1877),
.Y(n_12436)
);

INVx1_ASAP7_75t_L g12437 ( 
.A(n_12196),
.Y(n_12437)
);

AO32x2_ASAP7_75t_L g12438 ( 
.A1(n_12086),
.A2(n_1879),
.A3(n_1877),
.B1(n_1878),
.B2(n_1880),
.Y(n_12438)
);

INVx2_ASAP7_75t_L g12439 ( 
.A(n_11975),
.Y(n_12439)
);

AND2x2_ASAP7_75t_L g12440 ( 
.A(n_12082),
.B(n_1878),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_12019),
.Y(n_12441)
);

INVx1_ASAP7_75t_L g12442 ( 
.A(n_11918),
.Y(n_12442)
);

OR2x2_ASAP7_75t_L g12443 ( 
.A(n_12029),
.B(n_1880),
.Y(n_12443)
);

AO32x2_ASAP7_75t_L g12444 ( 
.A1(n_11878),
.A2(n_1883),
.A3(n_1881),
.B1(n_1882),
.B2(n_1884),
.Y(n_12444)
);

AOI22xp5_ASAP7_75t_L g12445 ( 
.A1(n_12188),
.A2(n_1885),
.B1(n_1881),
.B2(n_1884),
.Y(n_12445)
);

AOI22xp33_ASAP7_75t_L g12446 ( 
.A1(n_12017),
.A2(n_1888),
.B1(n_1885),
.B2(n_1887),
.Y(n_12446)
);

INVx1_ASAP7_75t_L g12447 ( 
.A(n_11924),
.Y(n_12447)
);

AND2x2_ASAP7_75t_L g12448 ( 
.A(n_12056),
.B(n_11866),
.Y(n_12448)
);

A2O1A1Ixp33_ASAP7_75t_L g12449 ( 
.A1(n_12128),
.A2(n_1890),
.B(n_1887),
.C(n_1888),
.Y(n_12449)
);

OR2x2_ASAP7_75t_L g12450 ( 
.A(n_12011),
.B(n_1890),
.Y(n_12450)
);

NAND2x1_ASAP7_75t_L g12451 ( 
.A(n_12221),
.B(n_11966),
.Y(n_12451)
);

INVx5_ASAP7_75t_L g12452 ( 
.A(n_12204),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_12247),
.Y(n_12453)
);

INVx1_ASAP7_75t_L g12454 ( 
.A(n_12258),
.Y(n_12454)
);

HB1xp67_ASAP7_75t_L g12455 ( 
.A(n_12241),
.Y(n_12455)
);

AND2x2_ASAP7_75t_L g12456 ( 
.A(n_12226),
.B(n_12076),
.Y(n_12456)
);

AND2x2_ASAP7_75t_L g12457 ( 
.A(n_12212),
.B(n_11933),
.Y(n_12457)
);

OR2x2_ASAP7_75t_L g12458 ( 
.A(n_12227),
.B(n_11935),
.Y(n_12458)
);

INVx2_ASAP7_75t_L g12459 ( 
.A(n_12212),
.Y(n_12459)
);

INVx1_ASAP7_75t_L g12460 ( 
.A(n_12240),
.Y(n_12460)
);

BUFx3_ASAP7_75t_L g12461 ( 
.A(n_12204),
.Y(n_12461)
);

INVx1_ASAP7_75t_L g12462 ( 
.A(n_12312),
.Y(n_12462)
);

HB1xp67_ASAP7_75t_L g12463 ( 
.A(n_12267),
.Y(n_12463)
);

INVx1_ASAP7_75t_L g12464 ( 
.A(n_12414),
.Y(n_12464)
);

OAI31xp33_ASAP7_75t_SL g12465 ( 
.A1(n_12209),
.A2(n_12248),
.A3(n_12249),
.B(n_12396),
.Y(n_12465)
);

INVx2_ASAP7_75t_SL g12466 ( 
.A(n_12388),
.Y(n_12466)
);

HB1xp67_ASAP7_75t_L g12467 ( 
.A(n_12275),
.Y(n_12467)
);

OR2x2_ASAP7_75t_L g12468 ( 
.A(n_12315),
.B(n_12006),
.Y(n_12468)
);

HB1xp67_ASAP7_75t_L g12469 ( 
.A(n_12253),
.Y(n_12469)
);

INVx1_ASAP7_75t_L g12470 ( 
.A(n_12433),
.Y(n_12470)
);

INVx2_ASAP7_75t_L g12471 ( 
.A(n_12370),
.Y(n_12471)
);

INVx1_ASAP7_75t_L g12472 ( 
.A(n_12233),
.Y(n_12472)
);

INVxp67_ASAP7_75t_L g12473 ( 
.A(n_12365),
.Y(n_12473)
);

INVx2_ASAP7_75t_L g12474 ( 
.A(n_12264),
.Y(n_12474)
);

INVx2_ASAP7_75t_L g12475 ( 
.A(n_12264),
.Y(n_12475)
);

INVx2_ASAP7_75t_L g12476 ( 
.A(n_12406),
.Y(n_12476)
);

INVx2_ASAP7_75t_SL g12477 ( 
.A(n_12377),
.Y(n_12477)
);

INVx2_ASAP7_75t_L g12478 ( 
.A(n_12207),
.Y(n_12478)
);

INVx3_ASAP7_75t_L g12479 ( 
.A(n_12362),
.Y(n_12479)
);

INVx3_ASAP7_75t_R g12480 ( 
.A(n_12292),
.Y(n_12480)
);

INVx1_ASAP7_75t_L g12481 ( 
.A(n_12245),
.Y(n_12481)
);

AND2x2_ASAP7_75t_L g12482 ( 
.A(n_12276),
.B(n_11899),
.Y(n_12482)
);

BUFx6f_ASAP7_75t_L g12483 ( 
.A(n_12199),
.Y(n_12483)
);

INVx2_ASAP7_75t_L g12484 ( 
.A(n_12356),
.Y(n_12484)
);

INVx3_ASAP7_75t_L g12485 ( 
.A(n_12371),
.Y(n_12485)
);

OR2x2_ASAP7_75t_L g12486 ( 
.A(n_12297),
.B(n_12009),
.Y(n_12486)
);

AOI21xp5_ASAP7_75t_L g12487 ( 
.A1(n_12359),
.A2(n_11972),
.B(n_11970),
.Y(n_12487)
);

INVxp67_ASAP7_75t_L g12488 ( 
.A(n_12284),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_12206),
.Y(n_12489)
);

INVx1_ASAP7_75t_L g12490 ( 
.A(n_12216),
.Y(n_12490)
);

AND2x2_ASAP7_75t_L g12491 ( 
.A(n_12323),
.B(n_11874),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_12225),
.Y(n_12492)
);

INVx2_ASAP7_75t_L g12493 ( 
.A(n_12389),
.Y(n_12493)
);

HB1xp67_ASAP7_75t_L g12494 ( 
.A(n_12373),
.Y(n_12494)
);

NAND2xp5_ASAP7_75t_L g12495 ( 
.A(n_12328),
.B(n_12005),
.Y(n_12495)
);

INVx3_ASAP7_75t_L g12496 ( 
.A(n_12431),
.Y(n_12496)
);

INVx1_ASAP7_75t_L g12497 ( 
.A(n_12291),
.Y(n_12497)
);

NAND2xp5_ASAP7_75t_L g12498 ( 
.A(n_12385),
.B(n_12127),
.Y(n_12498)
);

NOR2xp33_ASAP7_75t_L g12499 ( 
.A(n_12325),
.B(n_12032),
.Y(n_12499)
);

INVx1_ASAP7_75t_L g12500 ( 
.A(n_12335),
.Y(n_12500)
);

BUFx3_ASAP7_75t_L g12501 ( 
.A(n_12378),
.Y(n_12501)
);

NOR2xp67_ASAP7_75t_L g12502 ( 
.A(n_12333),
.B(n_11967),
.Y(n_12502)
);

INVx2_ASAP7_75t_SL g12503 ( 
.A(n_12401),
.Y(n_12503)
);

INVx3_ASAP7_75t_L g12504 ( 
.A(n_12298),
.Y(n_12504)
);

HB1xp67_ASAP7_75t_L g12505 ( 
.A(n_12215),
.Y(n_12505)
);

AND2x4_ASAP7_75t_L g12506 ( 
.A(n_12260),
.B(n_11919),
.Y(n_12506)
);

OR2x2_ASAP7_75t_L g12507 ( 
.A(n_12363),
.B(n_11944),
.Y(n_12507)
);

INVx5_ASAP7_75t_L g12508 ( 
.A(n_12326),
.Y(n_12508)
);

INVx1_ASAP7_75t_L g12509 ( 
.A(n_12251),
.Y(n_12509)
);

INVx2_ASAP7_75t_L g12510 ( 
.A(n_12266),
.Y(n_12510)
);

INVx1_ASAP7_75t_L g12511 ( 
.A(n_12281),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_12244),
.Y(n_12512)
);

INVx1_ASAP7_75t_L g12513 ( 
.A(n_12441),
.Y(n_12513)
);

INVx1_ASAP7_75t_L g12514 ( 
.A(n_12314),
.Y(n_12514)
);

INVx1_ASAP7_75t_L g12515 ( 
.A(n_12341),
.Y(n_12515)
);

AND2x2_ASAP7_75t_L g12516 ( 
.A(n_12203),
.B(n_12103),
.Y(n_12516)
);

AND2x4_ASAP7_75t_L g12517 ( 
.A(n_12210),
.B(n_11948),
.Y(n_12517)
);

INVx1_ASAP7_75t_L g12518 ( 
.A(n_12361),
.Y(n_12518)
);

INVx1_ASAP7_75t_L g12519 ( 
.A(n_12374),
.Y(n_12519)
);

INVx1_ASAP7_75t_L g12520 ( 
.A(n_12305),
.Y(n_12520)
);

AND2x2_ASAP7_75t_L g12521 ( 
.A(n_12237),
.B(n_12118),
.Y(n_12521)
);

BUFx2_ASAP7_75t_L g12522 ( 
.A(n_12326),
.Y(n_12522)
);

INVx1_ASAP7_75t_L g12523 ( 
.A(n_12353),
.Y(n_12523)
);

AND2x2_ASAP7_75t_L g12524 ( 
.A(n_12340),
.B(n_12124),
.Y(n_12524)
);

INVx2_ASAP7_75t_L g12525 ( 
.A(n_12290),
.Y(n_12525)
);

HB1xp67_ASAP7_75t_L g12526 ( 
.A(n_12339),
.Y(n_12526)
);

INVxp67_ASAP7_75t_SL g12527 ( 
.A(n_12409),
.Y(n_12527)
);

INVx1_ASAP7_75t_L g12528 ( 
.A(n_12402),
.Y(n_12528)
);

INVx2_ASAP7_75t_L g12529 ( 
.A(n_12346),
.Y(n_12529)
);

INVxp67_ASAP7_75t_L g12530 ( 
.A(n_12421),
.Y(n_12530)
);

INVx2_ASAP7_75t_L g12531 ( 
.A(n_12222),
.Y(n_12531)
);

AND2x2_ASAP7_75t_L g12532 ( 
.A(n_12200),
.B(n_11932),
.Y(n_12532)
);

HB1xp67_ASAP7_75t_L g12533 ( 
.A(n_12337),
.Y(n_12533)
);

INVxp67_ASAP7_75t_L g12534 ( 
.A(n_12265),
.Y(n_12534)
);

INVx1_ASAP7_75t_L g12535 ( 
.A(n_12211),
.Y(n_12535)
);

AND2x2_ASAP7_75t_L g12536 ( 
.A(n_12448),
.B(n_12093),
.Y(n_12536)
);

AND2x2_ASAP7_75t_L g12537 ( 
.A(n_12285),
.B(n_11979),
.Y(n_12537)
);

AND2x2_ASAP7_75t_L g12538 ( 
.A(n_12368),
.B(n_11981),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_12224),
.Y(n_12539)
);

INVx3_ASAP7_75t_L g12540 ( 
.A(n_12311),
.Y(n_12540)
);

OR2x2_ASAP7_75t_L g12541 ( 
.A(n_12321),
.B(n_11974),
.Y(n_12541)
);

INVx1_ASAP7_75t_L g12542 ( 
.A(n_12364),
.Y(n_12542)
);

INVx2_ASAP7_75t_L g12543 ( 
.A(n_12337),
.Y(n_12543)
);

NAND2xp5_ASAP7_75t_L g12544 ( 
.A(n_12302),
.B(n_12135),
.Y(n_12544)
);

INVx2_ASAP7_75t_L g12545 ( 
.A(n_12296),
.Y(n_12545)
);

AOI21xp33_ASAP7_75t_L g12546 ( 
.A1(n_12198),
.A2(n_11983),
.B(n_11985),
.Y(n_12546)
);

INVx1_ASAP7_75t_L g12547 ( 
.A(n_12289),
.Y(n_12547)
);

INVx3_ASAP7_75t_SL g12548 ( 
.A(n_12332),
.Y(n_12548)
);

OR2x2_ASAP7_75t_L g12549 ( 
.A(n_12255),
.B(n_11996),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_12416),
.B(n_11986),
.Y(n_12550)
);

INVx2_ASAP7_75t_L g12551 ( 
.A(n_12296),
.Y(n_12551)
);

AND2x2_ASAP7_75t_L g12552 ( 
.A(n_12205),
.B(n_11951),
.Y(n_12552)
);

INVxp67_ASAP7_75t_SL g12553 ( 
.A(n_12408),
.Y(n_12553)
);

NAND2xp5_ASAP7_75t_L g12554 ( 
.A(n_12263),
.B(n_12119),
.Y(n_12554)
);

INVx1_ASAP7_75t_L g12555 ( 
.A(n_12295),
.Y(n_12555)
);

BUFx3_ASAP7_75t_L g12556 ( 
.A(n_12378),
.Y(n_12556)
);

INVx1_ASAP7_75t_L g12557 ( 
.A(n_12324),
.Y(n_12557)
);

AND2x2_ASAP7_75t_L g12558 ( 
.A(n_12271),
.B(n_11978),
.Y(n_12558)
);

NAND2xp5_ASAP7_75t_L g12559 ( 
.A(n_12387),
.B(n_12101),
.Y(n_12559)
);

AND2x2_ASAP7_75t_L g12560 ( 
.A(n_12399),
.B(n_12044),
.Y(n_12560)
);

INVx4_ASAP7_75t_L g12561 ( 
.A(n_12310),
.Y(n_12561)
);

INVx1_ASAP7_75t_L g12562 ( 
.A(n_12329),
.Y(n_12562)
);

AND2x2_ASAP7_75t_L g12563 ( 
.A(n_12232),
.B(n_12047),
.Y(n_12563)
);

AND2x2_ASAP7_75t_L g12564 ( 
.A(n_12231),
.B(n_12055),
.Y(n_12564)
);

AND2x2_ASAP7_75t_L g12565 ( 
.A(n_12391),
.B(n_12064),
.Y(n_12565)
);

AND2x4_ASAP7_75t_L g12566 ( 
.A(n_12252),
.B(n_12087),
.Y(n_12566)
);

OR2x2_ASAP7_75t_L g12567 ( 
.A(n_12283),
.B(n_11998),
.Y(n_12567)
);

OR2x2_ASAP7_75t_L g12568 ( 
.A(n_12293),
.B(n_12004),
.Y(n_12568)
);

BUFx2_ASAP7_75t_L g12569 ( 
.A(n_12378),
.Y(n_12569)
);

INVx3_ASAP7_75t_SL g12570 ( 
.A(n_12304),
.Y(n_12570)
);

INVx2_ASAP7_75t_L g12571 ( 
.A(n_12213),
.Y(n_12571)
);

INVx1_ASAP7_75t_L g12572 ( 
.A(n_12345),
.Y(n_12572)
);

INVx2_ASAP7_75t_L g12573 ( 
.A(n_12300),
.Y(n_12573)
);

BUFx2_ASAP7_75t_L g12574 ( 
.A(n_12358),
.Y(n_12574)
);

INVx2_ASAP7_75t_L g12575 ( 
.A(n_12366),
.Y(n_12575)
);

INVx1_ASAP7_75t_L g12576 ( 
.A(n_12352),
.Y(n_12576)
);

NAND2xp5_ASAP7_75t_L g12577 ( 
.A(n_12308),
.B(n_11947),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_12379),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_12394),
.Y(n_12579)
);

INVxp33_ASAP7_75t_L g12580 ( 
.A(n_12423),
.Y(n_12580)
);

AND2x2_ASAP7_75t_L g12581 ( 
.A(n_12270),
.B(n_12025),
.Y(n_12581)
);

OR2x2_ASAP7_75t_L g12582 ( 
.A(n_12306),
.B(n_12007),
.Y(n_12582)
);

NAND2x1p5_ASAP7_75t_L g12583 ( 
.A(n_12230),
.B(n_12075),
.Y(n_12583)
);

OAI211xp5_ASAP7_75t_L g12584 ( 
.A1(n_12429),
.A2(n_12151),
.B(n_12185),
.C(n_12158),
.Y(n_12584)
);

NAND2xp5_ASAP7_75t_SL g12585 ( 
.A(n_12380),
.B(n_12094),
.Y(n_12585)
);

AOI22xp5_ASAP7_75t_L g12586 ( 
.A1(n_12282),
.A2(n_12164),
.B1(n_12133),
.B2(n_12043),
.Y(n_12586)
);

INVx3_ASAP7_75t_L g12587 ( 
.A(n_12398),
.Y(n_12587)
);

INVx2_ASAP7_75t_L g12588 ( 
.A(n_12288),
.Y(n_12588)
);

BUFx4f_ASAP7_75t_L g12589 ( 
.A(n_12383),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_12397),
.Y(n_12590)
);

AND2x4_ASAP7_75t_L g12591 ( 
.A(n_12234),
.B(n_12033),
.Y(n_12591)
);

INVx1_ASAP7_75t_L g12592 ( 
.A(n_12400),
.Y(n_12592)
);

INVx2_ASAP7_75t_L g12593 ( 
.A(n_12303),
.Y(n_12593)
);

INVx1_ASAP7_75t_L g12594 ( 
.A(n_12404),
.Y(n_12594)
);

OR2x2_ASAP7_75t_L g12595 ( 
.A(n_12318),
.B(n_11964),
.Y(n_12595)
);

INVx3_ASAP7_75t_L g12596 ( 
.A(n_12412),
.Y(n_12596)
);

INVx1_ASAP7_75t_L g12597 ( 
.A(n_12407),
.Y(n_12597)
);

INVx1_ASAP7_75t_L g12598 ( 
.A(n_12450),
.Y(n_12598)
);

INVx2_ASAP7_75t_L g12599 ( 
.A(n_12278),
.Y(n_12599)
);

BUFx3_ASAP7_75t_L g12600 ( 
.A(n_12228),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_12413),
.Y(n_12601)
);

INVx1_ASAP7_75t_L g12602 ( 
.A(n_12435),
.Y(n_12602)
);

HB1xp67_ASAP7_75t_L g12603 ( 
.A(n_12313),
.Y(n_12603)
);

AND2x2_ASAP7_75t_L g12604 ( 
.A(n_12235),
.B(n_12048),
.Y(n_12604)
);

OR2x2_ASAP7_75t_L g12605 ( 
.A(n_12331),
.B(n_12080),
.Y(n_12605)
);

OAI22xp5_ASAP7_75t_L g12606 ( 
.A1(n_12405),
.A2(n_11942),
.B1(n_12113),
.B2(n_12154),
.Y(n_12606)
);

BUFx2_ASAP7_75t_L g12607 ( 
.A(n_12358),
.Y(n_12607)
);

BUFx6f_ASAP7_75t_L g12608 ( 
.A(n_12272),
.Y(n_12608)
);

AND2x2_ASAP7_75t_L g12609 ( 
.A(n_12393),
.B(n_11927),
.Y(n_12609)
);

AND2x2_ASAP7_75t_L g12610 ( 
.A(n_12274),
.B(n_11992),
.Y(n_12610)
);

AOI22xp5_ASAP7_75t_L g12611 ( 
.A1(n_12280),
.A2(n_12116),
.B1(n_12126),
.B2(n_12162),
.Y(n_12611)
);

INVx1_ASAP7_75t_L g12612 ( 
.A(n_12440),
.Y(n_12612)
);

INVx2_ASAP7_75t_L g12613 ( 
.A(n_12348),
.Y(n_12613)
);

AOI22xp33_ASAP7_75t_L g12614 ( 
.A1(n_12223),
.A2(n_11952),
.B1(n_12039),
.B2(n_1893),
.Y(n_12614)
);

AND2x4_ASAP7_75t_L g12615 ( 
.A(n_12309),
.B(n_11952),
.Y(n_12615)
);

NAND2xp5_ASAP7_75t_L g12616 ( 
.A(n_12382),
.B(n_12386),
.Y(n_12616)
);

AND2x2_ASAP7_75t_L g12617 ( 
.A(n_12417),
.B(n_12039),
.Y(n_12617)
);

AOI22xp5_ASAP7_75t_L g12618 ( 
.A1(n_12242),
.A2(n_1893),
.B1(n_1891),
.B2(n_1892),
.Y(n_12618)
);

INVx1_ASAP7_75t_L g12619 ( 
.A(n_12410),
.Y(n_12619)
);

INVx2_ASAP7_75t_L g12620 ( 
.A(n_12355),
.Y(n_12620)
);

INVx4_ASAP7_75t_L g12621 ( 
.A(n_12392),
.Y(n_12621)
);

OR2x2_ASAP7_75t_L g12622 ( 
.A(n_12254),
.B(n_1892),
.Y(n_12622)
);

INVx2_ASAP7_75t_L g12623 ( 
.A(n_12338),
.Y(n_12623)
);

AND2x4_ASAP7_75t_SL g12624 ( 
.A(n_12229),
.B(n_1895),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12217),
.Y(n_12625)
);

INVx3_ASAP7_75t_L g12626 ( 
.A(n_12439),
.Y(n_12626)
);

AOI322xp5_ASAP7_75t_L g12627 ( 
.A1(n_12201),
.A2(n_1900),
.A3(n_1899),
.B1(n_1897),
.B2(n_1895),
.C1(n_1896),
.C2(n_1898),
.Y(n_12627)
);

OR2x2_ASAP7_75t_L g12628 ( 
.A(n_12437),
.B(n_1896),
.Y(n_12628)
);

INVx2_ASAP7_75t_L g12629 ( 
.A(n_12299),
.Y(n_12629)
);

INVx1_ASAP7_75t_L g12630 ( 
.A(n_12236),
.Y(n_12630)
);

INVx1_ASAP7_75t_L g12631 ( 
.A(n_12442),
.Y(n_12631)
);

AND2x4_ASAP7_75t_L g12632 ( 
.A(n_12420),
.B(n_1897),
.Y(n_12632)
);

NOR2xp67_ASAP7_75t_L g12633 ( 
.A(n_12218),
.B(n_1899),
.Y(n_12633)
);

INVx1_ASAP7_75t_L g12634 ( 
.A(n_12447),
.Y(n_12634)
);

INVx1_ASAP7_75t_L g12635 ( 
.A(n_12434),
.Y(n_12635)
);

HB1xp67_ASAP7_75t_L g12636 ( 
.A(n_12381),
.Y(n_12636)
);

AND2x4_ASAP7_75t_L g12637 ( 
.A(n_12219),
.B(n_1900),
.Y(n_12637)
);

AND2x2_ASAP7_75t_L g12638 ( 
.A(n_12369),
.B(n_1901),
.Y(n_12638)
);

INVx2_ASAP7_75t_L g12639 ( 
.A(n_12277),
.Y(n_12639)
);

INVx2_ASAP7_75t_L g12640 ( 
.A(n_12419),
.Y(n_12640)
);

INVxp67_ASAP7_75t_SL g12641 ( 
.A(n_12344),
.Y(n_12641)
);

HB1xp67_ASAP7_75t_L g12642 ( 
.A(n_12436),
.Y(n_12642)
);

HB1xp67_ASAP7_75t_L g12643 ( 
.A(n_12443),
.Y(n_12643)
);

BUFx2_ASAP7_75t_L g12644 ( 
.A(n_12342),
.Y(n_12644)
);

INVx1_ASAP7_75t_L g12645 ( 
.A(n_12357),
.Y(n_12645)
);

NAND2xp5_ASAP7_75t_L g12646 ( 
.A(n_12238),
.B(n_1901),
.Y(n_12646)
);

INVx2_ASAP7_75t_L g12647 ( 
.A(n_12307),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_12384),
.Y(n_12648)
);

INVx1_ASAP7_75t_L g12649 ( 
.A(n_12320),
.Y(n_12649)
);

INVx4_ASAP7_75t_L g12650 ( 
.A(n_12343),
.Y(n_12650)
);

NAND2xp5_ASAP7_75t_L g12651 ( 
.A(n_12208),
.B(n_12351),
.Y(n_12651)
);

NAND2xp5_ASAP7_75t_L g12652 ( 
.A(n_12250),
.B(n_1902),
.Y(n_12652)
);

AND2x2_ASAP7_75t_L g12653 ( 
.A(n_12461),
.B(n_12319),
.Y(n_12653)
);

NAND2xp5_ASAP7_75t_L g12654 ( 
.A(n_12644),
.B(n_12261),
.Y(n_12654)
);

NAND3xp33_ASAP7_75t_L g12655 ( 
.A(n_12553),
.B(n_12367),
.C(n_12214),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_12452),
.B(n_12259),
.Y(n_12656)
);

NOR3xp33_ASAP7_75t_L g12657 ( 
.A(n_12471),
.B(n_12334),
.C(n_12294),
.Y(n_12657)
);

AND2x2_ASAP7_75t_L g12658 ( 
.A(n_12452),
.B(n_12570),
.Y(n_12658)
);

AND2x2_ASAP7_75t_L g12659 ( 
.A(n_12466),
.B(n_12432),
.Y(n_12659)
);

OAI21xp5_ASAP7_75t_SL g12660 ( 
.A1(n_12465),
.A2(n_12322),
.B(n_12316),
.Y(n_12660)
);

INVx1_ASAP7_75t_L g12661 ( 
.A(n_12455),
.Y(n_12661)
);

OAI221xp5_ASAP7_75t_L g12662 ( 
.A1(n_12530),
.A2(n_12554),
.B1(n_12614),
.B2(n_12546),
.C(n_12487),
.Y(n_12662)
);

AND2x2_ASAP7_75t_L g12663 ( 
.A(n_12479),
.B(n_12415),
.Y(n_12663)
);

NAND2xp5_ASAP7_75t_L g12664 ( 
.A(n_12574),
.B(n_12430),
.Y(n_12664)
);

NAND2xp5_ASAP7_75t_SL g12665 ( 
.A(n_12508),
.B(n_12246),
.Y(n_12665)
);

AND2x2_ASAP7_75t_SL g12666 ( 
.A(n_12589),
.B(n_12427),
.Y(n_12666)
);

NAND3xp33_ASAP7_75t_L g12667 ( 
.A(n_12534),
.B(n_12422),
.C(n_12376),
.Y(n_12667)
);

NAND3xp33_ASAP7_75t_L g12668 ( 
.A(n_12526),
.B(n_12279),
.C(n_12445),
.Y(n_12668)
);

AOI22xp33_ASAP7_75t_L g12669 ( 
.A1(n_12650),
.A2(n_12607),
.B1(n_12485),
.B2(n_12476),
.Y(n_12669)
);

AND2x2_ASAP7_75t_L g12670 ( 
.A(n_12552),
.B(n_12418),
.Y(n_12670)
);

NAND4xp25_ASAP7_75t_L g12671 ( 
.A(n_12499),
.B(n_12350),
.C(n_12347),
.D(n_12317),
.Y(n_12671)
);

OR2x2_ASAP7_75t_L g12672 ( 
.A(n_12498),
.B(n_12531),
.Y(n_12672)
);

NAND2xp5_ASAP7_75t_L g12673 ( 
.A(n_12508),
.B(n_12202),
.Y(n_12673)
);

NAND2xp5_ASAP7_75t_L g12674 ( 
.A(n_12569),
.B(n_12522),
.Y(n_12674)
);

OAI221xp5_ASAP7_75t_L g12675 ( 
.A1(n_12611),
.A2(n_12586),
.B1(n_12584),
.B2(n_12488),
.C(n_12473),
.Y(n_12675)
);

NAND3xp33_ASAP7_75t_L g12676 ( 
.A(n_12603),
.B(n_12425),
.C(n_12354),
.Y(n_12676)
);

NAND2xp5_ASAP7_75t_L g12677 ( 
.A(n_12533),
.B(n_12372),
.Y(n_12677)
);

NAND4xp25_ASAP7_75t_L g12678 ( 
.A(n_12563),
.B(n_12403),
.C(n_12268),
.D(n_12390),
.Y(n_12678)
);

OA21x2_ASAP7_75t_L g12679 ( 
.A1(n_12460),
.A2(n_12462),
.B(n_12623),
.Y(n_12679)
);

NAND2xp5_ASAP7_75t_L g12680 ( 
.A(n_12469),
.B(n_12256),
.Y(n_12680)
);

NAND2xp5_ASAP7_75t_L g12681 ( 
.A(n_12527),
.B(n_12330),
.Y(n_12681)
);

AND2x2_ASAP7_75t_L g12682 ( 
.A(n_12456),
.B(n_12327),
.Y(n_12682)
);

OAI21xp5_ASAP7_75t_SL g12683 ( 
.A1(n_12616),
.A2(n_12428),
.B(n_12269),
.Y(n_12683)
);

NAND2xp5_ASAP7_75t_L g12684 ( 
.A(n_12558),
.B(n_12449),
.Y(n_12684)
);

AND2x2_ASAP7_75t_L g12685 ( 
.A(n_12560),
.B(n_12262),
.Y(n_12685)
);

AND2x2_ASAP7_75t_L g12686 ( 
.A(n_12482),
.B(n_12273),
.Y(n_12686)
);

AND2x2_ASAP7_75t_L g12687 ( 
.A(n_12565),
.B(n_12286),
.Y(n_12687)
);

NAND2xp5_ASAP7_75t_L g12688 ( 
.A(n_12502),
.B(n_12426),
.Y(n_12688)
);

NOR2xp33_ASAP7_75t_L g12689 ( 
.A(n_12548),
.B(n_12301),
.Y(n_12689)
);

AND2x2_ASAP7_75t_L g12690 ( 
.A(n_12496),
.B(n_12444),
.Y(n_12690)
);

OAI21xp5_ASAP7_75t_SL g12691 ( 
.A1(n_12618),
.A2(n_12287),
.B(n_12243),
.Y(n_12691)
);

NOR3xp33_ASAP7_75t_L g12692 ( 
.A(n_12478),
.B(n_12360),
.C(n_12424),
.Y(n_12692)
);

AND2x2_ASAP7_75t_L g12693 ( 
.A(n_12459),
.B(n_12543),
.Y(n_12693)
);

AOI22xp33_ASAP7_75t_L g12694 ( 
.A1(n_12493),
.A2(n_12349),
.B1(n_12336),
.B2(n_12395),
.Y(n_12694)
);

NAND2xp5_ASAP7_75t_L g12695 ( 
.A(n_12463),
.B(n_12220),
.Y(n_12695)
);

NAND2xp5_ASAP7_75t_L g12696 ( 
.A(n_12587),
.B(n_12545),
.Y(n_12696)
);

NAND2xp5_ASAP7_75t_L g12697 ( 
.A(n_12551),
.B(n_12375),
.Y(n_12697)
);

OAI22xp33_ASAP7_75t_SL g12698 ( 
.A1(n_12451),
.A2(n_12629),
.B1(n_12583),
.B2(n_12541),
.Y(n_12698)
);

NAND2xp5_ASAP7_75t_L g12699 ( 
.A(n_12591),
.B(n_12411),
.Y(n_12699)
);

OAI21xp5_ASAP7_75t_SL g12700 ( 
.A1(n_12580),
.A2(n_12446),
.B(n_12239),
.Y(n_12700)
);

AND2x2_ASAP7_75t_L g12701 ( 
.A(n_12564),
.B(n_12444),
.Y(n_12701)
);

NOR2xp33_ASAP7_75t_L g12702 ( 
.A(n_12561),
.B(n_12239),
.Y(n_12702)
);

NAND3xp33_ASAP7_75t_SL g12703 ( 
.A(n_12544),
.B(n_12257),
.C(n_12342),
.Y(n_12703)
);

AOI22xp33_ASAP7_75t_SL g12704 ( 
.A1(n_12636),
.A2(n_12438),
.B1(n_12257),
.B2(n_1904),
.Y(n_12704)
);

OA21x2_ASAP7_75t_L g12705 ( 
.A1(n_12494),
.A2(n_12438),
.B(n_1902),
.Y(n_12705)
);

NAND2xp5_ASAP7_75t_L g12706 ( 
.A(n_12566),
.B(n_1903),
.Y(n_12706)
);

NOR3xp33_ASAP7_75t_SL g12707 ( 
.A(n_12453),
.B(n_12454),
.C(n_12641),
.Y(n_12707)
);

AOI22xp33_ASAP7_75t_SL g12708 ( 
.A1(n_12606),
.A2(n_1906),
.B1(n_1904),
.B2(n_1905),
.Y(n_12708)
);

OA21x2_ASAP7_75t_L g12709 ( 
.A1(n_12577),
.A2(n_1905),
.B(n_1907),
.Y(n_12709)
);

AND2x2_ASAP7_75t_L g12710 ( 
.A(n_12491),
.B(n_12503),
.Y(n_12710)
);

NAND2xp5_ASAP7_75t_SL g12711 ( 
.A(n_12483),
.B(n_1908),
.Y(n_12711)
);

NAND2xp5_ASAP7_75t_L g12712 ( 
.A(n_12581),
.B(n_1909),
.Y(n_12712)
);

NAND2xp5_ASAP7_75t_L g12713 ( 
.A(n_12588),
.B(n_1909),
.Y(n_12713)
);

AND2x2_ASAP7_75t_L g12714 ( 
.A(n_12484),
.B(n_1911),
.Y(n_12714)
);

OAI21xp33_ASAP7_75t_L g12715 ( 
.A1(n_12477),
.A2(n_1911),
.B(n_1912),
.Y(n_12715)
);

AND2x2_ASAP7_75t_L g12716 ( 
.A(n_12536),
.B(n_1912),
.Y(n_12716)
);

OAI221xp5_ASAP7_75t_L g12717 ( 
.A1(n_12651),
.A2(n_1915),
.B1(n_1913),
.B2(n_1914),
.C(n_1916),
.Y(n_12717)
);

NOR2xp33_ASAP7_75t_L g12718 ( 
.A(n_12480),
.B(n_1913),
.Y(n_12718)
);

AND2x2_ASAP7_75t_L g12719 ( 
.A(n_12467),
.B(n_1914),
.Y(n_12719)
);

OAI221xp5_ASAP7_75t_L g12720 ( 
.A1(n_12585),
.A2(n_1918),
.B1(n_1916),
.B2(n_1917),
.C(n_1919),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_12501),
.B(n_1918),
.Y(n_12721)
);

NOR3xp33_ASAP7_75t_L g12722 ( 
.A(n_12509),
.B(n_1920),
.C(n_1921),
.Y(n_12722)
);

NAND2xp5_ASAP7_75t_L g12723 ( 
.A(n_12556),
.B(n_1920),
.Y(n_12723)
);

NAND2xp5_ASAP7_75t_SL g12724 ( 
.A(n_12483),
.B(n_1922),
.Y(n_12724)
);

AND2x2_ASAP7_75t_L g12725 ( 
.A(n_12504),
.B(n_1922),
.Y(n_12725)
);

NAND4xp25_ASAP7_75t_L g12726 ( 
.A(n_12500),
.B(n_1925),
.C(n_1923),
.D(n_1924),
.Y(n_12726)
);

OAI221xp5_ASAP7_75t_L g12727 ( 
.A1(n_12559),
.A2(n_1927),
.B1(n_1924),
.B2(n_1926),
.C(n_1928),
.Y(n_12727)
);

NAND2xp5_ASAP7_75t_L g12728 ( 
.A(n_12505),
.B(n_1929),
.Y(n_12728)
);

NOR3xp33_ASAP7_75t_L g12729 ( 
.A(n_12640),
.B(n_1929),
.C(n_1930),
.Y(n_12729)
);

AND2x2_ASAP7_75t_L g12730 ( 
.A(n_12540),
.B(n_1930),
.Y(n_12730)
);

AND2x2_ASAP7_75t_L g12731 ( 
.A(n_12521),
.B(n_1933),
.Y(n_12731)
);

OAI21xp5_ASAP7_75t_L g12732 ( 
.A1(n_12652),
.A2(n_1933),
.B(n_1934),
.Y(n_12732)
);

AOI221xp5_ASAP7_75t_L g12733 ( 
.A1(n_12464),
.A2(n_1937),
.B1(n_1935),
.B2(n_1936),
.C(n_1938),
.Y(n_12733)
);

NAND2xp5_ASAP7_75t_L g12734 ( 
.A(n_12596),
.B(n_1935),
.Y(n_12734)
);

OAI221xp5_ASAP7_75t_SL g12735 ( 
.A1(n_12605),
.A2(n_1938),
.B1(n_1936),
.B2(n_1937),
.C(n_1939),
.Y(n_12735)
);

NAND3xp33_ASAP7_75t_SL g12736 ( 
.A(n_12495),
.B(n_1939),
.C(n_1940),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_12633),
.B(n_1940),
.Y(n_12737)
);

NAND3xp33_ASAP7_75t_L g12738 ( 
.A(n_12470),
.B(n_1941),
.C(n_1942),
.Y(n_12738)
);

NAND2xp5_ASAP7_75t_L g12739 ( 
.A(n_12604),
.B(n_1941),
.Y(n_12739)
);

OAI21xp33_ASAP7_75t_L g12740 ( 
.A1(n_12457),
.A2(n_12510),
.B(n_12529),
.Y(n_12740)
);

OAI22xp5_ASAP7_75t_L g12741 ( 
.A1(n_12637),
.A2(n_1944),
.B1(n_1942),
.B2(n_1943),
.Y(n_12741)
);

OAI221xp5_ASAP7_75t_SL g12742 ( 
.A1(n_12627),
.A2(n_1946),
.B1(n_1944),
.B2(n_1945),
.C(n_1947),
.Y(n_12742)
);

NAND3xp33_ASAP7_75t_L g12743 ( 
.A(n_12571),
.B(n_1946),
.C(n_1947),
.Y(n_12743)
);

AND2x2_ASAP7_75t_L g12744 ( 
.A(n_12474),
.B(n_1948),
.Y(n_12744)
);

NAND2xp5_ASAP7_75t_SL g12745 ( 
.A(n_12608),
.B(n_1948),
.Y(n_12745)
);

NAND3xp33_ASAP7_75t_L g12746 ( 
.A(n_12642),
.B(n_1950),
.C(n_1951),
.Y(n_12746)
);

AND2x2_ASAP7_75t_L g12747 ( 
.A(n_12475),
.B(n_1950),
.Y(n_12747)
);

AOI22xp33_ASAP7_75t_L g12748 ( 
.A1(n_12539),
.A2(n_1954),
.B1(n_1951),
.B2(n_1952),
.Y(n_12748)
);

AND2x2_ASAP7_75t_L g12749 ( 
.A(n_12516),
.B(n_1955),
.Y(n_12749)
);

NAND2xp5_ASAP7_75t_L g12750 ( 
.A(n_12506),
.B(n_1955),
.Y(n_12750)
);

AND2x2_ASAP7_75t_L g12751 ( 
.A(n_12532),
.B(n_1956),
.Y(n_12751)
);

AND2x2_ASAP7_75t_L g12752 ( 
.A(n_12524),
.B(n_1956),
.Y(n_12752)
);

NAND3xp33_ASAP7_75t_L g12753 ( 
.A(n_12643),
.B(n_1957),
.C(n_1958),
.Y(n_12753)
);

OAI22xp5_ASAP7_75t_L g12754 ( 
.A1(n_12646),
.A2(n_1960),
.B1(n_1957),
.B2(n_1959),
.Y(n_12754)
);

NAND3xp33_ASAP7_75t_L g12755 ( 
.A(n_12458),
.B(n_1959),
.C(n_1960),
.Y(n_12755)
);

NAND3xp33_ASAP7_75t_L g12756 ( 
.A(n_12621),
.B(n_1961),
.C(n_1962),
.Y(n_12756)
);

AOI22xp5_ASAP7_75t_L g12757 ( 
.A1(n_12517),
.A2(n_1965),
.B1(n_1963),
.B2(n_1964),
.Y(n_12757)
);

AND2x2_ASAP7_75t_L g12758 ( 
.A(n_12600),
.B(n_1964),
.Y(n_12758)
);

AOI221xp5_ASAP7_75t_L g12759 ( 
.A1(n_12472),
.A2(n_1967),
.B1(n_1965),
.B2(n_1966),
.C(n_1968),
.Y(n_12759)
);

AND2x2_ASAP7_75t_L g12760 ( 
.A(n_12537),
.B(n_1966),
.Y(n_12760)
);

AOI22xp33_ASAP7_75t_L g12761 ( 
.A1(n_12608),
.A2(n_1970),
.B1(n_1967),
.B2(n_1969),
.Y(n_12761)
);

AND2x2_ASAP7_75t_L g12762 ( 
.A(n_12610),
.B(n_1970),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_12550),
.B(n_12593),
.Y(n_12763)
);

AND2x2_ASAP7_75t_L g12764 ( 
.A(n_12599),
.B(n_1972),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_12617),
.B(n_1972),
.Y(n_12765)
);

AOI22xp5_ASAP7_75t_L g12766 ( 
.A1(n_12601),
.A2(n_1975),
.B1(n_1973),
.B2(n_1974),
.Y(n_12766)
);

AND2x2_ASAP7_75t_L g12767 ( 
.A(n_12573),
.B(n_1973),
.Y(n_12767)
);

AND2x2_ASAP7_75t_L g12768 ( 
.A(n_12609),
.B(n_12575),
.Y(n_12768)
);

OAI22xp5_ASAP7_75t_L g12769 ( 
.A1(n_12639),
.A2(n_1977),
.B1(n_1974),
.B2(n_1976),
.Y(n_12769)
);

OAI21xp5_ASAP7_75t_SL g12770 ( 
.A1(n_12638),
.A2(n_1976),
.B(n_1977),
.Y(n_12770)
);

NAND3xp33_ASAP7_75t_L g12771 ( 
.A(n_12481),
.B(n_1978),
.C(n_1979),
.Y(n_12771)
);

AND2x2_ASAP7_75t_L g12772 ( 
.A(n_12613),
.B(n_1978),
.Y(n_12772)
);

NAND2xp5_ASAP7_75t_L g12773 ( 
.A(n_12615),
.B(n_1979),
.Y(n_12773)
);

AND2x2_ASAP7_75t_L g12774 ( 
.A(n_12620),
.B(n_1980),
.Y(n_12774)
);

NAND2xp5_ASAP7_75t_L g12775 ( 
.A(n_12647),
.B(n_1980),
.Y(n_12775)
);

AND2x2_ASAP7_75t_L g12776 ( 
.A(n_12602),
.B(n_12612),
.Y(n_12776)
);

OAI21xp5_ASAP7_75t_SL g12777 ( 
.A1(n_12514),
.A2(n_1981),
.B(n_1982),
.Y(n_12777)
);

AND2x2_ASAP7_75t_L g12778 ( 
.A(n_12538),
.B(n_1982),
.Y(n_12778)
);

OAI21xp5_ASAP7_75t_SL g12779 ( 
.A1(n_12515),
.A2(n_1983),
.B(n_1984),
.Y(n_12779)
);

INVx2_ASAP7_75t_L g12780 ( 
.A(n_12632),
.Y(n_12780)
);

OAI22xp5_ASAP7_75t_L g12781 ( 
.A1(n_12518),
.A2(n_1985),
.B1(n_1983),
.B2(n_1984),
.Y(n_12781)
);

AND2x2_ASAP7_75t_L g12782 ( 
.A(n_12519),
.B(n_1985),
.Y(n_12782)
);

NAND2xp5_ASAP7_75t_L g12783 ( 
.A(n_12542),
.B(n_1986),
.Y(n_12783)
);

NOR3xp33_ASAP7_75t_SL g12784 ( 
.A(n_12649),
.B(n_1986),
.C(n_1987),
.Y(n_12784)
);

AND2x2_ASAP7_75t_L g12785 ( 
.A(n_12547),
.B(n_12555),
.Y(n_12785)
);

OAI21xp33_ASAP7_75t_SL g12786 ( 
.A1(n_12486),
.A2(n_1988),
.B(n_1989),
.Y(n_12786)
);

NAND2xp5_ASAP7_75t_L g12787 ( 
.A(n_12528),
.B(n_1988),
.Y(n_12787)
);

AOI211xp5_ASAP7_75t_L g12788 ( 
.A1(n_12598),
.A2(n_1991),
.B(n_1989),
.C(n_1990),
.Y(n_12788)
);

NAND2xp5_ASAP7_75t_L g12789 ( 
.A(n_12520),
.B(n_1990),
.Y(n_12789)
);

OAI221xp5_ASAP7_75t_L g12790 ( 
.A1(n_12523),
.A2(n_1993),
.B1(n_1991),
.B2(n_1992),
.C(n_1994),
.Y(n_12790)
);

NAND3xp33_ASAP7_75t_L g12791 ( 
.A(n_12535),
.B(n_1992),
.C(n_1993),
.Y(n_12791)
);

AND2x2_ASAP7_75t_L g12792 ( 
.A(n_12489),
.B(n_1995),
.Y(n_12792)
);

AND2x2_ASAP7_75t_L g12793 ( 
.A(n_12490),
.B(n_1996),
.Y(n_12793)
);

AND2x2_ASAP7_75t_L g12794 ( 
.A(n_12492),
.B(n_1996),
.Y(n_12794)
);

NAND2xp5_ASAP7_75t_L g12795 ( 
.A(n_12625),
.B(n_1997),
.Y(n_12795)
);

OAI221xp5_ASAP7_75t_L g12796 ( 
.A1(n_12630),
.A2(n_2000),
.B1(n_1998),
.B2(n_1999),
.C(n_2001),
.Y(n_12796)
);

AND2x2_ASAP7_75t_L g12797 ( 
.A(n_12497),
.B(n_1998),
.Y(n_12797)
);

AND2x2_ASAP7_75t_L g12798 ( 
.A(n_12512),
.B(n_2000),
.Y(n_12798)
);

NAND2xp5_ASAP7_75t_L g12799 ( 
.A(n_12635),
.B(n_2001),
.Y(n_12799)
);

AND2x2_ASAP7_75t_SL g12800 ( 
.A(n_12507),
.B(n_2002),
.Y(n_12800)
);

NAND2xp5_ASAP7_75t_L g12801 ( 
.A(n_12525),
.B(n_2002),
.Y(n_12801)
);

NAND3xp33_ASAP7_75t_L g12802 ( 
.A(n_12645),
.B(n_2003),
.C(n_2005),
.Y(n_12802)
);

AOI22xp33_ASAP7_75t_SL g12803 ( 
.A1(n_12626),
.A2(n_12648),
.B1(n_12468),
.B2(n_12513),
.Y(n_12803)
);

NOR2xp33_ASAP7_75t_L g12804 ( 
.A(n_12622),
.B(n_2003),
.Y(n_12804)
);

AND2x2_ASAP7_75t_L g12805 ( 
.A(n_12624),
.B(n_2005),
.Y(n_12805)
);

HB1xp67_ASAP7_75t_L g12806 ( 
.A(n_12628),
.Y(n_12806)
);

OAI21xp5_ASAP7_75t_L g12807 ( 
.A1(n_12595),
.A2(n_2006),
.B(n_2007),
.Y(n_12807)
);

INVx1_ASAP7_75t_L g12808 ( 
.A(n_12674),
.Y(n_12808)
);

INVx2_ASAP7_75t_L g12809 ( 
.A(n_12658),
.Y(n_12809)
);

AND2x2_ASAP7_75t_L g12810 ( 
.A(n_12710),
.B(n_12619),
.Y(n_12810)
);

HB1xp67_ASAP7_75t_L g12811 ( 
.A(n_12679),
.Y(n_12811)
);

AND2x2_ASAP7_75t_L g12812 ( 
.A(n_12656),
.B(n_12631),
.Y(n_12812)
);

INVx2_ASAP7_75t_L g12813 ( 
.A(n_12693),
.Y(n_12813)
);

BUFx2_ASAP7_75t_L g12814 ( 
.A(n_12786),
.Y(n_12814)
);

AND2x2_ASAP7_75t_L g12815 ( 
.A(n_12653),
.B(n_12634),
.Y(n_12815)
);

AND2x2_ASAP7_75t_L g12816 ( 
.A(n_12663),
.B(n_12690),
.Y(n_12816)
);

OR2x2_ASAP7_75t_L g12817 ( 
.A(n_12654),
.B(n_12549),
.Y(n_12817)
);

AND2x2_ASAP7_75t_L g12818 ( 
.A(n_12763),
.B(n_12511),
.Y(n_12818)
);

NOR2x1_ASAP7_75t_L g12819 ( 
.A(n_12736),
.B(n_12557),
.Y(n_12819)
);

AND2x2_ASAP7_75t_L g12820 ( 
.A(n_12768),
.B(n_12562),
.Y(n_12820)
);

AND2x2_ASAP7_75t_L g12821 ( 
.A(n_12670),
.B(n_12572),
.Y(n_12821)
);

HB1xp67_ASAP7_75t_L g12822 ( 
.A(n_12679),
.Y(n_12822)
);

INVx1_ASAP7_75t_L g12823 ( 
.A(n_12719),
.Y(n_12823)
);

INVx2_ASAP7_75t_L g12824 ( 
.A(n_12725),
.Y(n_12824)
);

AND2x2_ASAP7_75t_L g12825 ( 
.A(n_12659),
.B(n_12576),
.Y(n_12825)
);

NAND2xp5_ASAP7_75t_L g12826 ( 
.A(n_12704),
.B(n_12578),
.Y(n_12826)
);

OR2x2_ASAP7_75t_L g12827 ( 
.A(n_12695),
.B(n_12567),
.Y(n_12827)
);

INVx1_ASAP7_75t_L g12828 ( 
.A(n_12661),
.Y(n_12828)
);

NAND2xp5_ASAP7_75t_L g12829 ( 
.A(n_12701),
.B(n_12579),
.Y(n_12829)
);

NAND2xp5_ASAP7_75t_L g12830 ( 
.A(n_12669),
.B(n_12800),
.Y(n_12830)
);

AND2x2_ASAP7_75t_L g12831 ( 
.A(n_12686),
.B(n_12590),
.Y(n_12831)
);

INVx1_ASAP7_75t_L g12832 ( 
.A(n_12806),
.Y(n_12832)
);

AND2x2_ASAP7_75t_L g12833 ( 
.A(n_12666),
.B(n_12592),
.Y(n_12833)
);

AND2x2_ASAP7_75t_L g12834 ( 
.A(n_12682),
.B(n_12594),
.Y(n_12834)
);

BUFx3_ASAP7_75t_L g12835 ( 
.A(n_12730),
.Y(n_12835)
);

INVx1_ASAP7_75t_L g12836 ( 
.A(n_12731),
.Y(n_12836)
);

AND2x2_ASAP7_75t_L g12837 ( 
.A(n_12780),
.B(n_12597),
.Y(n_12837)
);

AND2x4_ASAP7_75t_L g12838 ( 
.A(n_12749),
.B(n_12568),
.Y(n_12838)
);

INVx1_ASAP7_75t_L g12839 ( 
.A(n_12716),
.Y(n_12839)
);

INVx1_ASAP7_75t_L g12840 ( 
.A(n_12672),
.Y(n_12840)
);

NAND2xp5_ASAP7_75t_L g12841 ( 
.A(n_12685),
.B(n_12718),
.Y(n_12841)
);

AND2x2_ASAP7_75t_L g12842 ( 
.A(n_12687),
.B(n_12582),
.Y(n_12842)
);

OR2x2_ASAP7_75t_L g12843 ( 
.A(n_12664),
.B(n_2007),
.Y(n_12843)
);

AND2x4_ASAP7_75t_L g12844 ( 
.A(n_12776),
.B(n_2008),
.Y(n_12844)
);

AND2x2_ASAP7_75t_L g12845 ( 
.A(n_12785),
.B(n_2008),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_12702),
.B(n_2009),
.Y(n_12846)
);

AND2x2_ASAP7_75t_L g12847 ( 
.A(n_12707),
.B(n_2009),
.Y(n_12847)
);

INVx2_ASAP7_75t_L g12848 ( 
.A(n_12758),
.Y(n_12848)
);

INVx1_ASAP7_75t_L g12849 ( 
.A(n_12752),
.Y(n_12849)
);

AND2x4_ASAP7_75t_L g12850 ( 
.A(n_12778),
.B(n_2010),
.Y(n_12850)
);

AND2x2_ASAP7_75t_L g12851 ( 
.A(n_12760),
.B(n_2010),
.Y(n_12851)
);

INVx1_ASAP7_75t_L g12852 ( 
.A(n_12751),
.Y(n_12852)
);

AND2x4_ASAP7_75t_L g12853 ( 
.A(n_12762),
.B(n_2011),
.Y(n_12853)
);

AND2x2_ASAP7_75t_L g12854 ( 
.A(n_12689),
.B(n_2012),
.Y(n_12854)
);

CKINVDCx14_ASAP7_75t_R g12855 ( 
.A(n_12805),
.Y(n_12855)
);

INVx2_ASAP7_75t_L g12856 ( 
.A(n_12714),
.Y(n_12856)
);

INVx2_ASAP7_75t_L g12857 ( 
.A(n_12744),
.Y(n_12857)
);

INVx1_ASAP7_75t_L g12858 ( 
.A(n_12706),
.Y(n_12858)
);

OR2x2_ASAP7_75t_L g12859 ( 
.A(n_12677),
.B(n_2012),
.Y(n_12859)
);

INVx1_ASAP7_75t_L g12860 ( 
.A(n_12792),
.Y(n_12860)
);

INVx1_ASAP7_75t_L g12861 ( 
.A(n_12793),
.Y(n_12861)
);

AND2x2_ASAP7_75t_L g12862 ( 
.A(n_12696),
.B(n_12673),
.Y(n_12862)
);

INVx3_ASAP7_75t_L g12863 ( 
.A(n_12747),
.Y(n_12863)
);

INVx2_ASAP7_75t_L g12864 ( 
.A(n_12794),
.Y(n_12864)
);

INVx1_ASAP7_75t_SL g12865 ( 
.A(n_12688),
.Y(n_12865)
);

INVx1_ASAP7_75t_L g12866 ( 
.A(n_12797),
.Y(n_12866)
);

INVx2_ASAP7_75t_L g12867 ( 
.A(n_12798),
.Y(n_12867)
);

OR2x2_ASAP7_75t_L g12868 ( 
.A(n_12684),
.B(n_2013),
.Y(n_12868)
);

NOR2xp67_ASAP7_75t_L g12869 ( 
.A(n_12703),
.B(n_2014),
.Y(n_12869)
);

AND2x2_ASAP7_75t_L g12870 ( 
.A(n_12782),
.B(n_2015),
.Y(n_12870)
);

OR2x2_ASAP7_75t_L g12871 ( 
.A(n_12680),
.B(n_2015),
.Y(n_12871)
);

AND2x2_ASAP7_75t_L g12872 ( 
.A(n_12665),
.B(n_2016),
.Y(n_12872)
);

HB1xp67_ASAP7_75t_L g12873 ( 
.A(n_12705),
.Y(n_12873)
);

NAND2xp5_ASAP7_75t_L g12874 ( 
.A(n_12708),
.B(n_2016),
.Y(n_12874)
);

AND2x2_ASAP7_75t_L g12875 ( 
.A(n_12764),
.B(n_2017),
.Y(n_12875)
);

NAND2xp5_ASAP7_75t_L g12876 ( 
.A(n_12705),
.B(n_2018),
.Y(n_12876)
);

AND2x4_ASAP7_75t_L g12877 ( 
.A(n_12767),
.B(n_2018),
.Y(n_12877)
);

AND2x2_ASAP7_75t_L g12878 ( 
.A(n_12772),
.B(n_2019),
.Y(n_12878)
);

BUFx2_ASAP7_75t_L g12879 ( 
.A(n_12709),
.Y(n_12879)
);

AND2x2_ASAP7_75t_L g12880 ( 
.A(n_12774),
.B(n_2019),
.Y(n_12880)
);

INVx1_ASAP7_75t_L g12881 ( 
.A(n_12734),
.Y(n_12881)
);

AND2x2_ASAP7_75t_L g12882 ( 
.A(n_12657),
.B(n_2020),
.Y(n_12882)
);

INVx2_ASAP7_75t_L g12883 ( 
.A(n_12721),
.Y(n_12883)
);

HB1xp67_ASAP7_75t_L g12884 ( 
.A(n_12709),
.Y(n_12884)
);

AND2x4_ASAP7_75t_L g12885 ( 
.A(n_12711),
.B(n_2021),
.Y(n_12885)
);

BUFx2_ASAP7_75t_L g12886 ( 
.A(n_12728),
.Y(n_12886)
);

INVx1_ASAP7_75t_L g12887 ( 
.A(n_12723),
.Y(n_12887)
);

OR2x2_ASAP7_75t_L g12888 ( 
.A(n_12681),
.B(n_2021),
.Y(n_12888)
);

INVx1_ASAP7_75t_L g12889 ( 
.A(n_12750),
.Y(n_12889)
);

AND2x2_ASAP7_75t_L g12890 ( 
.A(n_12694),
.B(n_2022),
.Y(n_12890)
);

AND2x4_ASAP7_75t_L g12891 ( 
.A(n_12724),
.B(n_2023),
.Y(n_12891)
);

OR2x2_ASAP7_75t_L g12892 ( 
.A(n_12671),
.B(n_2023),
.Y(n_12892)
);

INVx1_ASAP7_75t_L g12893 ( 
.A(n_12713),
.Y(n_12893)
);

AOI22xp33_ASAP7_75t_L g12894 ( 
.A1(n_12655),
.A2(n_2026),
.B1(n_2024),
.B2(n_2025),
.Y(n_12894)
);

AND2x2_ASAP7_75t_L g12895 ( 
.A(n_12692),
.B(n_2025),
.Y(n_12895)
);

NAND2xp5_ASAP7_75t_L g12896 ( 
.A(n_12660),
.B(n_2026),
.Y(n_12896)
);

OR2x2_ASAP7_75t_L g12897 ( 
.A(n_12765),
.B(n_2027),
.Y(n_12897)
);

NAND2xp5_ASAP7_75t_L g12898 ( 
.A(n_12770),
.B(n_2027),
.Y(n_12898)
);

AND2x2_ASAP7_75t_L g12899 ( 
.A(n_12740),
.B(n_2028),
.Y(n_12899)
);

AND2x2_ASAP7_75t_L g12900 ( 
.A(n_12699),
.B(n_12803),
.Y(n_12900)
);

INVx1_ASAP7_75t_L g12901 ( 
.A(n_12773),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12712),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_12739),
.Y(n_12903)
);

INVx1_ASAP7_75t_L g12904 ( 
.A(n_12737),
.Y(n_12904)
);

INVx1_ASAP7_75t_L g12905 ( 
.A(n_12801),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_12789),
.Y(n_12906)
);

AND2x2_ASAP7_75t_L g12907 ( 
.A(n_12732),
.B(n_12697),
.Y(n_12907)
);

INVx1_ASAP7_75t_L g12908 ( 
.A(n_12795),
.Y(n_12908)
);

NAND2xp5_ASAP7_75t_L g12909 ( 
.A(n_12729),
.B(n_2028),
.Y(n_12909)
);

AND2x2_ASAP7_75t_L g12910 ( 
.A(n_12807),
.B(n_2029),
.Y(n_12910)
);

INVx1_ASAP7_75t_L g12911 ( 
.A(n_12799),
.Y(n_12911)
);

NOR2x1_ASAP7_75t_L g12912 ( 
.A(n_12746),
.B(n_2029),
.Y(n_12912)
);

INVx1_ASAP7_75t_L g12913 ( 
.A(n_12783),
.Y(n_12913)
);

OR2x2_ASAP7_75t_L g12914 ( 
.A(n_12668),
.B(n_2030),
.Y(n_12914)
);

OR2x2_ASAP7_75t_L g12915 ( 
.A(n_12676),
.B(n_2031),
.Y(n_12915)
);

OR2x2_ASAP7_75t_L g12916 ( 
.A(n_12675),
.B(n_2031),
.Y(n_12916)
);

AND2x2_ASAP7_75t_L g12917 ( 
.A(n_12784),
.B(n_2032),
.Y(n_12917)
);

AND2x4_ASAP7_75t_L g12918 ( 
.A(n_12745),
.B(n_2032),
.Y(n_12918)
);

AND2x2_ASAP7_75t_L g12919 ( 
.A(n_12804),
.B(n_2033),
.Y(n_12919)
);

AND2x2_ASAP7_75t_L g12920 ( 
.A(n_12787),
.B(n_2033),
.Y(n_12920)
);

INVx1_ASAP7_75t_L g12921 ( 
.A(n_12775),
.Y(n_12921)
);

INVx3_ASAP7_75t_L g12922 ( 
.A(n_12698),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12769),
.Y(n_12923)
);

NOR2xp33_ASAP7_75t_L g12924 ( 
.A(n_12678),
.B(n_2034),
.Y(n_12924)
);

INVx2_ASAP7_75t_L g12925 ( 
.A(n_12756),
.Y(n_12925)
);

NAND2xp5_ASAP7_75t_L g12926 ( 
.A(n_12777),
.B(n_2035),
.Y(n_12926)
);

HB1xp67_ASAP7_75t_L g12927 ( 
.A(n_12755),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12738),
.Y(n_12928)
);

INVxp67_ASAP7_75t_L g12929 ( 
.A(n_12662),
.Y(n_12929)
);

INVx1_ASAP7_75t_L g12930 ( 
.A(n_12753),
.Y(n_12930)
);

AND2x2_ASAP7_75t_L g12931 ( 
.A(n_12722),
.B(n_2035),
.Y(n_12931)
);

INVx1_ASAP7_75t_L g12932 ( 
.A(n_12791),
.Y(n_12932)
);

AND2x4_ASAP7_75t_SL g12933 ( 
.A(n_12757),
.B(n_2036),
.Y(n_12933)
);

NAND2xp5_ASAP7_75t_L g12934 ( 
.A(n_12779),
.B(n_2036),
.Y(n_12934)
);

INVx2_ASAP7_75t_L g12935 ( 
.A(n_12743),
.Y(n_12935)
);

AND2x2_ASAP7_75t_L g12936 ( 
.A(n_12715),
.B(n_2037),
.Y(n_12936)
);

INVx1_ASAP7_75t_L g12937 ( 
.A(n_12771),
.Y(n_12937)
);

INVx1_ASAP7_75t_L g12938 ( 
.A(n_12802),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12766),
.Y(n_12939)
);

INVx1_ASAP7_75t_L g12940 ( 
.A(n_12811),
.Y(n_12940)
);

INVx1_ASAP7_75t_L g12941 ( 
.A(n_12822),
.Y(n_12941)
);

INVx2_ASAP7_75t_SL g12942 ( 
.A(n_12838),
.Y(n_12942)
);

NAND2xp5_ASAP7_75t_L g12943 ( 
.A(n_12873),
.B(n_12683),
.Y(n_12943)
);

INVx1_ASAP7_75t_L g12944 ( 
.A(n_12884),
.Y(n_12944)
);

OAI21xp5_ASAP7_75t_L g12945 ( 
.A1(n_12869),
.A2(n_12667),
.B(n_12700),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12879),
.Y(n_12946)
);

NAND2xp5_ASAP7_75t_L g12947 ( 
.A(n_12816),
.B(n_12691),
.Y(n_12947)
);

INVx1_ASAP7_75t_L g12948 ( 
.A(n_12845),
.Y(n_12948)
);

INVx2_ASAP7_75t_SL g12949 ( 
.A(n_12810),
.Y(n_12949)
);

NAND2xp5_ASAP7_75t_SL g12950 ( 
.A(n_12814),
.B(n_12788),
.Y(n_12950)
);

INVx1_ASAP7_75t_L g12951 ( 
.A(n_12823),
.Y(n_12951)
);

INVx1_ASAP7_75t_L g12952 ( 
.A(n_12831),
.Y(n_12952)
);

INVx1_ASAP7_75t_L g12953 ( 
.A(n_12825),
.Y(n_12953)
);

INVx4_ASAP7_75t_SL g12954 ( 
.A(n_12844),
.Y(n_12954)
);

HB1xp67_ASAP7_75t_L g12955 ( 
.A(n_12855),
.Y(n_12955)
);

INVx1_ASAP7_75t_L g12956 ( 
.A(n_12818),
.Y(n_12956)
);

AND2x2_ASAP7_75t_L g12957 ( 
.A(n_12809),
.B(n_12754),
.Y(n_12957)
);

OAI21x1_ASAP7_75t_L g12958 ( 
.A1(n_12922),
.A2(n_12741),
.B(n_12781),
.Y(n_12958)
);

NOR2x1p5_ASAP7_75t_L g12959 ( 
.A(n_12841),
.B(n_12726),
.Y(n_12959)
);

BUFx2_ASAP7_75t_L g12960 ( 
.A(n_12842),
.Y(n_12960)
);

INVx1_ASAP7_75t_L g12961 ( 
.A(n_12820),
.Y(n_12961)
);

INVx1_ASAP7_75t_L g12962 ( 
.A(n_12851),
.Y(n_12962)
);

OA21x2_ASAP7_75t_L g12963 ( 
.A1(n_12876),
.A2(n_12733),
.B(n_12727),
.Y(n_12963)
);

INVx2_ASAP7_75t_L g12964 ( 
.A(n_12835),
.Y(n_12964)
);

NAND2xp5_ASAP7_75t_L g12965 ( 
.A(n_12865),
.B(n_12759),
.Y(n_12965)
);

HB1xp67_ASAP7_75t_L g12966 ( 
.A(n_12833),
.Y(n_12966)
);

INVx1_ASAP7_75t_L g12967 ( 
.A(n_12870),
.Y(n_12967)
);

HB1xp67_ASAP7_75t_L g12968 ( 
.A(n_12832),
.Y(n_12968)
);

AND2x2_ASAP7_75t_L g12969 ( 
.A(n_12813),
.B(n_12761),
.Y(n_12969)
);

INVx4_ASAP7_75t_L g12970 ( 
.A(n_12877),
.Y(n_12970)
);

OA21x2_ASAP7_75t_L g12971 ( 
.A1(n_12826),
.A2(n_12717),
.B(n_12748),
.Y(n_12971)
);

AOI21x1_ASAP7_75t_L g12972 ( 
.A1(n_12900),
.A2(n_12735),
.B(n_12742),
.Y(n_12972)
);

INVx2_ASAP7_75t_L g12973 ( 
.A(n_12863),
.Y(n_12973)
);

INVx1_ASAP7_75t_L g12974 ( 
.A(n_12875),
.Y(n_12974)
);

NOR2x1_ASAP7_75t_L g12975 ( 
.A(n_12915),
.B(n_12720),
.Y(n_12975)
);

NAND2xp5_ASAP7_75t_L g12976 ( 
.A(n_12890),
.B(n_12862),
.Y(n_12976)
);

INVx1_ASAP7_75t_L g12977 ( 
.A(n_12878),
.Y(n_12977)
);

NOR2xp67_ASAP7_75t_SL g12978 ( 
.A(n_12843),
.B(n_12790),
.Y(n_12978)
);

INVx1_ASAP7_75t_L g12979 ( 
.A(n_12880),
.Y(n_12979)
);

BUFx6f_ASAP7_75t_L g12980 ( 
.A(n_12850),
.Y(n_12980)
);

OAI21xp5_ASAP7_75t_L g12981 ( 
.A1(n_12929),
.A2(n_12796),
.B(n_2038),
.Y(n_12981)
);

NOR2x1p5_ASAP7_75t_L g12982 ( 
.A(n_12830),
.B(n_2038),
.Y(n_12982)
);

AND2x2_ASAP7_75t_L g12983 ( 
.A(n_12834),
.B(n_2039),
.Y(n_12983)
);

OAI21x1_ASAP7_75t_L g12984 ( 
.A1(n_12819),
.A2(n_2039),
.B(n_2040),
.Y(n_12984)
);

AND2x2_ASAP7_75t_L g12985 ( 
.A(n_12815),
.B(n_2040),
.Y(n_12985)
);

AND2x2_ASAP7_75t_L g12986 ( 
.A(n_12821),
.B(n_2041),
.Y(n_12986)
);

NOR2x1p5_ASAP7_75t_L g12987 ( 
.A(n_12829),
.B(n_2042),
.Y(n_12987)
);

OAI21x1_ASAP7_75t_L g12988 ( 
.A1(n_12912),
.A2(n_2042),
.B(n_2043),
.Y(n_12988)
);

INVx1_ASAP7_75t_L g12989 ( 
.A(n_12836),
.Y(n_12989)
);

INVx4_ASAP7_75t_SL g12990 ( 
.A(n_12872),
.Y(n_12990)
);

AND2x4_ASAP7_75t_L g12991 ( 
.A(n_12812),
.B(n_2043),
.Y(n_12991)
);

INVx2_ASAP7_75t_L g12992 ( 
.A(n_12853),
.Y(n_12992)
);

INVxp67_ASAP7_75t_L g12993 ( 
.A(n_12924),
.Y(n_12993)
);

OAI21x1_ASAP7_75t_L g12994 ( 
.A1(n_12817),
.A2(n_2044),
.B(n_2045),
.Y(n_12994)
);

INVxp67_ASAP7_75t_SL g12995 ( 
.A(n_12927),
.Y(n_12995)
);

INVx2_ASAP7_75t_L g12996 ( 
.A(n_12824),
.Y(n_12996)
);

INVx3_ASAP7_75t_L g12997 ( 
.A(n_12885),
.Y(n_12997)
);

INVx1_ASAP7_75t_SL g12998 ( 
.A(n_12891),
.Y(n_12998)
);

INVx2_ASAP7_75t_L g12999 ( 
.A(n_12848),
.Y(n_12999)
);

INVx1_ASAP7_75t_L g13000 ( 
.A(n_12839),
.Y(n_13000)
);

INVx2_ASAP7_75t_L g13001 ( 
.A(n_12864),
.Y(n_13001)
);

BUFx8_ASAP7_75t_L g13002 ( 
.A(n_12854),
.Y(n_13002)
);

BUFx8_ASAP7_75t_L g13003 ( 
.A(n_12919),
.Y(n_13003)
);

INVx1_ASAP7_75t_L g13004 ( 
.A(n_12837),
.Y(n_13004)
);

INVx1_ASAP7_75t_L g13005 ( 
.A(n_12849),
.Y(n_13005)
);

INVx1_ASAP7_75t_L g13006 ( 
.A(n_12852),
.Y(n_13006)
);

INVx3_ASAP7_75t_L g13007 ( 
.A(n_12918),
.Y(n_13007)
);

HB1xp67_ASAP7_75t_L g13008 ( 
.A(n_12840),
.Y(n_13008)
);

OA21x2_ASAP7_75t_L g13009 ( 
.A1(n_12896),
.A2(n_2044),
.B(n_2046),
.Y(n_13009)
);

INVx2_ASAP7_75t_L g13010 ( 
.A(n_12867),
.Y(n_13010)
);

INVxp67_ASAP7_75t_SL g13011 ( 
.A(n_12827),
.Y(n_13011)
);

INVx1_ASAP7_75t_L g13012 ( 
.A(n_12860),
.Y(n_13012)
);

INVx2_ASAP7_75t_L g13013 ( 
.A(n_12857),
.Y(n_13013)
);

AND2x2_ASAP7_75t_L g13014 ( 
.A(n_12856),
.B(n_2046),
.Y(n_13014)
);

INVx4_ASAP7_75t_SL g13015 ( 
.A(n_12920),
.Y(n_13015)
);

NAND4xp25_ASAP7_75t_L g13016 ( 
.A(n_12923),
.B(n_2051),
.C(n_2047),
.D(n_2050),
.Y(n_13016)
);

NAND3xp33_ASAP7_75t_SL g13017 ( 
.A(n_12914),
.B(n_12916),
.C(n_12847),
.Y(n_13017)
);

OA21x2_ASAP7_75t_L g13018 ( 
.A1(n_12846),
.A2(n_2047),
.B(n_2051),
.Y(n_13018)
);

INVx1_ASAP7_75t_L g13019 ( 
.A(n_12861),
.Y(n_13019)
);

INVx2_ASAP7_75t_L g13020 ( 
.A(n_12866),
.Y(n_13020)
);

AO21x1_ASAP7_75t_L g13021 ( 
.A1(n_12882),
.A2(n_2052),
.B(n_2053),
.Y(n_13021)
);

AO21x1_ASAP7_75t_L g13022 ( 
.A1(n_12895),
.A2(n_12892),
.B(n_12871),
.Y(n_13022)
);

AO21x2_ASAP7_75t_L g13023 ( 
.A1(n_12899),
.A2(n_2052),
.B(n_2053),
.Y(n_13023)
);

INVx2_ASAP7_75t_L g13024 ( 
.A(n_12808),
.Y(n_13024)
);

INVx2_ASAP7_75t_L g13025 ( 
.A(n_12897),
.Y(n_13025)
);

AND2x2_ASAP7_75t_L g13026 ( 
.A(n_12925),
.B(n_2054),
.Y(n_13026)
);

INVx1_ASAP7_75t_L g13027 ( 
.A(n_12828),
.Y(n_13027)
);

NOR2xp33_ASAP7_75t_L g13028 ( 
.A(n_12868),
.B(n_2054),
.Y(n_13028)
);

OAI21xp5_ASAP7_75t_L g13029 ( 
.A1(n_12928),
.A2(n_12907),
.B(n_12932),
.Y(n_13029)
);

OA21x2_ASAP7_75t_L g13030 ( 
.A1(n_12874),
.A2(n_2055),
.B(n_2056),
.Y(n_13030)
);

NAND2xp5_ASAP7_75t_SL g13031 ( 
.A(n_12935),
.B(n_2056),
.Y(n_13031)
);

OAI21xp5_ASAP7_75t_L g13032 ( 
.A1(n_12930),
.A2(n_12937),
.B(n_12938),
.Y(n_13032)
);

BUFx2_ASAP7_75t_L g13033 ( 
.A(n_12886),
.Y(n_13033)
);

INVxp67_ASAP7_75t_L g13034 ( 
.A(n_12917),
.Y(n_13034)
);

INVx1_ASAP7_75t_L g13035 ( 
.A(n_12904),
.Y(n_13035)
);

HB1xp67_ASAP7_75t_L g13036 ( 
.A(n_12888),
.Y(n_13036)
);

AND2x2_ASAP7_75t_L g13037 ( 
.A(n_12933),
.B(n_2057),
.Y(n_13037)
);

INVxp67_ASAP7_75t_L g13038 ( 
.A(n_12936),
.Y(n_13038)
);

INVx1_ASAP7_75t_SL g13039 ( 
.A(n_12859),
.Y(n_13039)
);

INVxp67_ASAP7_75t_SL g13040 ( 
.A(n_12909),
.Y(n_13040)
);

INVx1_ASAP7_75t_L g13041 ( 
.A(n_12887),
.Y(n_13041)
);

INVx1_ASAP7_75t_L g13042 ( 
.A(n_12883),
.Y(n_13042)
);

INVx1_ASAP7_75t_L g13043 ( 
.A(n_12902),
.Y(n_13043)
);

OA21x2_ASAP7_75t_L g13044 ( 
.A1(n_12898),
.A2(n_2057),
.B(n_2058),
.Y(n_13044)
);

HB1xp67_ASAP7_75t_L g13045 ( 
.A(n_12910),
.Y(n_13045)
);

INVx1_ASAP7_75t_L g13046 ( 
.A(n_12903),
.Y(n_13046)
);

INVx3_ASAP7_75t_L g13047 ( 
.A(n_12901),
.Y(n_13047)
);

AND2x2_ASAP7_75t_L g13048 ( 
.A(n_12939),
.B(n_2058),
.Y(n_13048)
);

AND2x2_ASAP7_75t_L g13049 ( 
.A(n_12858),
.B(n_2059),
.Y(n_13049)
);

INVx2_ASAP7_75t_SL g13050 ( 
.A(n_12931),
.Y(n_13050)
);

INVx2_ASAP7_75t_SL g13051 ( 
.A(n_12926),
.Y(n_13051)
);

NOR3xp33_ASAP7_75t_SL g13052 ( 
.A(n_12889),
.B(n_2059),
.C(n_2060),
.Y(n_13052)
);

AOI21x1_ASAP7_75t_L g13053 ( 
.A1(n_12934),
.A2(n_2060),
.B(n_2061),
.Y(n_13053)
);

BUFx8_ASAP7_75t_L g13054 ( 
.A(n_12893),
.Y(n_13054)
);

OR2x2_ASAP7_75t_L g13055 ( 
.A(n_12960),
.B(n_12881),
.Y(n_13055)
);

INVx1_ASAP7_75t_L g13056 ( 
.A(n_12955),
.Y(n_13056)
);

INVx1_ASAP7_75t_L g13057 ( 
.A(n_12966),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12968),
.Y(n_13058)
);

INVx2_ASAP7_75t_L g13059 ( 
.A(n_12954),
.Y(n_13059)
);

INVx2_ASAP7_75t_L g13060 ( 
.A(n_12954),
.Y(n_13060)
);

AND2x2_ASAP7_75t_L g13061 ( 
.A(n_12942),
.B(n_12913),
.Y(n_13061)
);

AND2x2_ASAP7_75t_L g13062 ( 
.A(n_13015),
.B(n_12906),
.Y(n_13062)
);

NAND2xp5_ASAP7_75t_L g13063 ( 
.A(n_12949),
.B(n_12894),
.Y(n_13063)
);

INVx1_ASAP7_75t_L g13064 ( 
.A(n_13033),
.Y(n_13064)
);

NAND2x1_ASAP7_75t_L g13065 ( 
.A(n_12970),
.B(n_12921),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_13008),
.Y(n_13066)
);

AND2x2_ASAP7_75t_L g13067 ( 
.A(n_13015),
.B(n_12908),
.Y(n_13067)
);

AND2x2_ASAP7_75t_L g13068 ( 
.A(n_12990),
.B(n_12911),
.Y(n_13068)
);

INVx1_ASAP7_75t_L g13069 ( 
.A(n_12944),
.Y(n_13069)
);

INVx1_ASAP7_75t_L g13070 ( 
.A(n_12946),
.Y(n_13070)
);

AND2x2_ASAP7_75t_L g13071 ( 
.A(n_12990),
.B(n_12905),
.Y(n_13071)
);

HB1xp67_ASAP7_75t_L g13072 ( 
.A(n_13023),
.Y(n_13072)
);

NAND2xp5_ASAP7_75t_L g13073 ( 
.A(n_13002),
.B(n_2062),
.Y(n_13073)
);

NOR2x1p5_ASAP7_75t_L g13074 ( 
.A(n_13011),
.B(n_2062),
.Y(n_13074)
);

NAND2xp5_ASAP7_75t_L g13075 ( 
.A(n_13003),
.B(n_2063),
.Y(n_13075)
);

AND2x2_ASAP7_75t_L g13076 ( 
.A(n_12952),
.B(n_12995),
.Y(n_13076)
);

NAND2xp5_ASAP7_75t_L g13077 ( 
.A(n_12956),
.B(n_2065),
.Y(n_13077)
);

OR2x2_ASAP7_75t_L g13078 ( 
.A(n_12943),
.B(n_2065),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12983),
.Y(n_13079)
);

OR2x2_ASAP7_75t_L g13080 ( 
.A(n_12947),
.B(n_2066),
.Y(n_13080)
);

AND2x4_ASAP7_75t_L g13081 ( 
.A(n_12964),
.B(n_2066),
.Y(n_13081)
);

BUFx2_ASAP7_75t_L g13082 ( 
.A(n_12980),
.Y(n_13082)
);

INVx1_ASAP7_75t_L g13083 ( 
.A(n_12940),
.Y(n_13083)
);

AND2x2_ASAP7_75t_L g13084 ( 
.A(n_12992),
.B(n_2067),
.Y(n_13084)
);

INVx2_ASAP7_75t_L g13085 ( 
.A(n_12980),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12941),
.Y(n_13086)
);

INVxp67_ASAP7_75t_SL g13087 ( 
.A(n_13021),
.Y(n_13087)
);

AND2x2_ASAP7_75t_L g13088 ( 
.A(n_12961),
.B(n_2067),
.Y(n_13088)
);

INVx2_ASAP7_75t_L g13089 ( 
.A(n_12997),
.Y(n_13089)
);

BUFx2_ASAP7_75t_L g13090 ( 
.A(n_13018),
.Y(n_13090)
);

INVx1_ASAP7_75t_L g13091 ( 
.A(n_12985),
.Y(n_13091)
);

INVx1_ASAP7_75t_L g13092 ( 
.A(n_12986),
.Y(n_13092)
);

AND2x2_ASAP7_75t_L g13093 ( 
.A(n_12953),
.B(n_12973),
.Y(n_13093)
);

OR2x6_ASAP7_75t_L g13094 ( 
.A(n_12999),
.B(n_2068),
.Y(n_13094)
);

NAND2xp5_ASAP7_75t_L g13095 ( 
.A(n_13007),
.B(n_2068),
.Y(n_13095)
);

AND2x2_ASAP7_75t_L g13096 ( 
.A(n_12957),
.B(n_2069),
.Y(n_13096)
);

INVx1_ASAP7_75t_L g13097 ( 
.A(n_13037),
.Y(n_13097)
);

INVx4_ASAP7_75t_L g13098 ( 
.A(n_12991),
.Y(n_13098)
);

INVx1_ASAP7_75t_L g13099 ( 
.A(n_13045),
.Y(n_13099)
);

OR2x2_ASAP7_75t_L g13100 ( 
.A(n_12950),
.B(n_12976),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_13048),
.Y(n_13101)
);

AND2x2_ASAP7_75t_L g13102 ( 
.A(n_12998),
.B(n_2069),
.Y(n_13102)
);

OR2x2_ASAP7_75t_L g13103 ( 
.A(n_13017),
.B(n_2070),
.Y(n_13103)
);

NAND2xp5_ASAP7_75t_L g13104 ( 
.A(n_13004),
.B(n_2071),
.Y(n_13104)
);

AND2x2_ASAP7_75t_L g13105 ( 
.A(n_12962),
.B(n_2071),
.Y(n_13105)
);

INVx2_ASAP7_75t_L g13106 ( 
.A(n_12984),
.Y(n_13106)
);

NAND2xp5_ASAP7_75t_L g13107 ( 
.A(n_13034),
.B(n_2072),
.Y(n_13107)
);

INVx1_ASAP7_75t_L g13108 ( 
.A(n_13026),
.Y(n_13108)
);

INVx2_ASAP7_75t_L g13109 ( 
.A(n_12994),
.Y(n_13109)
);

INVx1_ASAP7_75t_L g13110 ( 
.A(n_13014),
.Y(n_13110)
);

NAND2xp5_ASAP7_75t_L g13111 ( 
.A(n_12948),
.B(n_2073),
.Y(n_13111)
);

INVx2_ASAP7_75t_L g13112 ( 
.A(n_12988),
.Y(n_13112)
);

OR2x2_ASAP7_75t_L g13113 ( 
.A(n_12967),
.B(n_2074),
.Y(n_13113)
);

INVx2_ASAP7_75t_L g13114 ( 
.A(n_12996),
.Y(n_13114)
);

AND2x2_ASAP7_75t_L g13115 ( 
.A(n_12969),
.B(n_2074),
.Y(n_13115)
);

AND2x2_ASAP7_75t_SL g13116 ( 
.A(n_12971),
.B(n_2075),
.Y(n_13116)
);

AND2x2_ASAP7_75t_L g13117 ( 
.A(n_12974),
.B(n_2076),
.Y(n_13117)
);

INVx1_ASAP7_75t_L g13118 ( 
.A(n_13036),
.Y(n_13118)
);

NAND2xp5_ASAP7_75t_L g13119 ( 
.A(n_12977),
.B(n_2076),
.Y(n_13119)
);

AND2x2_ASAP7_75t_L g13120 ( 
.A(n_12979),
.B(n_2077),
.Y(n_13120)
);

AND2x2_ASAP7_75t_L g13121 ( 
.A(n_12982),
.B(n_2077),
.Y(n_13121)
);

AND2x2_ASAP7_75t_L g13122 ( 
.A(n_13001),
.B(n_2078),
.Y(n_13122)
);

AND2x2_ASAP7_75t_L g13123 ( 
.A(n_13010),
.B(n_2078),
.Y(n_13123)
);

AND2x2_ASAP7_75t_L g13124 ( 
.A(n_13013),
.B(n_2079),
.Y(n_13124)
);

NOR2xp33_ASAP7_75t_SL g13125 ( 
.A(n_13039),
.B(n_2080),
.Y(n_13125)
);

AND2x4_ASAP7_75t_SL g13126 ( 
.A(n_13025),
.B(n_2081),
.Y(n_13126)
);

INVx1_ASAP7_75t_L g13127 ( 
.A(n_13049),
.Y(n_13127)
);

BUFx2_ASAP7_75t_L g13128 ( 
.A(n_13054),
.Y(n_13128)
);

INVx2_ASAP7_75t_L g13129 ( 
.A(n_12987),
.Y(n_13129)
);

OR2x2_ASAP7_75t_L g13130 ( 
.A(n_12965),
.B(n_2082),
.Y(n_13130)
);

BUFx2_ASAP7_75t_SL g13131 ( 
.A(n_13020),
.Y(n_13131)
);

AND2x2_ASAP7_75t_L g13132 ( 
.A(n_12958),
.B(n_2082),
.Y(n_13132)
);

AND2x2_ASAP7_75t_L g13133 ( 
.A(n_13029),
.B(n_2083),
.Y(n_13133)
);

NAND2xp5_ASAP7_75t_L g13134 ( 
.A(n_12945),
.B(n_2083),
.Y(n_13134)
);

INVx1_ASAP7_75t_L g13135 ( 
.A(n_12989),
.Y(n_13135)
);

HB1xp67_ASAP7_75t_L g13136 ( 
.A(n_13009),
.Y(n_13136)
);

AND2x2_ASAP7_75t_L g13137 ( 
.A(n_13038),
.B(n_2084),
.Y(n_13137)
);

AND2x2_ASAP7_75t_SL g13138 ( 
.A(n_12963),
.B(n_2084),
.Y(n_13138)
);

NOR2xp67_ASAP7_75t_L g13139 ( 
.A(n_13047),
.B(n_2085),
.Y(n_13139)
);

INVx1_ASAP7_75t_SL g13140 ( 
.A(n_13030),
.Y(n_13140)
);

AND2x2_ASAP7_75t_L g13141 ( 
.A(n_13050),
.B(n_2086),
.Y(n_13141)
);

INVx2_ASAP7_75t_L g13142 ( 
.A(n_13000),
.Y(n_13142)
);

INVx1_ASAP7_75t_L g13143 ( 
.A(n_13005),
.Y(n_13143)
);

NAND2xp5_ASAP7_75t_L g13144 ( 
.A(n_12978),
.B(n_2086),
.Y(n_13144)
);

AND2x4_ASAP7_75t_SL g13145 ( 
.A(n_13052),
.B(n_2087),
.Y(n_13145)
);

OR2x2_ASAP7_75t_L g13146 ( 
.A(n_13006),
.B(n_2087),
.Y(n_13146)
);

AND2x4_ASAP7_75t_L g13147 ( 
.A(n_13012),
.B(n_2088),
.Y(n_13147)
);

AND2x2_ASAP7_75t_L g13148 ( 
.A(n_13032),
.B(n_2088),
.Y(n_13148)
);

NAND2xp5_ASAP7_75t_L g13149 ( 
.A(n_12959),
.B(n_2089),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_13022),
.Y(n_13150)
);

INVx1_ASAP7_75t_L g13151 ( 
.A(n_12951),
.Y(n_13151)
);

INVx1_ASAP7_75t_L g13152 ( 
.A(n_13019),
.Y(n_13152)
);

AND2x2_ASAP7_75t_L g13153 ( 
.A(n_12975),
.B(n_2090),
.Y(n_13153)
);

AOI22xp33_ASAP7_75t_L g13154 ( 
.A1(n_13051),
.A2(n_2092),
.B1(n_2090),
.B2(n_2091),
.Y(n_13154)
);

AND2x2_ASAP7_75t_L g13155 ( 
.A(n_12993),
.B(n_2091),
.Y(n_13155)
);

INVx1_ASAP7_75t_L g13156 ( 
.A(n_13031),
.Y(n_13156)
);

NAND2xp5_ASAP7_75t_L g13157 ( 
.A(n_13028),
.B(n_2092),
.Y(n_13157)
);

INVx1_ASAP7_75t_L g13158 ( 
.A(n_13044),
.Y(n_13158)
);

OR2x2_ASAP7_75t_L g13159 ( 
.A(n_13016),
.B(n_2093),
.Y(n_13159)
);

NAND2xp5_ASAP7_75t_L g13160 ( 
.A(n_13040),
.B(n_2093),
.Y(n_13160)
);

AND2x2_ASAP7_75t_L g13161 ( 
.A(n_13024),
.B(n_2094),
.Y(n_13161)
);

INVx3_ASAP7_75t_L g13162 ( 
.A(n_13053),
.Y(n_13162)
);

NAND2xp5_ASAP7_75t_L g13163 ( 
.A(n_13027),
.B(n_2094),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_12981),
.B(n_2095),
.Y(n_13164)
);

NAND2xp5_ASAP7_75t_L g13165 ( 
.A(n_13042),
.B(n_2095),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_13035),
.Y(n_13166)
);

INVx2_ASAP7_75t_SL g13167 ( 
.A(n_13043),
.Y(n_13167)
);

OR2x2_ASAP7_75t_L g13168 ( 
.A(n_13046),
.B(n_2096),
.Y(n_13168)
);

INVx2_ASAP7_75t_L g13169 ( 
.A(n_13041),
.Y(n_13169)
);

AND2x2_ASAP7_75t_L g13170 ( 
.A(n_12972),
.B(n_2096),
.Y(n_13170)
);

INVxp67_ASAP7_75t_L g13171 ( 
.A(n_12955),
.Y(n_13171)
);

AND2x2_ASAP7_75t_L g13172 ( 
.A(n_12955),
.B(n_2097),
.Y(n_13172)
);

AND2x2_ASAP7_75t_L g13173 ( 
.A(n_12955),
.B(n_2097),
.Y(n_13173)
);

OR2x2_ASAP7_75t_L g13174 ( 
.A(n_12960),
.B(n_2098),
.Y(n_13174)
);

INVx2_ASAP7_75t_L g13175 ( 
.A(n_12960),
.Y(n_13175)
);

NAND2xp5_ASAP7_75t_L g13176 ( 
.A(n_12955),
.B(n_2098),
.Y(n_13176)
);

INVx1_ASAP7_75t_L g13177 ( 
.A(n_12960),
.Y(n_13177)
);

AND2x2_ASAP7_75t_L g13178 ( 
.A(n_12955),
.B(n_2099),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_12960),
.Y(n_13179)
);

AND2x2_ASAP7_75t_L g13180 ( 
.A(n_13128),
.B(n_2099),
.Y(n_13180)
);

INVx1_ASAP7_75t_L g13181 ( 
.A(n_13072),
.Y(n_13181)
);

OR2x2_ASAP7_75t_L g13182 ( 
.A(n_13059),
.B(n_2100),
.Y(n_13182)
);

NAND2xp5_ASAP7_75t_L g13183 ( 
.A(n_13060),
.B(n_2101),
.Y(n_13183)
);

INVx2_ASAP7_75t_L g13184 ( 
.A(n_13175),
.Y(n_13184)
);

INVx1_ASAP7_75t_L g13185 ( 
.A(n_13073),
.Y(n_13185)
);

INVx2_ASAP7_75t_L g13186 ( 
.A(n_13074),
.Y(n_13186)
);

HB1xp67_ASAP7_75t_L g13187 ( 
.A(n_13139),
.Y(n_13187)
);

INVx1_ASAP7_75t_L g13188 ( 
.A(n_13075),
.Y(n_13188)
);

AND2x2_ASAP7_75t_L g13189 ( 
.A(n_13132),
.B(n_2101),
.Y(n_13189)
);

INVx2_ASAP7_75t_L g13190 ( 
.A(n_13174),
.Y(n_13190)
);

AND2x2_ASAP7_75t_L g13191 ( 
.A(n_13082),
.B(n_2102),
.Y(n_13191)
);

AND2x2_ASAP7_75t_L g13192 ( 
.A(n_13177),
.B(n_2102),
.Y(n_13192)
);

BUFx3_ASAP7_75t_L g13193 ( 
.A(n_13065),
.Y(n_13193)
);

NOR3xp33_ASAP7_75t_L g13194 ( 
.A(n_13171),
.B(n_2103),
.C(n_2104),
.Y(n_13194)
);

AND2x2_ASAP7_75t_L g13195 ( 
.A(n_13179),
.B(n_2103),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_13136),
.Y(n_13196)
);

INVx1_ASAP7_75t_L g13197 ( 
.A(n_13172),
.Y(n_13197)
);

INVxp67_ASAP7_75t_SL g13198 ( 
.A(n_13162),
.Y(n_13198)
);

OR2x6_ASAP7_75t_L g13199 ( 
.A(n_13131),
.B(n_2105),
.Y(n_13199)
);

INVx2_ASAP7_75t_L g13200 ( 
.A(n_13173),
.Y(n_13200)
);

AND2x2_ASAP7_75t_L g13201 ( 
.A(n_13178),
.B(n_13170),
.Y(n_13201)
);

INVx2_ASAP7_75t_L g13202 ( 
.A(n_13094),
.Y(n_13202)
);

INVx2_ASAP7_75t_SL g13203 ( 
.A(n_13126),
.Y(n_13203)
);

AND2x2_ASAP7_75t_L g13204 ( 
.A(n_13056),
.B(n_2105),
.Y(n_13204)
);

AND2x2_ASAP7_75t_L g13205 ( 
.A(n_13145),
.B(n_2106),
.Y(n_13205)
);

NAND2xp67_ASAP7_75t_L g13206 ( 
.A(n_13153),
.B(n_2107),
.Y(n_13206)
);

AND2x2_ASAP7_75t_L g13207 ( 
.A(n_13098),
.B(n_2108),
.Y(n_13207)
);

AND2x2_ASAP7_75t_L g13208 ( 
.A(n_13096),
.B(n_2108),
.Y(n_13208)
);

NAND2xp5_ASAP7_75t_L g13209 ( 
.A(n_13087),
.B(n_2109),
.Y(n_13209)
);

NAND2xp5_ASAP7_75t_L g13210 ( 
.A(n_13138),
.B(n_2109),
.Y(n_13210)
);

INVx2_ASAP7_75t_L g13211 ( 
.A(n_13094),
.Y(n_13211)
);

INVx1_ASAP7_75t_L g13212 ( 
.A(n_13090),
.Y(n_13212)
);

INVx1_ASAP7_75t_SL g13213 ( 
.A(n_13140),
.Y(n_13213)
);

INVx1_ASAP7_75t_L g13214 ( 
.A(n_13076),
.Y(n_13214)
);

NAND2xp5_ASAP7_75t_L g13215 ( 
.A(n_13057),
.B(n_2110),
.Y(n_13215)
);

AND2x2_ASAP7_75t_L g13216 ( 
.A(n_13061),
.B(n_2110),
.Y(n_13216)
);

INVx1_ASAP7_75t_SL g13217 ( 
.A(n_13116),
.Y(n_13217)
);

NAND2xp5_ASAP7_75t_L g13218 ( 
.A(n_13064),
.B(n_2111),
.Y(n_13218)
);

INVx1_ASAP7_75t_L g13219 ( 
.A(n_13062),
.Y(n_13219)
);

INVxp67_ASAP7_75t_SL g13220 ( 
.A(n_13158),
.Y(n_13220)
);

INVx2_ASAP7_75t_L g13221 ( 
.A(n_13055),
.Y(n_13221)
);

NAND2x1p5_ASAP7_75t_L g13222 ( 
.A(n_13067),
.B(n_2112),
.Y(n_13222)
);

INVx2_ASAP7_75t_L g13223 ( 
.A(n_13071),
.Y(n_13223)
);

INVx1_ASAP7_75t_L g13224 ( 
.A(n_13121),
.Y(n_13224)
);

INVx1_ASAP7_75t_L g13225 ( 
.A(n_13068),
.Y(n_13225)
);

INVx2_ASAP7_75t_L g13226 ( 
.A(n_13085),
.Y(n_13226)
);

AND2x4_ASAP7_75t_L g13227 ( 
.A(n_13089),
.B(n_2112),
.Y(n_13227)
);

NOR2xp67_ASAP7_75t_SL g13228 ( 
.A(n_13066),
.B(n_2113),
.Y(n_13228)
);

NAND2xp5_ASAP7_75t_L g13229 ( 
.A(n_13150),
.B(n_2113),
.Y(n_13229)
);

OAI21xp33_ASAP7_75t_L g13230 ( 
.A1(n_13063),
.A2(n_2114),
.B(n_2115),
.Y(n_13230)
);

INVx1_ASAP7_75t_L g13231 ( 
.A(n_13102),
.Y(n_13231)
);

INVx1_ASAP7_75t_L g13232 ( 
.A(n_13084),
.Y(n_13232)
);

NAND2x1_ASAP7_75t_SL g13233 ( 
.A(n_13106),
.B(n_2114),
.Y(n_13233)
);

OR2x2_ASAP7_75t_L g13234 ( 
.A(n_13100),
.B(n_2116),
.Y(n_13234)
);

AND2x4_ASAP7_75t_SL g13235 ( 
.A(n_13093),
.B(n_2116),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_13144),
.Y(n_13236)
);

OR2x2_ASAP7_75t_L g13237 ( 
.A(n_13176),
.B(n_2117),
.Y(n_13237)
);

OR2x2_ASAP7_75t_L g13238 ( 
.A(n_13129),
.B(n_2117),
.Y(n_13238)
);

AND2x2_ASAP7_75t_L g13239 ( 
.A(n_13115),
.B(n_2118),
.Y(n_13239)
);

INVx1_ASAP7_75t_L g13240 ( 
.A(n_13105),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_13117),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_13120),
.Y(n_13242)
);

INVx1_ASAP7_75t_L g13243 ( 
.A(n_13141),
.Y(n_13243)
);

BUFx2_ASAP7_75t_L g13244 ( 
.A(n_13109),
.Y(n_13244)
);

INVx1_ASAP7_75t_L g13245 ( 
.A(n_13058),
.Y(n_13245)
);

OR2x2_ASAP7_75t_L g13246 ( 
.A(n_13103),
.B(n_2119),
.Y(n_13246)
);

INVxp67_ASAP7_75t_SL g13247 ( 
.A(n_13125),
.Y(n_13247)
);

NAND2x1_ASAP7_75t_L g13248 ( 
.A(n_13112),
.B(n_2119),
.Y(n_13248)
);

INVx1_ASAP7_75t_L g13249 ( 
.A(n_13088),
.Y(n_13249)
);

INVx1_ASAP7_75t_L g13250 ( 
.A(n_13113),
.Y(n_13250)
);

INVx1_ASAP7_75t_L g13251 ( 
.A(n_13122),
.Y(n_13251)
);

AND2x2_ASAP7_75t_L g13252 ( 
.A(n_13097),
.B(n_2120),
.Y(n_13252)
);

INVx2_ASAP7_75t_L g13253 ( 
.A(n_13081),
.Y(n_13253)
);

INVx1_ASAP7_75t_L g13254 ( 
.A(n_13123),
.Y(n_13254)
);

AND2x2_ASAP7_75t_L g13255 ( 
.A(n_13079),
.B(n_2121),
.Y(n_13255)
);

AND2x2_ASAP7_75t_L g13256 ( 
.A(n_13091),
.B(n_2122),
.Y(n_13256)
);

INVx2_ASAP7_75t_SL g13257 ( 
.A(n_13147),
.Y(n_13257)
);

AND2x2_ASAP7_75t_L g13258 ( 
.A(n_13092),
.B(n_2122),
.Y(n_13258)
);

OAI21xp33_ASAP7_75t_L g13259 ( 
.A1(n_13099),
.A2(n_13156),
.B(n_13118),
.Y(n_13259)
);

INVx1_ASAP7_75t_L g13260 ( 
.A(n_13124),
.Y(n_13260)
);

NAND2xp5_ASAP7_75t_L g13261 ( 
.A(n_13070),
.B(n_2123),
.Y(n_13261)
);

OR2x2_ASAP7_75t_L g13262 ( 
.A(n_13080),
.B(n_2124),
.Y(n_13262)
);

INVx2_ASAP7_75t_L g13263 ( 
.A(n_13146),
.Y(n_13263)
);

AOI211xp5_ASAP7_75t_SL g13264 ( 
.A1(n_13134),
.A2(n_2128),
.B(n_2124),
.C(n_2127),
.Y(n_13264)
);

AND2x2_ASAP7_75t_L g13265 ( 
.A(n_13101),
.B(n_2127),
.Y(n_13265)
);

OR2x2_ASAP7_75t_L g13266 ( 
.A(n_13078),
.B(n_2128),
.Y(n_13266)
);

NAND2xp5_ASAP7_75t_L g13267 ( 
.A(n_13133),
.B(n_13137),
.Y(n_13267)
);

INVx1_ASAP7_75t_L g13268 ( 
.A(n_13095),
.Y(n_13268)
);

INVx2_ASAP7_75t_L g13269 ( 
.A(n_13168),
.Y(n_13269)
);

NOR2xp33_ASAP7_75t_SL g13270 ( 
.A(n_13127),
.B(n_2129),
.Y(n_13270)
);

NAND2xp5_ASAP7_75t_L g13271 ( 
.A(n_13148),
.B(n_2129),
.Y(n_13271)
);

AND2x2_ASAP7_75t_L g13272 ( 
.A(n_13164),
.B(n_2130),
.Y(n_13272)
);

INVx1_ASAP7_75t_SL g13273 ( 
.A(n_13159),
.Y(n_13273)
);

NAND2xp5_ASAP7_75t_L g13274 ( 
.A(n_13108),
.B(n_2131),
.Y(n_13274)
);

CKINVDCx16_ASAP7_75t_R g13275 ( 
.A(n_13130),
.Y(n_13275)
);

AND2x2_ASAP7_75t_L g13276 ( 
.A(n_13110),
.B(n_2132),
.Y(n_13276)
);

NAND2xp5_ASAP7_75t_L g13277 ( 
.A(n_13069),
.B(n_2133),
.Y(n_13277)
);

INVx1_ASAP7_75t_L g13278 ( 
.A(n_13155),
.Y(n_13278)
);

AND2x2_ASAP7_75t_L g13279 ( 
.A(n_13114),
.B(n_2133),
.Y(n_13279)
);

INVx1_ASAP7_75t_L g13280 ( 
.A(n_13149),
.Y(n_13280)
);

AND2x4_ASAP7_75t_SL g13281 ( 
.A(n_13142),
.B(n_2134),
.Y(n_13281)
);

INVx1_ASAP7_75t_SL g13282 ( 
.A(n_13161),
.Y(n_13282)
);

OR2x2_ASAP7_75t_L g13283 ( 
.A(n_13111),
.B(n_2134),
.Y(n_13283)
);

INVx2_ASAP7_75t_SL g13284 ( 
.A(n_13167),
.Y(n_13284)
);

OAI21xp33_ASAP7_75t_L g13285 ( 
.A1(n_13083),
.A2(n_13086),
.B(n_13135),
.Y(n_13285)
);

AOI21xp33_ASAP7_75t_L g13286 ( 
.A1(n_13143),
.A2(n_2135),
.B(n_2136),
.Y(n_13286)
);

INVx1_ASAP7_75t_SL g13287 ( 
.A(n_13119),
.Y(n_13287)
);

INVx1_ASAP7_75t_L g13288 ( 
.A(n_13077),
.Y(n_13288)
);

INVx1_ASAP7_75t_L g13289 ( 
.A(n_13104),
.Y(n_13289)
);

INVx2_ASAP7_75t_L g13290 ( 
.A(n_13169),
.Y(n_13290)
);

NOR2x1p5_ASAP7_75t_L g13291 ( 
.A(n_13107),
.B(n_2135),
.Y(n_13291)
);

OR2x2_ASAP7_75t_L g13292 ( 
.A(n_13160),
.B(n_2136),
.Y(n_13292)
);

NAND2xp5_ASAP7_75t_L g13293 ( 
.A(n_13151),
.B(n_2137),
.Y(n_13293)
);

INVx1_ASAP7_75t_L g13294 ( 
.A(n_13165),
.Y(n_13294)
);

INVx2_ASAP7_75t_L g13295 ( 
.A(n_13152),
.Y(n_13295)
);

INVx1_ASAP7_75t_L g13296 ( 
.A(n_13157),
.Y(n_13296)
);

INVx4_ASAP7_75t_L g13297 ( 
.A(n_13166),
.Y(n_13297)
);

INVx1_ASAP7_75t_L g13298 ( 
.A(n_13163),
.Y(n_13298)
);

INVx1_ASAP7_75t_L g13299 ( 
.A(n_13154),
.Y(n_13299)
);

INVx1_ASAP7_75t_L g13300 ( 
.A(n_13072),
.Y(n_13300)
);

AND2x2_ASAP7_75t_L g13301 ( 
.A(n_13128),
.B(n_2137),
.Y(n_13301)
);

HB1xp67_ASAP7_75t_L g13302 ( 
.A(n_13139),
.Y(n_13302)
);

AND2x2_ASAP7_75t_L g13303 ( 
.A(n_13128),
.B(n_2138),
.Y(n_13303)
);

NAND2xp5_ASAP7_75t_L g13304 ( 
.A(n_13059),
.B(n_2138),
.Y(n_13304)
);

INVx1_ASAP7_75t_L g13305 ( 
.A(n_13072),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_13072),
.Y(n_13306)
);

INVx2_ASAP7_75t_L g13307 ( 
.A(n_13059),
.Y(n_13307)
);

NAND2xp5_ASAP7_75t_L g13308 ( 
.A(n_13059),
.B(n_2139),
.Y(n_13308)
);

AND2x2_ASAP7_75t_L g13309 ( 
.A(n_13128),
.B(n_2139),
.Y(n_13309)
);

OAI32xp33_ASAP7_75t_L g13310 ( 
.A1(n_13150),
.A2(n_2142),
.A3(n_2140),
.B1(n_2141),
.B2(n_2143),
.Y(n_13310)
);

INVx1_ASAP7_75t_L g13311 ( 
.A(n_13072),
.Y(n_13311)
);

NAND2xp5_ASAP7_75t_L g13312 ( 
.A(n_13059),
.B(n_2140),
.Y(n_13312)
);

INVx1_ASAP7_75t_L g13313 ( 
.A(n_13072),
.Y(n_13313)
);

NOR3x1_ASAP7_75t_L g13314 ( 
.A(n_13128),
.B(n_2141),
.C(n_2143),
.Y(n_13314)
);

OR2x2_ASAP7_75t_L g13315 ( 
.A(n_13059),
.B(n_2144),
.Y(n_13315)
);

AND2x2_ASAP7_75t_L g13316 ( 
.A(n_13128),
.B(n_2145),
.Y(n_13316)
);

AND2x2_ASAP7_75t_L g13317 ( 
.A(n_13128),
.B(n_2145),
.Y(n_13317)
);

INVx2_ASAP7_75t_L g13318 ( 
.A(n_13059),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_13072),
.Y(n_13319)
);

INVx2_ASAP7_75t_L g13320 ( 
.A(n_13059),
.Y(n_13320)
);

INVx1_ASAP7_75t_L g13321 ( 
.A(n_13072),
.Y(n_13321)
);

AND2x4_ASAP7_75t_L g13322 ( 
.A(n_13175),
.B(n_2147),
.Y(n_13322)
);

INVx1_ASAP7_75t_L g13323 ( 
.A(n_13072),
.Y(n_13323)
);

AND2x2_ASAP7_75t_L g13324 ( 
.A(n_13128),
.B(n_2149),
.Y(n_13324)
);

AND2x4_ASAP7_75t_L g13325 ( 
.A(n_13175),
.B(n_2149),
.Y(n_13325)
);

NOR2xp33_ASAP7_75t_L g13326 ( 
.A(n_13098),
.B(n_2150),
.Y(n_13326)
);

NAND2xp5_ASAP7_75t_L g13327 ( 
.A(n_13059),
.B(n_2151),
.Y(n_13327)
);

NAND2xp5_ASAP7_75t_L g13328 ( 
.A(n_13059),
.B(n_2151),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_13072),
.Y(n_13329)
);

INVx1_ASAP7_75t_L g13330 ( 
.A(n_13072),
.Y(n_13330)
);

NAND2xp33_ASAP7_75t_SL g13331 ( 
.A(n_13233),
.B(n_2152),
.Y(n_13331)
);

INVx1_ASAP7_75t_L g13332 ( 
.A(n_13187),
.Y(n_13332)
);

INVx2_ASAP7_75t_L g13333 ( 
.A(n_13193),
.Y(n_13333)
);

INVx1_ASAP7_75t_L g13334 ( 
.A(n_13302),
.Y(n_13334)
);

AND2x2_ASAP7_75t_L g13335 ( 
.A(n_13201),
.B(n_2152),
.Y(n_13335)
);

INVx2_ASAP7_75t_L g13336 ( 
.A(n_13222),
.Y(n_13336)
);

AND2x2_ASAP7_75t_L g13337 ( 
.A(n_13180),
.B(n_2153),
.Y(n_13337)
);

AOI22xp5_ASAP7_75t_L g13338 ( 
.A1(n_13184),
.A2(n_2155),
.B1(n_2153),
.B2(n_2154),
.Y(n_13338)
);

AND2x2_ASAP7_75t_L g13339 ( 
.A(n_13301),
.B(n_2154),
.Y(n_13339)
);

AND2x2_ASAP7_75t_L g13340 ( 
.A(n_13303),
.B(n_2155),
.Y(n_13340)
);

INVx2_ASAP7_75t_L g13341 ( 
.A(n_13199),
.Y(n_13341)
);

INVx2_ASAP7_75t_SL g13342 ( 
.A(n_13235),
.Y(n_13342)
);

OR2x2_ASAP7_75t_L g13343 ( 
.A(n_13217),
.B(n_13223),
.Y(n_13343)
);

NAND2xp5_ASAP7_75t_L g13344 ( 
.A(n_13219),
.B(n_2156),
.Y(n_13344)
);

AND2x2_ASAP7_75t_L g13345 ( 
.A(n_13309),
.B(n_2156),
.Y(n_13345)
);

AND2x4_ASAP7_75t_L g13346 ( 
.A(n_13203),
.B(n_2157),
.Y(n_13346)
);

NAND2xp5_ASAP7_75t_L g13347 ( 
.A(n_13225),
.B(n_2157),
.Y(n_13347)
);

AOI21xp33_ASAP7_75t_SL g13348 ( 
.A1(n_13275),
.A2(n_2158),
.B(n_2159),
.Y(n_13348)
);

NAND2xp5_ASAP7_75t_L g13349 ( 
.A(n_13212),
.B(n_2158),
.Y(n_13349)
);

NAND2xp5_ASAP7_75t_L g13350 ( 
.A(n_13316),
.B(n_2159),
.Y(n_13350)
);

INVx1_ASAP7_75t_L g13351 ( 
.A(n_13317),
.Y(n_13351)
);

INVx1_ASAP7_75t_L g13352 ( 
.A(n_13324),
.Y(n_13352)
);

AND2x2_ASAP7_75t_L g13353 ( 
.A(n_13205),
.B(n_2160),
.Y(n_13353)
);

AND2x2_ASAP7_75t_L g13354 ( 
.A(n_13221),
.B(n_2160),
.Y(n_13354)
);

INVx2_ASAP7_75t_L g13355 ( 
.A(n_13199),
.Y(n_13355)
);

INVx1_ASAP7_75t_L g13356 ( 
.A(n_13206),
.Y(n_13356)
);

NAND2xp5_ASAP7_75t_L g13357 ( 
.A(n_13198),
.B(n_2161),
.Y(n_13357)
);

INVx2_ASAP7_75t_L g13358 ( 
.A(n_13207),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_13186),
.B(n_2161),
.Y(n_13359)
);

INVx2_ASAP7_75t_L g13360 ( 
.A(n_13189),
.Y(n_13360)
);

AOI222xp33_ASAP7_75t_L g13361 ( 
.A1(n_13196),
.A2(n_2164),
.B1(n_2167),
.B2(n_2162),
.C1(n_2163),
.C2(n_2166),
.Y(n_13361)
);

NAND2xp5_ASAP7_75t_L g13362 ( 
.A(n_13220),
.B(n_2162),
.Y(n_13362)
);

INVx1_ASAP7_75t_L g13363 ( 
.A(n_13216),
.Y(n_13363)
);

NAND2xp5_ASAP7_75t_L g13364 ( 
.A(n_13214),
.B(n_13191),
.Y(n_13364)
);

AND2x4_ASAP7_75t_L g13365 ( 
.A(n_13307),
.B(n_2168),
.Y(n_13365)
);

AND2x2_ASAP7_75t_L g13366 ( 
.A(n_13200),
.B(n_2168),
.Y(n_13366)
);

INVx2_ASAP7_75t_L g13367 ( 
.A(n_13239),
.Y(n_13367)
);

INVx3_ASAP7_75t_L g13368 ( 
.A(n_13297),
.Y(n_13368)
);

INVx1_ASAP7_75t_L g13369 ( 
.A(n_13210),
.Y(n_13369)
);

NAND2x1p5_ASAP7_75t_L g13370 ( 
.A(n_13314),
.B(n_2169),
.Y(n_13370)
);

NAND2x2_ASAP7_75t_L g13371 ( 
.A(n_13257),
.B(n_2169),
.Y(n_13371)
);

INVx1_ASAP7_75t_L g13372 ( 
.A(n_13208),
.Y(n_13372)
);

INVx1_ASAP7_75t_L g13373 ( 
.A(n_13248),
.Y(n_13373)
);

OR2x2_ASAP7_75t_L g13374 ( 
.A(n_13213),
.B(n_2170),
.Y(n_13374)
);

INVx1_ASAP7_75t_SL g13375 ( 
.A(n_13234),
.Y(n_13375)
);

NAND3x2_ASAP7_75t_L g13376 ( 
.A(n_13244),
.B(n_2171),
.C(n_2173),
.Y(n_13376)
);

NAND2xp5_ASAP7_75t_L g13377 ( 
.A(n_13318),
.B(n_2171),
.Y(n_13377)
);

NAND2xp5_ASAP7_75t_L g13378 ( 
.A(n_13320),
.B(n_2173),
.Y(n_13378)
);

AND2x2_ASAP7_75t_L g13379 ( 
.A(n_13197),
.B(n_2174),
.Y(n_13379)
);

INVxp67_ASAP7_75t_L g13380 ( 
.A(n_13270),
.Y(n_13380)
);

NAND2xp5_ASAP7_75t_L g13381 ( 
.A(n_13322),
.B(n_13325),
.Y(n_13381)
);

INVx1_ASAP7_75t_L g13382 ( 
.A(n_13228),
.Y(n_13382)
);

INVx1_ASAP7_75t_L g13383 ( 
.A(n_13182),
.Y(n_13383)
);

NAND2xp5_ASAP7_75t_L g13384 ( 
.A(n_13264),
.B(n_2174),
.Y(n_13384)
);

INVx1_ASAP7_75t_L g13385 ( 
.A(n_13315),
.Y(n_13385)
);

INVx1_ASAP7_75t_L g13386 ( 
.A(n_13204),
.Y(n_13386)
);

AND2x4_ASAP7_75t_SL g13387 ( 
.A(n_13253),
.B(n_13202),
.Y(n_13387)
);

AND2x2_ASAP7_75t_L g13388 ( 
.A(n_13247),
.B(n_2175),
.Y(n_13388)
);

INVx1_ASAP7_75t_L g13389 ( 
.A(n_13252),
.Y(n_13389)
);

INVx2_ASAP7_75t_L g13390 ( 
.A(n_13211),
.Y(n_13390)
);

NAND2xp5_ASAP7_75t_L g13391 ( 
.A(n_13281),
.B(n_2175),
.Y(n_13391)
);

OR2x2_ASAP7_75t_L g13392 ( 
.A(n_13209),
.B(n_2176),
.Y(n_13392)
);

INVx1_ASAP7_75t_L g13393 ( 
.A(n_13255),
.Y(n_13393)
);

INVxp67_ASAP7_75t_SL g13394 ( 
.A(n_13291),
.Y(n_13394)
);

AND2x2_ASAP7_75t_L g13395 ( 
.A(n_13231),
.B(n_2176),
.Y(n_13395)
);

AND2x4_ASAP7_75t_L g13396 ( 
.A(n_13284),
.B(n_2177),
.Y(n_13396)
);

OR2x2_ASAP7_75t_L g13397 ( 
.A(n_13246),
.B(n_2178),
.Y(n_13397)
);

INVx1_ASAP7_75t_L g13398 ( 
.A(n_13256),
.Y(n_13398)
);

AND2x2_ASAP7_75t_L g13399 ( 
.A(n_13243),
.B(n_2178),
.Y(n_13399)
);

HB1xp67_ASAP7_75t_L g13400 ( 
.A(n_13181),
.Y(n_13400)
);

INVx1_ASAP7_75t_L g13401 ( 
.A(n_13258),
.Y(n_13401)
);

AND2x2_ASAP7_75t_L g13402 ( 
.A(n_13226),
.B(n_2179),
.Y(n_13402)
);

AND2x2_ASAP7_75t_L g13403 ( 
.A(n_13224),
.B(n_2179),
.Y(n_13403)
);

INVxp67_ASAP7_75t_SL g13404 ( 
.A(n_13326),
.Y(n_13404)
);

INVx1_ASAP7_75t_SL g13405 ( 
.A(n_13262),
.Y(n_13405)
);

AND2x4_ASAP7_75t_L g13406 ( 
.A(n_13190),
.B(n_2180),
.Y(n_13406)
);

AND2x4_ASAP7_75t_L g13407 ( 
.A(n_13240),
.B(n_2180),
.Y(n_13407)
);

OR2x2_ASAP7_75t_L g13408 ( 
.A(n_13183),
.B(n_2181),
.Y(n_13408)
);

AOI21xp5_ASAP7_75t_SL g13409 ( 
.A1(n_13300),
.A2(n_2181),
.B(n_2182),
.Y(n_13409)
);

NAND2xp5_ASAP7_75t_SL g13410 ( 
.A(n_13263),
.B(n_2182),
.Y(n_13410)
);

NOR2xp67_ASAP7_75t_SL g13411 ( 
.A(n_13266),
.B(n_2184),
.Y(n_13411)
);

AND3x1_ASAP7_75t_L g13412 ( 
.A(n_13259),
.B(n_2185),
.C(n_2186),
.Y(n_13412)
);

INVx1_ASAP7_75t_L g13413 ( 
.A(n_13192),
.Y(n_13413)
);

AND2x2_ASAP7_75t_L g13414 ( 
.A(n_13241),
.B(n_2186),
.Y(n_13414)
);

AND2x2_ASAP7_75t_L g13415 ( 
.A(n_13242),
.B(n_2187),
.Y(n_13415)
);

OR2x2_ASAP7_75t_L g13416 ( 
.A(n_13304),
.B(n_2187),
.Y(n_13416)
);

AND2x2_ASAP7_75t_L g13417 ( 
.A(n_13249),
.B(n_2188),
.Y(n_13417)
);

NAND2xp5_ASAP7_75t_L g13418 ( 
.A(n_13195),
.B(n_2188),
.Y(n_13418)
);

INVx2_ASAP7_75t_L g13419 ( 
.A(n_13227),
.Y(n_13419)
);

HB1xp67_ASAP7_75t_L g13420 ( 
.A(n_13305),
.Y(n_13420)
);

INVxp33_ASAP7_75t_L g13421 ( 
.A(n_13267),
.Y(n_13421)
);

AOI21xp33_ASAP7_75t_L g13422 ( 
.A1(n_13306),
.A2(n_2189),
.B(n_2190),
.Y(n_13422)
);

NAND2xp5_ASAP7_75t_L g13423 ( 
.A(n_13265),
.B(n_2191),
.Y(n_13423)
);

NAND2xp5_ASAP7_75t_L g13424 ( 
.A(n_13276),
.B(n_2191),
.Y(n_13424)
);

OAI211xp5_ASAP7_75t_L g13425 ( 
.A1(n_13285),
.A2(n_2194),
.B(n_2192),
.C(n_2193),
.Y(n_13425)
);

AND2x2_ASAP7_75t_L g13426 ( 
.A(n_13272),
.B(n_2192),
.Y(n_13426)
);

INVxp67_ASAP7_75t_L g13427 ( 
.A(n_13238),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_13308),
.Y(n_13428)
);

INVx1_ASAP7_75t_L g13429 ( 
.A(n_13312),
.Y(n_13429)
);

NAND2x1_ASAP7_75t_L g13430 ( 
.A(n_13311),
.B(n_2193),
.Y(n_13430)
);

INVx2_ASAP7_75t_L g13431 ( 
.A(n_13237),
.Y(n_13431)
);

INVx1_ASAP7_75t_L g13432 ( 
.A(n_13327),
.Y(n_13432)
);

OR2x2_ASAP7_75t_L g13433 ( 
.A(n_13328),
.B(n_2194),
.Y(n_13433)
);

OR2x2_ASAP7_75t_L g13434 ( 
.A(n_13282),
.B(n_2195),
.Y(n_13434)
);

AND2x4_ASAP7_75t_L g13435 ( 
.A(n_13232),
.B(n_2195),
.Y(n_13435)
);

AND2x2_ASAP7_75t_L g13436 ( 
.A(n_13185),
.B(n_2196),
.Y(n_13436)
);

NOR2xp33_ASAP7_75t_L g13437 ( 
.A(n_13230),
.B(n_2196),
.Y(n_13437)
);

HB1xp67_ASAP7_75t_L g13438 ( 
.A(n_13313),
.Y(n_13438)
);

INVx1_ASAP7_75t_SL g13439 ( 
.A(n_13279),
.Y(n_13439)
);

INVx1_ASAP7_75t_L g13440 ( 
.A(n_13319),
.Y(n_13440)
);

INVx1_ASAP7_75t_L g13441 ( 
.A(n_13321),
.Y(n_13441)
);

OR2x2_ASAP7_75t_L g13442 ( 
.A(n_13218),
.B(n_2197),
.Y(n_13442)
);

INVx1_ASAP7_75t_L g13443 ( 
.A(n_13323),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_13188),
.B(n_2197),
.Y(n_13444)
);

AND2x2_ASAP7_75t_L g13445 ( 
.A(n_13278),
.B(n_13251),
.Y(n_13445)
);

OR2x2_ASAP7_75t_L g13446 ( 
.A(n_13215),
.B(n_2198),
.Y(n_13446)
);

INVx1_ASAP7_75t_L g13447 ( 
.A(n_13329),
.Y(n_13447)
);

NAND2xp5_ASAP7_75t_L g13448 ( 
.A(n_13254),
.B(n_2199),
.Y(n_13448)
);

OR2x2_ASAP7_75t_L g13449 ( 
.A(n_13274),
.B(n_2199),
.Y(n_13449)
);

AND2x2_ASAP7_75t_L g13450 ( 
.A(n_13260),
.B(n_13269),
.Y(n_13450)
);

INVx1_ASAP7_75t_L g13451 ( 
.A(n_13330),
.Y(n_13451)
);

INVx1_ASAP7_75t_SL g13452 ( 
.A(n_13292),
.Y(n_13452)
);

AND2x2_ASAP7_75t_L g13453 ( 
.A(n_13273),
.B(n_2200),
.Y(n_13453)
);

AOI22xp33_ASAP7_75t_SL g13454 ( 
.A1(n_13245),
.A2(n_2202),
.B1(n_2200),
.B2(n_2201),
.Y(n_13454)
);

OR2x2_ASAP7_75t_L g13455 ( 
.A(n_13271),
.B(n_2202),
.Y(n_13455)
);

OR2x2_ASAP7_75t_L g13456 ( 
.A(n_13250),
.B(n_2203),
.Y(n_13456)
);

NAND2x1p5_ASAP7_75t_L g13457 ( 
.A(n_13290),
.B(n_2203),
.Y(n_13457)
);

OR2x2_ASAP7_75t_L g13458 ( 
.A(n_13229),
.B(n_2204),
.Y(n_13458)
);

INVx1_ASAP7_75t_SL g13459 ( 
.A(n_13283),
.Y(n_13459)
);

AND2x2_ASAP7_75t_SL g13460 ( 
.A(n_13194),
.B(n_2204),
.Y(n_13460)
);

AND2x2_ASAP7_75t_L g13461 ( 
.A(n_13299),
.B(n_2205),
.Y(n_13461)
);

INVx1_ASAP7_75t_L g13462 ( 
.A(n_13261),
.Y(n_13462)
);

INVx1_ASAP7_75t_L g13463 ( 
.A(n_13277),
.Y(n_13463)
);

BUFx2_ASAP7_75t_L g13464 ( 
.A(n_13295),
.Y(n_13464)
);

AND2x2_ASAP7_75t_L g13465 ( 
.A(n_13236),
.B(n_2206),
.Y(n_13465)
);

AND2x4_ASAP7_75t_L g13466 ( 
.A(n_13268),
.B(n_2206),
.Y(n_13466)
);

INVx1_ASAP7_75t_L g13467 ( 
.A(n_13293),
.Y(n_13467)
);

NOR2x2_ASAP7_75t_L g13468 ( 
.A(n_13287),
.B(n_2207),
.Y(n_13468)
);

AOI22xp5_ASAP7_75t_L g13469 ( 
.A1(n_13280),
.A2(n_2210),
.B1(n_2208),
.B2(n_2209),
.Y(n_13469)
);

INVx1_ASAP7_75t_L g13470 ( 
.A(n_13310),
.Y(n_13470)
);

AOI221xp5_ASAP7_75t_L g13471 ( 
.A1(n_13288),
.A2(n_2211),
.B1(n_2209),
.B2(n_2210),
.C(n_2212),
.Y(n_13471)
);

NAND2xp5_ASAP7_75t_L g13472 ( 
.A(n_13296),
.B(n_2211),
.Y(n_13472)
);

OA21x2_ASAP7_75t_L g13473 ( 
.A1(n_13286),
.A2(n_2212),
.B(n_2213),
.Y(n_13473)
);

OAI322xp33_ASAP7_75t_L g13474 ( 
.A1(n_13343),
.A2(n_13289),
.A3(n_13294),
.B1(n_13298),
.B2(n_2215),
.C1(n_2218),
.C2(n_2217),
.Y(n_13474)
);

OR2x2_ASAP7_75t_L g13475 ( 
.A(n_13370),
.B(n_2213),
.Y(n_13475)
);

INVx1_ASAP7_75t_L g13476 ( 
.A(n_13430),
.Y(n_13476)
);

OAI22xp5_ASAP7_75t_L g13477 ( 
.A1(n_13371),
.A2(n_2216),
.B1(n_2214),
.B2(n_2215),
.Y(n_13477)
);

OAI21xp33_ASAP7_75t_L g13478 ( 
.A1(n_13421),
.A2(n_2214),
.B(n_2216),
.Y(n_13478)
);

OAI21xp33_ASAP7_75t_L g13479 ( 
.A1(n_13387),
.A2(n_2218),
.B(n_2219),
.Y(n_13479)
);

INVxp67_ASAP7_75t_SL g13480 ( 
.A(n_13457),
.Y(n_13480)
);

INVx1_ASAP7_75t_L g13481 ( 
.A(n_13337),
.Y(n_13481)
);

INVxp67_ASAP7_75t_L g13482 ( 
.A(n_13331),
.Y(n_13482)
);

NAND2xp5_ASAP7_75t_L g13483 ( 
.A(n_13346),
.B(n_2219),
.Y(n_13483)
);

INVx1_ASAP7_75t_L g13484 ( 
.A(n_13339),
.Y(n_13484)
);

O2A1O1Ixp5_ASAP7_75t_SL g13485 ( 
.A1(n_13368),
.A2(n_2222),
.B(n_2220),
.C(n_2221),
.Y(n_13485)
);

INVx1_ASAP7_75t_SL g13486 ( 
.A(n_13468),
.Y(n_13486)
);

NAND2xp5_ASAP7_75t_L g13487 ( 
.A(n_13340),
.B(n_2220),
.Y(n_13487)
);

INVx2_ASAP7_75t_L g13488 ( 
.A(n_13345),
.Y(n_13488)
);

NAND2xp5_ASAP7_75t_L g13489 ( 
.A(n_13396),
.B(n_2221),
.Y(n_13489)
);

INVx1_ASAP7_75t_L g13490 ( 
.A(n_13353),
.Y(n_13490)
);

NAND2xp5_ASAP7_75t_L g13491 ( 
.A(n_13342),
.B(n_2222),
.Y(n_13491)
);

NAND2xp5_ASAP7_75t_L g13492 ( 
.A(n_13373),
.B(n_2223),
.Y(n_13492)
);

INVx1_ASAP7_75t_L g13493 ( 
.A(n_13335),
.Y(n_13493)
);

NAND2xp5_ASAP7_75t_L g13494 ( 
.A(n_13365),
.B(n_2224),
.Y(n_13494)
);

INVx1_ASAP7_75t_L g13495 ( 
.A(n_13400),
.Y(n_13495)
);

INVx1_ASAP7_75t_L g13496 ( 
.A(n_13420),
.Y(n_13496)
);

NOR2x1p5_ASAP7_75t_L g13497 ( 
.A(n_13394),
.B(n_2224),
.Y(n_13497)
);

INVx2_ASAP7_75t_SL g13498 ( 
.A(n_13341),
.Y(n_13498)
);

INVx1_ASAP7_75t_SL g13499 ( 
.A(n_13426),
.Y(n_13499)
);

INVx1_ASAP7_75t_SL g13500 ( 
.A(n_13434),
.Y(n_13500)
);

OR2x2_ASAP7_75t_L g13501 ( 
.A(n_13355),
.B(n_13384),
.Y(n_13501)
);

AND2x2_ASAP7_75t_L g13502 ( 
.A(n_13358),
.B(n_2225),
.Y(n_13502)
);

INVx1_ASAP7_75t_L g13503 ( 
.A(n_13438),
.Y(n_13503)
);

AOI22xp33_ASAP7_75t_L g13504 ( 
.A1(n_13333),
.A2(n_2228),
.B1(n_2226),
.B2(n_2227),
.Y(n_13504)
);

INVx2_ASAP7_75t_L g13505 ( 
.A(n_13397),
.Y(n_13505)
);

AOI21xp5_ASAP7_75t_L g13506 ( 
.A1(n_13381),
.A2(n_2226),
.B(n_2227),
.Y(n_13506)
);

AOI22xp5_ASAP7_75t_L g13507 ( 
.A1(n_13470),
.A2(n_2230),
.B1(n_2228),
.B2(n_2229),
.Y(n_13507)
);

AND2x2_ASAP7_75t_L g13508 ( 
.A(n_13336),
.B(n_2229),
.Y(n_13508)
);

INVx2_ASAP7_75t_L g13509 ( 
.A(n_13407),
.Y(n_13509)
);

AND2x2_ASAP7_75t_L g13510 ( 
.A(n_13388),
.B(n_2230),
.Y(n_13510)
);

NAND3xp33_ASAP7_75t_L g13511 ( 
.A(n_13412),
.B(n_2231),
.C(n_2232),
.Y(n_13511)
);

NAND2xp5_ASAP7_75t_L g13512 ( 
.A(n_13406),
.B(n_2231),
.Y(n_13512)
);

NOR3xp33_ASAP7_75t_L g13513 ( 
.A(n_13332),
.B(n_2233),
.C(n_2234),
.Y(n_13513)
);

OAI21xp33_ASAP7_75t_L g13514 ( 
.A1(n_13390),
.A2(n_2235),
.B(n_2237),
.Y(n_13514)
);

NOR3xp33_ASAP7_75t_L g13515 ( 
.A(n_13334),
.B(n_2235),
.C(n_2237),
.Y(n_13515)
);

INVxp67_ASAP7_75t_L g13516 ( 
.A(n_13411),
.Y(n_13516)
);

NAND2xp5_ASAP7_75t_L g13517 ( 
.A(n_13351),
.B(n_2238),
.Y(n_13517)
);

INVx1_ASAP7_75t_L g13518 ( 
.A(n_13354),
.Y(n_13518)
);

HB1xp67_ASAP7_75t_L g13519 ( 
.A(n_13473),
.Y(n_13519)
);

INVx2_ASAP7_75t_L g13520 ( 
.A(n_13456),
.Y(n_13520)
);

AOI32xp33_ASAP7_75t_L g13521 ( 
.A1(n_13461),
.A2(n_2240),
.A3(n_2238),
.B1(n_2239),
.B2(n_2241),
.Y(n_13521)
);

OR2x2_ASAP7_75t_L g13522 ( 
.A(n_13376),
.B(n_2239),
.Y(n_13522)
);

INVx1_ASAP7_75t_L g13523 ( 
.A(n_13379),
.Y(n_13523)
);

NAND3xp33_ASAP7_75t_L g13524 ( 
.A(n_13409),
.B(n_2241),
.C(n_2242),
.Y(n_13524)
);

OAI211xp5_ASAP7_75t_SL g13525 ( 
.A1(n_13380),
.A2(n_2244),
.B(n_2242),
.C(n_2243),
.Y(n_13525)
);

AND2x2_ASAP7_75t_L g13526 ( 
.A(n_13360),
.B(n_2243),
.Y(n_13526)
);

O2A1O1Ixp33_ASAP7_75t_L g13527 ( 
.A1(n_13362),
.A2(n_2246),
.B(n_2244),
.C(n_2245),
.Y(n_13527)
);

AND2x2_ASAP7_75t_L g13528 ( 
.A(n_13352),
.B(n_2245),
.Y(n_13528)
);

HB1xp67_ASAP7_75t_L g13529 ( 
.A(n_13356),
.Y(n_13529)
);

AOI21xp5_ASAP7_75t_L g13530 ( 
.A1(n_13410),
.A2(n_2247),
.B(n_2248),
.Y(n_13530)
);

AOI21xp5_ASAP7_75t_L g13531 ( 
.A1(n_13364),
.A2(n_2247),
.B(n_2248),
.Y(n_13531)
);

NAND2xp5_ASAP7_75t_L g13532 ( 
.A(n_13348),
.B(n_2249),
.Y(n_13532)
);

NAND2xp5_ASAP7_75t_L g13533 ( 
.A(n_13454),
.B(n_2249),
.Y(n_13533)
);

INVx1_ASAP7_75t_L g13534 ( 
.A(n_13399),
.Y(n_13534)
);

INVx1_ASAP7_75t_L g13535 ( 
.A(n_13350),
.Y(n_13535)
);

AOI32xp33_ASAP7_75t_L g13536 ( 
.A1(n_13450),
.A2(n_2253),
.A3(n_2251),
.B1(n_2252),
.B2(n_2254),
.Y(n_13536)
);

NAND2xp33_ASAP7_75t_SL g13537 ( 
.A(n_13382),
.B(n_2251),
.Y(n_13537)
);

AOI22xp5_ASAP7_75t_L g13538 ( 
.A1(n_13445),
.A2(n_2255),
.B1(n_2252),
.B2(n_2254),
.Y(n_13538)
);

AND2x2_ASAP7_75t_L g13539 ( 
.A(n_13367),
.B(n_2255),
.Y(n_13539)
);

INVx3_ASAP7_75t_L g13540 ( 
.A(n_13435),
.Y(n_13540)
);

INVx1_ASAP7_75t_L g13541 ( 
.A(n_13403),
.Y(n_13541)
);

INVx1_ASAP7_75t_L g13542 ( 
.A(n_13414),
.Y(n_13542)
);

INVx2_ASAP7_75t_L g13543 ( 
.A(n_13374),
.Y(n_13543)
);

NOR2xp33_ASAP7_75t_L g13544 ( 
.A(n_13363),
.B(n_2256),
.Y(n_13544)
);

OR2x2_ASAP7_75t_L g13545 ( 
.A(n_13344),
.B(n_2256),
.Y(n_13545)
);

OAI21xp5_ASAP7_75t_L g13546 ( 
.A1(n_13427),
.A2(n_13453),
.B(n_13347),
.Y(n_13546)
);

NAND2xp5_ASAP7_75t_L g13547 ( 
.A(n_13415),
.B(n_2257),
.Y(n_13547)
);

INVx1_ASAP7_75t_L g13548 ( 
.A(n_13417),
.Y(n_13548)
);

INVxp67_ASAP7_75t_L g13549 ( 
.A(n_13391),
.Y(n_13549)
);

AOI22xp33_ASAP7_75t_L g13550 ( 
.A1(n_13464),
.A2(n_2259),
.B1(n_2257),
.B2(n_2258),
.Y(n_13550)
);

NOR2xp33_ASAP7_75t_L g13551 ( 
.A(n_13372),
.B(n_2259),
.Y(n_13551)
);

OR2x2_ASAP7_75t_L g13552 ( 
.A(n_13377),
.B(n_2260),
.Y(n_13552)
);

NAND2x1_ASAP7_75t_L g13553 ( 
.A(n_13402),
.B(n_2260),
.Y(n_13553)
);

INVx3_ASAP7_75t_L g13554 ( 
.A(n_13466),
.Y(n_13554)
);

INVx1_ASAP7_75t_L g13555 ( 
.A(n_13395),
.Y(n_13555)
);

NAND2xp5_ASAP7_75t_L g13556 ( 
.A(n_13359),
.B(n_13366),
.Y(n_13556)
);

O2A1O1Ixp33_ASAP7_75t_L g13557 ( 
.A1(n_13349),
.A2(n_2263),
.B(n_2261),
.C(n_2262),
.Y(n_13557)
);

INVx2_ASAP7_75t_SL g13558 ( 
.A(n_13419),
.Y(n_13558)
);

INVx1_ASAP7_75t_L g13559 ( 
.A(n_13418),
.Y(n_13559)
);

NAND2xp5_ASAP7_75t_L g13560 ( 
.A(n_13375),
.B(n_2261),
.Y(n_13560)
);

INVx1_ASAP7_75t_L g13561 ( 
.A(n_13357),
.Y(n_13561)
);

INVx1_ASAP7_75t_L g13562 ( 
.A(n_13423),
.Y(n_13562)
);

INVx1_ASAP7_75t_L g13563 ( 
.A(n_13424),
.Y(n_13563)
);

AO22x1_ASAP7_75t_L g13564 ( 
.A1(n_13404),
.A2(n_2264),
.B1(n_2262),
.B2(n_2263),
.Y(n_13564)
);

INVx2_ASAP7_75t_SL g13565 ( 
.A(n_13436),
.Y(n_13565)
);

OR4x1_ASAP7_75t_L g13566 ( 
.A(n_13440),
.B(n_2266),
.C(n_2264),
.D(n_2265),
.Y(n_13566)
);

INVx2_ASAP7_75t_L g13567 ( 
.A(n_13455),
.Y(n_13567)
);

NOR2x1_ASAP7_75t_L g13568 ( 
.A(n_13425),
.B(n_2265),
.Y(n_13568)
);

INVx1_ASAP7_75t_L g13569 ( 
.A(n_13378),
.Y(n_13569)
);

AND2x2_ASAP7_75t_L g13570 ( 
.A(n_13413),
.B(n_2266),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_13444),
.Y(n_13571)
);

OAI22xp5_ASAP7_75t_L g13572 ( 
.A1(n_13439),
.A2(n_2269),
.B1(n_2267),
.B2(n_2268),
.Y(n_13572)
);

INVx1_ASAP7_75t_L g13573 ( 
.A(n_13465),
.Y(n_13573)
);

OAI211xp5_ASAP7_75t_L g13574 ( 
.A1(n_13441),
.A2(n_13447),
.B(n_13451),
.C(n_13443),
.Y(n_13574)
);

OAI31xp33_ASAP7_75t_L g13575 ( 
.A1(n_13405),
.A2(n_2269),
.A3(n_2267),
.B(n_2268),
.Y(n_13575)
);

OAI22xp5_ASAP7_75t_L g13576 ( 
.A1(n_13389),
.A2(n_2272),
.B1(n_2270),
.B2(n_2271),
.Y(n_13576)
);

AOI32xp33_ASAP7_75t_L g13577 ( 
.A1(n_13393),
.A2(n_2272),
.A3(n_2270),
.B1(n_2271),
.B2(n_2273),
.Y(n_13577)
);

NAND2xp5_ASAP7_75t_L g13578 ( 
.A(n_13361),
.B(n_2273),
.Y(n_13578)
);

NAND2xp5_ASAP7_75t_L g13579 ( 
.A(n_13398),
.B(n_2275),
.Y(n_13579)
);

OR2x2_ASAP7_75t_L g13580 ( 
.A(n_13392),
.B(n_2275),
.Y(n_13580)
);

NAND3xp33_ASAP7_75t_L g13581 ( 
.A(n_13448),
.B(n_2276),
.C(n_2277),
.Y(n_13581)
);

INVx1_ASAP7_75t_L g13582 ( 
.A(n_13408),
.Y(n_13582)
);

AOI211xp5_ASAP7_75t_L g13583 ( 
.A1(n_13422),
.A2(n_2278),
.B(n_2276),
.C(n_2277),
.Y(n_13583)
);

AOI221xp5_ASAP7_75t_L g13584 ( 
.A1(n_13401),
.A2(n_2281),
.B1(n_2279),
.B2(n_2280),
.C(n_2282),
.Y(n_13584)
);

INVx2_ASAP7_75t_SL g13585 ( 
.A(n_13416),
.Y(n_13585)
);

NAND2xp5_ASAP7_75t_L g13586 ( 
.A(n_13460),
.B(n_2279),
.Y(n_13586)
);

NAND2xp5_ASAP7_75t_L g13587 ( 
.A(n_13386),
.B(n_2281),
.Y(n_13587)
);

INVx2_ASAP7_75t_SL g13588 ( 
.A(n_13433),
.Y(n_13588)
);

INVx1_ASAP7_75t_L g13589 ( 
.A(n_13458),
.Y(n_13589)
);

AOI22xp5_ASAP7_75t_L g13590 ( 
.A1(n_13437),
.A2(n_2285),
.B1(n_2283),
.B2(n_2284),
.Y(n_13590)
);

AOI32xp33_ASAP7_75t_L g13591 ( 
.A1(n_13369),
.A2(n_2285),
.A3(n_2283),
.B1(n_2284),
.B2(n_2286),
.Y(n_13591)
);

INVx1_ASAP7_75t_L g13592 ( 
.A(n_13442),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_13449),
.Y(n_13593)
);

AOI322xp5_ASAP7_75t_L g13594 ( 
.A1(n_13452),
.A2(n_2291),
.A3(n_2290),
.B1(n_2288),
.B2(n_2286),
.C1(n_2287),
.C2(n_2289),
.Y(n_13594)
);

OAI22xp5_ASAP7_75t_L g13595 ( 
.A1(n_13383),
.A2(n_2290),
.B1(n_2288),
.B2(n_2289),
.Y(n_13595)
);

INVx2_ASAP7_75t_L g13596 ( 
.A(n_13446),
.Y(n_13596)
);

AOI22xp5_ASAP7_75t_L g13597 ( 
.A1(n_13459),
.A2(n_13385),
.B1(n_13431),
.B2(n_13429),
.Y(n_13597)
);

INVx2_ASAP7_75t_SL g13598 ( 
.A(n_13428),
.Y(n_13598)
);

NAND2xp5_ASAP7_75t_L g13599 ( 
.A(n_13338),
.B(n_2291),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_13472),
.Y(n_13600)
);

AND2x2_ASAP7_75t_L g13601 ( 
.A(n_13432),
.B(n_2292),
.Y(n_13601)
);

OAI22xp33_ASAP7_75t_L g13602 ( 
.A1(n_13462),
.A2(n_13467),
.B1(n_13463),
.B2(n_13469),
.Y(n_13602)
);

INVx2_ASAP7_75t_L g13603 ( 
.A(n_13471),
.Y(n_13603)
);

INVx1_ASAP7_75t_L g13604 ( 
.A(n_13370),
.Y(n_13604)
);

NAND2xp5_ASAP7_75t_L g13605 ( 
.A(n_13346),
.B(n_2292),
.Y(n_13605)
);

INVx2_ASAP7_75t_L g13606 ( 
.A(n_13468),
.Y(n_13606)
);

NAND2x1p5_ASAP7_75t_L g13607 ( 
.A(n_13368),
.B(n_2293),
.Y(n_13607)
);

HB1xp67_ASAP7_75t_L g13608 ( 
.A(n_13430),
.Y(n_13608)
);

INVx1_ASAP7_75t_SL g13609 ( 
.A(n_13486),
.Y(n_13609)
);

INVx2_ASAP7_75t_L g13610 ( 
.A(n_13607),
.Y(n_13610)
);

OAI22xp5_ASAP7_75t_L g13611 ( 
.A1(n_13507),
.A2(n_13495),
.B1(n_13503),
.B2(n_13496),
.Y(n_13611)
);

OAI22xp5_ASAP7_75t_L g13612 ( 
.A1(n_13516),
.A2(n_2296),
.B1(n_2294),
.B2(n_2295),
.Y(n_13612)
);

AND2x2_ASAP7_75t_L g13613 ( 
.A(n_13606),
.B(n_2294),
.Y(n_13613)
);

INVxp67_ASAP7_75t_SL g13614 ( 
.A(n_13608),
.Y(n_13614)
);

OAI22xp5_ASAP7_75t_L g13615 ( 
.A1(n_13482),
.A2(n_2297),
.B1(n_2295),
.B2(n_2296),
.Y(n_13615)
);

OR2x2_ASAP7_75t_L g13616 ( 
.A(n_13476),
.B(n_2297),
.Y(n_13616)
);

INVx2_ASAP7_75t_L g13617 ( 
.A(n_13497),
.Y(n_13617)
);

INVx1_ASAP7_75t_L g13618 ( 
.A(n_13510),
.Y(n_13618)
);

NAND2xp5_ASAP7_75t_SL g13619 ( 
.A(n_13575),
.B(n_13540),
.Y(n_13619)
);

NAND2xp5_ASAP7_75t_L g13620 ( 
.A(n_13564),
.B(n_2298),
.Y(n_13620)
);

INVx1_ASAP7_75t_L g13621 ( 
.A(n_13475),
.Y(n_13621)
);

INVx1_ASAP7_75t_SL g13622 ( 
.A(n_13537),
.Y(n_13622)
);

AND2x2_ASAP7_75t_L g13623 ( 
.A(n_13540),
.B(n_2298),
.Y(n_13623)
);

OAI33xp33_ASAP7_75t_L g13624 ( 
.A1(n_13602),
.A2(n_2303),
.A3(n_2305),
.B1(n_2299),
.B2(n_2301),
.B3(n_2304),
.Y(n_13624)
);

AOI21xp33_ASAP7_75t_L g13625 ( 
.A1(n_13498),
.A2(n_13480),
.B(n_13604),
.Y(n_13625)
);

OR2x2_ASAP7_75t_L g13626 ( 
.A(n_13553),
.B(n_2299),
.Y(n_13626)
);

OA21x2_ASAP7_75t_SL g13627 ( 
.A1(n_13499),
.A2(n_2301),
.B(n_2303),
.Y(n_13627)
);

INVx2_ASAP7_75t_L g13628 ( 
.A(n_13566),
.Y(n_13628)
);

NAND2xp5_ASAP7_75t_L g13629 ( 
.A(n_13554),
.B(n_2305),
.Y(n_13629)
);

AND2x2_ASAP7_75t_L g13630 ( 
.A(n_13554),
.B(n_2306),
.Y(n_13630)
);

OAI22xp33_ASAP7_75t_L g13631 ( 
.A1(n_13522),
.A2(n_2309),
.B1(n_2306),
.B2(n_2308),
.Y(n_13631)
);

OAI21xp33_ASAP7_75t_L g13632 ( 
.A1(n_13558),
.A2(n_2308),
.B(n_2310),
.Y(n_13632)
);

AOI21xp5_ASAP7_75t_L g13633 ( 
.A1(n_13586),
.A2(n_2310),
.B(n_2312),
.Y(n_13633)
);

NOR2xp33_ASAP7_75t_L g13634 ( 
.A(n_13479),
.B(n_2313),
.Y(n_13634)
);

AOI22xp5_ASAP7_75t_L g13635 ( 
.A1(n_13493),
.A2(n_2315),
.B1(n_2313),
.B2(n_2314),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_13528),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_13519),
.Y(n_13637)
);

INVx1_ASAP7_75t_L g13638 ( 
.A(n_13570),
.Y(n_13638)
);

NAND2xp5_ASAP7_75t_L g13639 ( 
.A(n_13502),
.B(n_2314),
.Y(n_13639)
);

AND2x2_ASAP7_75t_L g13640 ( 
.A(n_13509),
.B(n_2316),
.Y(n_13640)
);

INVxp67_ASAP7_75t_L g13641 ( 
.A(n_13544),
.Y(n_13641)
);

OAI21xp5_ASAP7_75t_L g13642 ( 
.A1(n_13511),
.A2(n_2316),
.B(n_2317),
.Y(n_13642)
);

AND2x2_ASAP7_75t_L g13643 ( 
.A(n_13488),
.B(n_2318),
.Y(n_13643)
);

AND2x2_ASAP7_75t_L g13644 ( 
.A(n_13490),
.B(n_2319),
.Y(n_13644)
);

OAI32xp33_ASAP7_75t_L g13645 ( 
.A1(n_13492),
.A2(n_2323),
.A3(n_2321),
.B1(n_2322),
.B2(n_2324),
.Y(n_13645)
);

INVx1_ASAP7_75t_L g13646 ( 
.A(n_13526),
.Y(n_13646)
);

AOI22xp5_ASAP7_75t_L g13647 ( 
.A1(n_13565),
.A2(n_2323),
.B1(n_2321),
.B2(n_2322),
.Y(n_13647)
);

AND2x2_ASAP7_75t_L g13648 ( 
.A(n_13481),
.B(n_2325),
.Y(n_13648)
);

AOI21xp5_ASAP7_75t_L g13649 ( 
.A1(n_13556),
.A2(n_2325),
.B(n_2326),
.Y(n_13649)
);

NOR2xp33_ASAP7_75t_SL g13650 ( 
.A(n_13524),
.B(n_2326),
.Y(n_13650)
);

NAND2xp5_ASAP7_75t_L g13651 ( 
.A(n_13539),
.B(n_2328),
.Y(n_13651)
);

NAND2xp5_ASAP7_75t_L g13652 ( 
.A(n_13508),
.B(n_2329),
.Y(n_13652)
);

AND2x2_ASAP7_75t_L g13653 ( 
.A(n_13484),
.B(n_2329),
.Y(n_13653)
);

O2A1O1Ixp5_ASAP7_75t_L g13654 ( 
.A1(n_13574),
.A2(n_2332),
.B(n_2330),
.C(n_2331),
.Y(n_13654)
);

OR2x2_ASAP7_75t_L g13655 ( 
.A(n_13491),
.B(n_2330),
.Y(n_13655)
);

NAND2xp5_ASAP7_75t_L g13656 ( 
.A(n_13536),
.B(n_2331),
.Y(n_13656)
);

NAND2xp5_ASAP7_75t_L g13657 ( 
.A(n_13577),
.B(n_2332),
.Y(n_13657)
);

AND2x4_ASAP7_75t_L g13658 ( 
.A(n_13505),
.B(n_2333),
.Y(n_13658)
);

INVx1_ASAP7_75t_L g13659 ( 
.A(n_13605),
.Y(n_13659)
);

OR2x2_ASAP7_75t_L g13660 ( 
.A(n_13532),
.B(n_2333),
.Y(n_13660)
);

OAI322xp33_ASAP7_75t_L g13661 ( 
.A1(n_13501),
.A2(n_2339),
.A3(n_2338),
.B1(n_2336),
.B2(n_2334),
.C1(n_2335),
.C2(n_2337),
.Y(n_13661)
);

OAI21xp5_ASAP7_75t_L g13662 ( 
.A1(n_13568),
.A2(n_2334),
.B(n_2335),
.Y(n_13662)
);

AO21x1_ASAP7_75t_L g13663 ( 
.A1(n_13477),
.A2(n_2336),
.B(n_2337),
.Y(n_13663)
);

NAND2xp5_ASAP7_75t_L g13664 ( 
.A(n_13551),
.B(n_2338),
.Y(n_13664)
);

INVx1_ASAP7_75t_L g13665 ( 
.A(n_13483),
.Y(n_13665)
);

NAND2x1_ASAP7_75t_SL g13666 ( 
.A(n_13529),
.B(n_2339),
.Y(n_13666)
);

NAND2x1_ASAP7_75t_SL g13667 ( 
.A(n_13523),
.B(n_2340),
.Y(n_13667)
);

INVx1_ASAP7_75t_SL g13668 ( 
.A(n_13580),
.Y(n_13668)
);

NAND2xp5_ASAP7_75t_L g13669 ( 
.A(n_13521),
.B(n_2340),
.Y(n_13669)
);

INVx1_ASAP7_75t_L g13670 ( 
.A(n_13489),
.Y(n_13670)
);

NAND2xp5_ASAP7_75t_L g13671 ( 
.A(n_13591),
.B(n_2341),
.Y(n_13671)
);

OAI21xp5_ASAP7_75t_L g13672 ( 
.A1(n_13597),
.A2(n_2341),
.B(n_2342),
.Y(n_13672)
);

OAI21xp33_ASAP7_75t_L g13673 ( 
.A1(n_13603),
.A2(n_2342),
.B(n_2343),
.Y(n_13673)
);

NOR2x1_ASAP7_75t_L g13674 ( 
.A(n_13474),
.B(n_2344),
.Y(n_13674)
);

OAI21xp33_ASAP7_75t_L g13675 ( 
.A1(n_13500),
.A2(n_13541),
.B(n_13534),
.Y(n_13675)
);

HB1xp67_ASAP7_75t_L g13676 ( 
.A(n_13560),
.Y(n_13676)
);

AOI21xp33_ASAP7_75t_SL g13677 ( 
.A1(n_13527),
.A2(n_2344),
.B(n_2345),
.Y(n_13677)
);

OAI22xp5_ASAP7_75t_L g13678 ( 
.A1(n_13590),
.A2(n_2348),
.B1(n_2345),
.B2(n_2347),
.Y(n_13678)
);

AOI21xp5_ASAP7_75t_SL g13679 ( 
.A1(n_13557),
.A2(n_2348),
.B(n_2349),
.Y(n_13679)
);

INVx1_ASAP7_75t_L g13680 ( 
.A(n_13487),
.Y(n_13680)
);

INVx2_ASAP7_75t_L g13681 ( 
.A(n_13545),
.Y(n_13681)
);

AOI22xp5_ASAP7_75t_L g13682 ( 
.A1(n_13542),
.A2(n_13555),
.B1(n_13548),
.B2(n_13571),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_13547),
.Y(n_13683)
);

OAI32xp33_ASAP7_75t_L g13684 ( 
.A1(n_13578),
.A2(n_2351),
.A3(n_2349),
.B1(n_2350),
.B2(n_2352),
.Y(n_13684)
);

INVx1_ASAP7_75t_L g13685 ( 
.A(n_13512),
.Y(n_13685)
);

AND2x2_ASAP7_75t_L g13686 ( 
.A(n_13573),
.B(n_2350),
.Y(n_13686)
);

INVx1_ASAP7_75t_L g13687 ( 
.A(n_13494),
.Y(n_13687)
);

OR2x2_ASAP7_75t_L g13688 ( 
.A(n_13533),
.B(n_2351),
.Y(n_13688)
);

NOR2xp33_ASAP7_75t_SL g13689 ( 
.A(n_13478),
.B(n_2352),
.Y(n_13689)
);

O2A1O1Ixp5_ASAP7_75t_L g13690 ( 
.A1(n_13546),
.A2(n_2356),
.B(n_2353),
.C(n_2355),
.Y(n_13690)
);

AOI21xp33_ASAP7_75t_L g13691 ( 
.A1(n_13598),
.A2(n_2356),
.B(n_2357),
.Y(n_13691)
);

NAND2xp5_ASAP7_75t_L g13692 ( 
.A(n_13601),
.B(n_2357),
.Y(n_13692)
);

OAI322xp33_ASAP7_75t_L g13693 ( 
.A1(n_13518),
.A2(n_2365),
.A3(n_2363),
.B1(n_2361),
.B2(n_2359),
.C1(n_2360),
.C2(n_2362),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_13517),
.Y(n_13694)
);

AND2x2_ASAP7_75t_L g13695 ( 
.A(n_13520),
.B(n_13543),
.Y(n_13695)
);

OAI221xp5_ASAP7_75t_L g13696 ( 
.A1(n_13579),
.A2(n_13587),
.B1(n_13583),
.B2(n_13549),
.C(n_13514),
.Y(n_13696)
);

AND2x4_ASAP7_75t_L g13697 ( 
.A(n_13585),
.B(n_2359),
.Y(n_13697)
);

INVx1_ASAP7_75t_L g13698 ( 
.A(n_13552),
.Y(n_13698)
);

INVx1_ASAP7_75t_L g13699 ( 
.A(n_13599),
.Y(n_13699)
);

OAI32xp33_ASAP7_75t_L g13700 ( 
.A1(n_13561),
.A2(n_2363),
.A3(n_2361),
.B1(n_2362),
.B2(n_2365),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_13581),
.Y(n_13701)
);

INVxp67_ASAP7_75t_L g13702 ( 
.A(n_13572),
.Y(n_13702)
);

NAND3xp33_ASAP7_75t_L g13703 ( 
.A(n_13485),
.B(n_2366),
.C(n_2368),
.Y(n_13703)
);

AND2x2_ASAP7_75t_L g13704 ( 
.A(n_13567),
.B(n_2366),
.Y(n_13704)
);

OAI22xp5_ASAP7_75t_L g13705 ( 
.A1(n_13550),
.A2(n_2370),
.B1(n_2368),
.B2(n_2369),
.Y(n_13705)
);

AND2x2_ASAP7_75t_L g13706 ( 
.A(n_13596),
.B(n_2369),
.Y(n_13706)
);

AOI211xp5_ASAP7_75t_L g13707 ( 
.A1(n_13525),
.A2(n_2373),
.B(n_2370),
.C(n_2372),
.Y(n_13707)
);

INVx1_ASAP7_75t_L g13708 ( 
.A(n_13513),
.Y(n_13708)
);

INVx1_ASAP7_75t_L g13709 ( 
.A(n_13515),
.Y(n_13709)
);

INVx3_ASAP7_75t_L g13710 ( 
.A(n_13588),
.Y(n_13710)
);

NAND2xp5_ASAP7_75t_L g13711 ( 
.A(n_13506),
.B(n_2372),
.Y(n_13711)
);

INVxp67_ASAP7_75t_L g13712 ( 
.A(n_13576),
.Y(n_13712)
);

AOI21xp5_ASAP7_75t_L g13713 ( 
.A1(n_13531),
.A2(n_2374),
.B(n_2375),
.Y(n_13713)
);

INVx1_ASAP7_75t_L g13714 ( 
.A(n_13595),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_13589),
.Y(n_13715)
);

BUFx2_ASAP7_75t_L g13716 ( 
.A(n_13592),
.Y(n_13716)
);

AOI221xp5_ASAP7_75t_L g13717 ( 
.A1(n_13582),
.A2(n_2376),
.B1(n_2374),
.B2(n_2375),
.C(n_2377),
.Y(n_13717)
);

NOR2xp67_ASAP7_75t_L g13718 ( 
.A(n_13530),
.B(n_2376),
.Y(n_13718)
);

NAND2xp5_ASAP7_75t_L g13719 ( 
.A(n_13504),
.B(n_2377),
.Y(n_13719)
);

AND2x2_ASAP7_75t_L g13720 ( 
.A(n_13593),
.B(n_2378),
.Y(n_13720)
);

AND2x4_ASAP7_75t_L g13721 ( 
.A(n_13535),
.B(n_2378),
.Y(n_13721)
);

NAND2xp5_ASAP7_75t_L g13722 ( 
.A(n_13594),
.B(n_2379),
.Y(n_13722)
);

NAND2xp5_ASAP7_75t_L g13723 ( 
.A(n_13538),
.B(n_2379),
.Y(n_13723)
);

OAI22xp5_ASAP7_75t_L g13724 ( 
.A1(n_13559),
.A2(n_2382),
.B1(n_2380),
.B2(n_2381),
.Y(n_13724)
);

AOI221xp5_ASAP7_75t_L g13725 ( 
.A1(n_13569),
.A2(n_2383),
.B1(n_2381),
.B2(n_2382),
.C(n_2385),
.Y(n_13725)
);

AOI21xp5_ASAP7_75t_L g13726 ( 
.A1(n_13562),
.A2(n_2383),
.B(n_2385),
.Y(n_13726)
);

NAND2xp5_ASAP7_75t_L g13727 ( 
.A(n_13584),
.B(n_2386),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_13563),
.Y(n_13728)
);

INVx1_ASAP7_75t_L g13729 ( 
.A(n_13600),
.Y(n_13729)
);

INVx1_ASAP7_75t_L g13730 ( 
.A(n_13608),
.Y(n_13730)
);

INVx1_ASAP7_75t_L g13731 ( 
.A(n_13608),
.Y(n_13731)
);

AND2x4_ASAP7_75t_L g13732 ( 
.A(n_13540),
.B(n_2386),
.Y(n_13732)
);

INVxp67_ASAP7_75t_L g13733 ( 
.A(n_13608),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_13608),
.Y(n_13734)
);

NAND2xp5_ASAP7_75t_SL g13735 ( 
.A(n_13663),
.B(n_2387),
.Y(n_13735)
);

AOI22xp5_ASAP7_75t_L g13736 ( 
.A1(n_13609),
.A2(n_13614),
.B1(n_13733),
.B2(n_13731),
.Y(n_13736)
);

NOR3xp33_ASAP7_75t_L g13737 ( 
.A(n_13625),
.B(n_2387),
.C(n_2388),
.Y(n_13737)
);

AOI221xp5_ASAP7_75t_L g13738 ( 
.A1(n_13611),
.A2(n_2391),
.B1(n_2389),
.B2(n_2390),
.C(n_2392),
.Y(n_13738)
);

AOI22xp33_ASAP7_75t_L g13739 ( 
.A1(n_13730),
.A2(n_2392),
.B1(n_2390),
.B2(n_2391),
.Y(n_13739)
);

OR2x2_ASAP7_75t_L g13740 ( 
.A(n_13626),
.B(n_2393),
.Y(n_13740)
);

AO22x1_ASAP7_75t_L g13741 ( 
.A1(n_13662),
.A2(n_2395),
.B1(n_2393),
.B2(n_2394),
.Y(n_13741)
);

INVx1_ASAP7_75t_L g13742 ( 
.A(n_13666),
.Y(n_13742)
);

AOI21xp5_ASAP7_75t_L g13743 ( 
.A1(n_13619),
.A2(n_2395),
.B(n_2396),
.Y(n_13743)
);

NAND2xp5_ASAP7_75t_SL g13744 ( 
.A(n_13734),
.B(n_2396),
.Y(n_13744)
);

AO22x1_ASAP7_75t_L g13745 ( 
.A1(n_13674),
.A2(n_2399),
.B1(n_2397),
.B2(n_2398),
.Y(n_13745)
);

OAI21xp5_ASAP7_75t_SL g13746 ( 
.A1(n_13682),
.A2(n_2397),
.B(n_2398),
.Y(n_13746)
);

NAND4xp25_ASAP7_75t_SL g13747 ( 
.A(n_13707),
.B(n_13622),
.C(n_13722),
.D(n_13679),
.Y(n_13747)
);

AOI22xp5_ASAP7_75t_L g13748 ( 
.A1(n_13675),
.A2(n_2401),
.B1(n_2399),
.B2(n_2400),
.Y(n_13748)
);

INVx1_ASAP7_75t_L g13749 ( 
.A(n_13667),
.Y(n_13749)
);

AND3x2_ASAP7_75t_L g13750 ( 
.A(n_13716),
.B(n_13697),
.C(n_13630),
.Y(n_13750)
);

AOI22xp5_ASAP7_75t_L g13751 ( 
.A1(n_13710),
.A2(n_2402),
.B1(n_2400),
.B2(n_2401),
.Y(n_13751)
);

OAI22xp5_ASAP7_75t_L g13752 ( 
.A1(n_13712),
.A2(n_2404),
.B1(n_2402),
.B2(n_2403),
.Y(n_13752)
);

INVx1_ASAP7_75t_L g13753 ( 
.A(n_13623),
.Y(n_13753)
);

OR2x2_ASAP7_75t_L g13754 ( 
.A(n_13629),
.B(n_2403),
.Y(n_13754)
);

OAI21xp5_ASAP7_75t_L g13755 ( 
.A1(n_13654),
.A2(n_2404),
.B(n_2405),
.Y(n_13755)
);

NOR3xp33_ASAP7_75t_L g13756 ( 
.A(n_13696),
.B(n_2413),
.C(n_2405),
.Y(n_13756)
);

INVxp67_ASAP7_75t_L g13757 ( 
.A(n_13650),
.Y(n_13757)
);

INVx1_ASAP7_75t_SL g13758 ( 
.A(n_13616),
.Y(n_13758)
);

INVx1_ASAP7_75t_L g13759 ( 
.A(n_13732),
.Y(n_13759)
);

INVx1_ASAP7_75t_L g13760 ( 
.A(n_13697),
.Y(n_13760)
);

OAI21xp33_ASAP7_75t_SL g13761 ( 
.A1(n_13637),
.A2(n_3463),
.B(n_3455),
.Y(n_13761)
);

NAND2xp5_ASAP7_75t_L g13762 ( 
.A(n_13644),
.B(n_2406),
.Y(n_13762)
);

NAND2x1_ASAP7_75t_L g13763 ( 
.A(n_13658),
.B(n_13610),
.Y(n_13763)
);

AND2x2_ASAP7_75t_L g13764 ( 
.A(n_13613),
.B(n_2406),
.Y(n_13764)
);

AOI22xp5_ASAP7_75t_L g13765 ( 
.A1(n_13689),
.A2(n_2409),
.B1(n_2407),
.B2(n_2408),
.Y(n_13765)
);

OAI221xp5_ASAP7_75t_L g13766 ( 
.A1(n_13672),
.A2(n_2425),
.B1(n_2433),
.B2(n_2416),
.C(n_2407),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_13648),
.Y(n_13767)
);

INVx1_ASAP7_75t_L g13768 ( 
.A(n_13653),
.Y(n_13768)
);

OR2x2_ASAP7_75t_L g13769 ( 
.A(n_13620),
.B(n_2408),
.Y(n_13769)
);

AOI22xp5_ASAP7_75t_L g13770 ( 
.A1(n_13695),
.A2(n_2411),
.B1(n_2409),
.B2(n_2410),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_13658),
.Y(n_13771)
);

OR2x2_ASAP7_75t_L g13772 ( 
.A(n_13628),
.B(n_2410),
.Y(n_13772)
);

INVx1_ASAP7_75t_L g13773 ( 
.A(n_13640),
.Y(n_13773)
);

OR2x2_ASAP7_75t_L g13774 ( 
.A(n_13692),
.B(n_2411),
.Y(n_13774)
);

OAI221xp5_ASAP7_75t_L g13775 ( 
.A1(n_13642),
.A2(n_2430),
.B1(n_2439),
.B2(n_2421),
.C(n_2412),
.Y(n_13775)
);

AOI21xp5_ASAP7_75t_SL g13776 ( 
.A1(n_13661),
.A2(n_2412),
.B(n_2414),
.Y(n_13776)
);

INVx2_ASAP7_75t_L g13777 ( 
.A(n_13721),
.Y(n_13777)
);

NAND2xp33_ASAP7_75t_L g13778 ( 
.A(n_13632),
.B(n_2415),
.Y(n_13778)
);

AND2x2_ASAP7_75t_L g13779 ( 
.A(n_13617),
.B(n_2415),
.Y(n_13779)
);

INVx2_ASAP7_75t_L g13780 ( 
.A(n_13721),
.Y(n_13780)
);

NAND2xp5_ASAP7_75t_L g13781 ( 
.A(n_13686),
.B(n_2416),
.Y(n_13781)
);

INVx1_ASAP7_75t_L g13782 ( 
.A(n_13643),
.Y(n_13782)
);

AOI221xp5_ASAP7_75t_SL g13783 ( 
.A1(n_13677),
.A2(n_2419),
.B1(n_2417),
.B2(n_2418),
.C(n_2420),
.Y(n_13783)
);

OR2x2_ASAP7_75t_L g13784 ( 
.A(n_13639),
.B(n_2418),
.Y(n_13784)
);

INVx1_ASAP7_75t_L g13785 ( 
.A(n_13720),
.Y(n_13785)
);

AOI21xp33_ASAP7_75t_SL g13786 ( 
.A1(n_13703),
.A2(n_2424),
.B(n_2422),
.Y(n_13786)
);

INVx1_ASAP7_75t_L g13787 ( 
.A(n_13704),
.Y(n_13787)
);

INVx2_ASAP7_75t_L g13788 ( 
.A(n_13706),
.Y(n_13788)
);

NAND4xp25_ASAP7_75t_L g13789 ( 
.A(n_13627),
.B(n_13718),
.C(n_13702),
.D(n_13714),
.Y(n_13789)
);

INVx1_ASAP7_75t_SL g13790 ( 
.A(n_13668),
.Y(n_13790)
);

AND2x2_ASAP7_75t_L g13791 ( 
.A(n_13618),
.B(n_2420),
.Y(n_13791)
);

A2O1A1Ixp33_ASAP7_75t_L g13792 ( 
.A1(n_13690),
.A2(n_2426),
.B(n_2424),
.C(n_2425),
.Y(n_13792)
);

INVx1_ASAP7_75t_L g13793 ( 
.A(n_13652),
.Y(n_13793)
);

NAND3xp33_ASAP7_75t_SL g13794 ( 
.A(n_13713),
.B(n_2426),
.C(n_2427),
.Y(n_13794)
);

INVx2_ASAP7_75t_L g13795 ( 
.A(n_13655),
.Y(n_13795)
);

NAND2xp5_ASAP7_75t_L g13796 ( 
.A(n_13726),
.B(n_2427),
.Y(n_13796)
);

AOI21xp33_ASAP7_75t_SL g13797 ( 
.A1(n_13631),
.A2(n_2431),
.B(n_2429),
.Y(n_13797)
);

NAND2xp5_ASAP7_75t_L g13798 ( 
.A(n_13636),
.B(n_2428),
.Y(n_13798)
);

OAI21xp33_ASAP7_75t_L g13799 ( 
.A1(n_13715),
.A2(n_2428),
.B(n_2429),
.Y(n_13799)
);

OR2x2_ASAP7_75t_L g13800 ( 
.A(n_13651),
.B(n_2431),
.Y(n_13800)
);

INVx1_ASAP7_75t_L g13801 ( 
.A(n_13711),
.Y(n_13801)
);

OAI22xp5_ASAP7_75t_L g13802 ( 
.A1(n_13657),
.A2(n_2435),
.B1(n_2432),
.B2(n_2434),
.Y(n_13802)
);

OAI22xp5_ASAP7_75t_L g13803 ( 
.A1(n_13671),
.A2(n_2436),
.B1(n_2432),
.B2(n_2435),
.Y(n_13803)
);

OAI21xp5_ASAP7_75t_L g13804 ( 
.A1(n_13656),
.A2(n_2437),
.B(n_2438),
.Y(n_13804)
);

OR2x2_ASAP7_75t_L g13805 ( 
.A(n_13688),
.B(n_2437),
.Y(n_13805)
);

AOI22xp5_ASAP7_75t_L g13806 ( 
.A1(n_13634),
.A2(n_2441),
.B1(n_2438),
.B2(n_2440),
.Y(n_13806)
);

OAI31xp33_ASAP7_75t_L g13807 ( 
.A1(n_13673),
.A2(n_2442),
.A3(n_2440),
.B(n_2441),
.Y(n_13807)
);

AOI22xp5_ASAP7_75t_L g13808 ( 
.A1(n_13638),
.A2(n_2445),
.B1(n_2443),
.B2(n_2444),
.Y(n_13808)
);

NAND2xp33_ASAP7_75t_L g13809 ( 
.A(n_13646),
.B(n_2444),
.Y(n_13809)
);

AOI22xp33_ASAP7_75t_L g13810 ( 
.A1(n_13708),
.A2(n_2448),
.B1(n_2446),
.B2(n_2447),
.Y(n_13810)
);

INVx1_ASAP7_75t_L g13811 ( 
.A(n_13669),
.Y(n_13811)
);

NAND2xp5_ASAP7_75t_L g13812 ( 
.A(n_13649),
.B(n_2446),
.Y(n_13812)
);

INVx1_ASAP7_75t_L g13813 ( 
.A(n_13660),
.Y(n_13813)
);

INVxp67_ASAP7_75t_L g13814 ( 
.A(n_13624),
.Y(n_13814)
);

NAND2xp5_ASAP7_75t_L g13815 ( 
.A(n_13647),
.B(n_2447),
.Y(n_13815)
);

INVx2_ASAP7_75t_SL g13816 ( 
.A(n_13621),
.Y(n_13816)
);

INVx1_ASAP7_75t_L g13817 ( 
.A(n_13664),
.Y(n_13817)
);

AOI22xp5_ASAP7_75t_L g13818 ( 
.A1(n_13709),
.A2(n_2450),
.B1(n_2448),
.B2(n_2449),
.Y(n_13818)
);

AND2x2_ASAP7_75t_L g13819 ( 
.A(n_13701),
.B(n_2449),
.Y(n_13819)
);

AND2x2_ASAP7_75t_L g13820 ( 
.A(n_13676),
.B(n_2451),
.Y(n_13820)
);

OAI22xp33_ASAP7_75t_L g13821 ( 
.A1(n_13719),
.A2(n_2454),
.B1(n_2452),
.B2(n_2453),
.Y(n_13821)
);

NAND2xp5_ASAP7_75t_L g13822 ( 
.A(n_13633),
.B(n_2452),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_13681),
.B(n_13698),
.Y(n_13823)
);

AOI21xp33_ASAP7_75t_L g13824 ( 
.A1(n_13727),
.A2(n_2453),
.B(n_2454),
.Y(n_13824)
);

INVx1_ASAP7_75t_L g13825 ( 
.A(n_13723),
.Y(n_13825)
);

NAND2xp5_ASAP7_75t_SL g13826 ( 
.A(n_13691),
.B(n_2455),
.Y(n_13826)
);

OAI21xp33_ASAP7_75t_L g13827 ( 
.A1(n_13680),
.A2(n_2455),
.B(n_2456),
.Y(n_13827)
);

AND2x2_ASAP7_75t_L g13828 ( 
.A(n_13641),
.B(n_2456),
.Y(n_13828)
);

NOR2xp33_ASAP7_75t_L g13829 ( 
.A(n_13684),
.B(n_13705),
.Y(n_13829)
);

NOR2xp33_ASAP7_75t_L g13830 ( 
.A(n_13645),
.B(n_2457),
.Y(n_13830)
);

OAI21xp5_ASAP7_75t_L g13831 ( 
.A1(n_13728),
.A2(n_13729),
.B(n_13665),
.Y(n_13831)
);

INVx1_ASAP7_75t_L g13832 ( 
.A(n_13615),
.Y(n_13832)
);

NOR2xp33_ASAP7_75t_L g13833 ( 
.A(n_13678),
.B(n_2457),
.Y(n_13833)
);

OAI221xp5_ASAP7_75t_L g13834 ( 
.A1(n_13699),
.A2(n_2474),
.B1(n_2483),
.B2(n_2466),
.C(n_2458),
.Y(n_13834)
);

AOI22xp33_ASAP7_75t_L g13835 ( 
.A1(n_13694),
.A2(n_2460),
.B1(n_2458),
.B2(n_2459),
.Y(n_13835)
);

NOR2xp33_ASAP7_75t_L g13836 ( 
.A(n_13693),
.B(n_2459),
.Y(n_13836)
);

NAND2xp5_ASAP7_75t_L g13837 ( 
.A(n_13635),
.B(n_13612),
.Y(n_13837)
);

INVx1_ASAP7_75t_L g13838 ( 
.A(n_13683),
.Y(n_13838)
);

NAND2xp33_ASAP7_75t_SL g13839 ( 
.A(n_13659),
.B(n_2460),
.Y(n_13839)
);

OR2x2_ASAP7_75t_L g13840 ( 
.A(n_13670),
.B(n_2461),
.Y(n_13840)
);

INVx1_ASAP7_75t_L g13841 ( 
.A(n_13724),
.Y(n_13841)
);

AND2x2_ASAP7_75t_L g13842 ( 
.A(n_13685),
.B(n_2462),
.Y(n_13842)
);

BUFx2_ASAP7_75t_L g13843 ( 
.A(n_13687),
.Y(n_13843)
);

OAI22xp5_ASAP7_75t_L g13844 ( 
.A1(n_13717),
.A2(n_2464),
.B1(n_2462),
.B2(n_2463),
.Y(n_13844)
);

NAND2xp5_ASAP7_75t_L g13845 ( 
.A(n_13725),
.B(n_2463),
.Y(n_13845)
);

INVx1_ASAP7_75t_L g13846 ( 
.A(n_13700),
.Y(n_13846)
);

NAND2xp5_ASAP7_75t_SL g13847 ( 
.A(n_13663),
.B(n_2464),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_13666),
.Y(n_13848)
);

INVx1_ASAP7_75t_L g13849 ( 
.A(n_13666),
.Y(n_13849)
);

INVx1_ASAP7_75t_L g13850 ( 
.A(n_13666),
.Y(n_13850)
);

OAI22xp5_ASAP7_75t_L g13851 ( 
.A1(n_13733),
.A2(n_2467),
.B1(n_2465),
.B2(n_2466),
.Y(n_13851)
);

NAND2xp5_ASAP7_75t_L g13852 ( 
.A(n_13614),
.B(n_2465),
.Y(n_13852)
);

INVx2_ASAP7_75t_L g13853 ( 
.A(n_13666),
.Y(n_13853)
);

INVx1_ASAP7_75t_SL g13854 ( 
.A(n_13667),
.Y(n_13854)
);

AOI221xp5_ASAP7_75t_L g13855 ( 
.A1(n_13625),
.A2(n_2470),
.B1(n_2468),
.B2(n_2469),
.C(n_2471),
.Y(n_13855)
);

AOI21xp5_ASAP7_75t_L g13856 ( 
.A1(n_13614),
.A2(n_2469),
.B(n_2470),
.Y(n_13856)
);

NOR2xp33_ASAP7_75t_L g13857 ( 
.A(n_13609),
.B(n_2471),
.Y(n_13857)
);

OAI322xp33_ASAP7_75t_L g13858 ( 
.A1(n_13733),
.A2(n_2477),
.A3(n_2476),
.B1(n_2474),
.B2(n_2472),
.C1(n_2473),
.C2(n_2475),
.Y(n_13858)
);

INVx2_ASAP7_75t_SL g13859 ( 
.A(n_13667),
.Y(n_13859)
);

XOR2x2_ASAP7_75t_L g13860 ( 
.A(n_13667),
.B(n_2472),
.Y(n_13860)
);

NAND2xp5_ASAP7_75t_SL g13861 ( 
.A(n_13663),
.B(n_2473),
.Y(n_13861)
);

AOI21xp5_ASAP7_75t_L g13862 ( 
.A1(n_13614),
.A2(n_2475),
.B(n_2476),
.Y(n_13862)
);

INVxp67_ASAP7_75t_L g13863 ( 
.A(n_13623),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_13614),
.B(n_2478),
.Y(n_13864)
);

OR2x2_ASAP7_75t_L g13865 ( 
.A(n_13859),
.B(n_2478),
.Y(n_13865)
);

NAND2xp5_ASAP7_75t_L g13866 ( 
.A(n_13750),
.B(n_2481),
.Y(n_13866)
);

AOI221xp5_ASAP7_75t_L g13867 ( 
.A1(n_13786),
.A2(n_13797),
.B1(n_13824),
.B2(n_13839),
.C(n_13745),
.Y(n_13867)
);

NAND2xp5_ASAP7_75t_L g13868 ( 
.A(n_13791),
.B(n_2481),
.Y(n_13868)
);

INVxp33_ASAP7_75t_L g13869 ( 
.A(n_13857),
.Y(n_13869)
);

NAND2xp5_ASAP7_75t_SL g13870 ( 
.A(n_13736),
.B(n_2480),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_13860),
.Y(n_13871)
);

AOI321xp33_ASAP7_75t_L g13872 ( 
.A1(n_13747),
.A2(n_2483),
.A3(n_2485),
.B1(n_2480),
.B2(n_2482),
.C(n_2484),
.Y(n_13872)
);

OAI32xp33_ASAP7_75t_L g13873 ( 
.A1(n_13761),
.A2(n_13864),
.A3(n_13852),
.B1(n_13854),
.B2(n_13737),
.Y(n_13873)
);

OAI22xp5_ASAP7_75t_L g13874 ( 
.A1(n_13748),
.A2(n_2486),
.B1(n_2482),
.B2(n_2484),
.Y(n_13874)
);

NAND3xp33_ASAP7_75t_L g13875 ( 
.A(n_13756),
.B(n_2486),
.C(n_2487),
.Y(n_13875)
);

OAI22xp33_ASAP7_75t_L g13876 ( 
.A1(n_13765),
.A2(n_13790),
.B1(n_13749),
.B2(n_13853),
.Y(n_13876)
);

AOI21xp5_ASAP7_75t_L g13877 ( 
.A1(n_13763),
.A2(n_13847),
.B(n_13735),
.Y(n_13877)
);

AOI322xp5_ASAP7_75t_L g13878 ( 
.A1(n_13846),
.A2(n_13836),
.A3(n_13829),
.B1(n_13814),
.B2(n_13816),
.C1(n_13758),
.C2(n_13778),
.Y(n_13878)
);

INVx1_ASAP7_75t_L g13879 ( 
.A(n_13764),
.Y(n_13879)
);

NAND2xp5_ASAP7_75t_L g13880 ( 
.A(n_13779),
.B(n_2489),
.Y(n_13880)
);

OAI32xp33_ASAP7_75t_L g13881 ( 
.A1(n_13769),
.A2(n_2490),
.A3(n_2488),
.B1(n_2489),
.B2(n_2491),
.Y(n_13881)
);

OAI32xp33_ASAP7_75t_L g13882 ( 
.A1(n_13796),
.A2(n_2492),
.A3(n_2488),
.B1(n_2490),
.B2(n_2493),
.Y(n_13882)
);

INVx1_ASAP7_75t_L g13883 ( 
.A(n_13772),
.Y(n_13883)
);

AOI222xp33_ASAP7_75t_L g13884 ( 
.A1(n_13861),
.A2(n_2495),
.B1(n_2497),
.B2(n_2492),
.C1(n_2494),
.C2(n_2496),
.Y(n_13884)
);

AOI22xp5_ASAP7_75t_L g13885 ( 
.A1(n_13823),
.A2(n_2496),
.B1(n_2494),
.B2(n_2495),
.Y(n_13885)
);

INVx2_ASAP7_75t_L g13886 ( 
.A(n_13740),
.Y(n_13886)
);

AOI311xp33_ASAP7_75t_L g13887 ( 
.A1(n_13742),
.A2(n_2499),
.A3(n_2497),
.B(n_2498),
.C(n_2500),
.Y(n_13887)
);

INVx1_ASAP7_75t_L g13888 ( 
.A(n_13840),
.Y(n_13888)
);

AOI22xp5_ASAP7_75t_L g13889 ( 
.A1(n_13759),
.A2(n_2500),
.B1(n_2498),
.B2(n_2499),
.Y(n_13889)
);

OR2x2_ASAP7_75t_L g13890 ( 
.A(n_13848),
.B(n_2501),
.Y(n_13890)
);

AOI32xp33_ASAP7_75t_L g13891 ( 
.A1(n_13849),
.A2(n_2503),
.A3(n_2501),
.B1(n_2502),
.B2(n_2505),
.Y(n_13891)
);

AND3x1_ASAP7_75t_L g13892 ( 
.A(n_13807),
.B(n_2502),
.C(n_2503),
.Y(n_13892)
);

INVx2_ASAP7_75t_L g13893 ( 
.A(n_13805),
.Y(n_13893)
);

INVx2_ASAP7_75t_L g13894 ( 
.A(n_13842),
.Y(n_13894)
);

INVx1_ASAP7_75t_L g13895 ( 
.A(n_13760),
.Y(n_13895)
);

AOI22xp5_ASAP7_75t_L g13896 ( 
.A1(n_13753),
.A2(n_2508),
.B1(n_2506),
.B2(n_2507),
.Y(n_13896)
);

NAND2xp5_ASAP7_75t_L g13897 ( 
.A(n_13741),
.B(n_2507),
.Y(n_13897)
);

NAND2xp5_ASAP7_75t_L g13898 ( 
.A(n_13820),
.B(n_2508),
.Y(n_13898)
);

AOI21xp5_ASAP7_75t_L g13899 ( 
.A1(n_13809),
.A2(n_2506),
.B(n_2509),
.Y(n_13899)
);

NOR2x1_ASAP7_75t_L g13900 ( 
.A(n_13789),
.B(n_13850),
.Y(n_13900)
);

AOI21xp5_ASAP7_75t_L g13901 ( 
.A1(n_13822),
.A2(n_2509),
.B(n_2510),
.Y(n_13901)
);

AOI322xp5_ASAP7_75t_L g13902 ( 
.A1(n_13832),
.A2(n_13841),
.A3(n_13757),
.B1(n_13830),
.B2(n_13768),
.C1(n_13767),
.C2(n_13785),
.Y(n_13902)
);

NAND2xp5_ASAP7_75t_L g13903 ( 
.A(n_13777),
.B(n_2512),
.Y(n_13903)
);

OAI221xp5_ASAP7_75t_SL g13904 ( 
.A1(n_13743),
.A2(n_2514),
.B1(n_2511),
.B2(n_2512),
.C(n_2515),
.Y(n_13904)
);

NOR2xp33_ASAP7_75t_L g13905 ( 
.A(n_13780),
.B(n_2515),
.Y(n_13905)
);

A2O1A1Ixp33_ASAP7_75t_L g13906 ( 
.A1(n_13856),
.A2(n_2520),
.B(n_2518),
.C(n_2519),
.Y(n_13906)
);

OAI21xp5_ASAP7_75t_SL g13907 ( 
.A1(n_13746),
.A2(n_2518),
.B(n_2521),
.Y(n_13907)
);

A2O1A1O1Ixp25_ASAP7_75t_L g13908 ( 
.A1(n_13771),
.A2(n_2523),
.B(n_2521),
.C(n_2522),
.D(n_2524),
.Y(n_13908)
);

OAI221xp5_ASAP7_75t_SL g13909 ( 
.A1(n_13776),
.A2(n_2524),
.B1(n_2522),
.B2(n_2523),
.C(n_2525),
.Y(n_13909)
);

OAI22xp33_ASAP7_75t_L g13910 ( 
.A1(n_13798),
.A2(n_13806),
.B1(n_13815),
.B2(n_13775),
.Y(n_13910)
);

INVx1_ASAP7_75t_L g13911 ( 
.A(n_13819),
.Y(n_13911)
);

AOI221xp5_ASAP7_75t_L g13912 ( 
.A1(n_13755),
.A2(n_2528),
.B1(n_2526),
.B2(n_2527),
.C(n_2530),
.Y(n_13912)
);

OAI21xp5_ASAP7_75t_L g13913 ( 
.A1(n_13792),
.A2(n_2526),
.B(n_2527),
.Y(n_13913)
);

NAND2xp5_ASAP7_75t_L g13914 ( 
.A(n_13862),
.B(n_2530),
.Y(n_13914)
);

AND2x2_ASAP7_75t_L g13915 ( 
.A(n_13828),
.B(n_2528),
.Y(n_13915)
);

AOI211xp5_ASAP7_75t_L g13916 ( 
.A1(n_13844),
.A2(n_2533),
.B(n_2531),
.C(n_2532),
.Y(n_13916)
);

OAI211xp5_ASAP7_75t_SL g13917 ( 
.A1(n_13831),
.A2(n_3462),
.B(n_3463),
.C(n_3461),
.Y(n_13917)
);

NAND2xp5_ASAP7_75t_L g13918 ( 
.A(n_13783),
.B(n_2533),
.Y(n_13918)
);

AOI22xp33_ASAP7_75t_L g13919 ( 
.A1(n_13843),
.A2(n_13794),
.B1(n_13788),
.B2(n_13773),
.Y(n_13919)
);

OAI22xp5_ASAP7_75t_L g13920 ( 
.A1(n_13863),
.A2(n_2535),
.B1(n_2532),
.B2(n_2534),
.Y(n_13920)
);

AOI31xp33_ASAP7_75t_L g13921 ( 
.A1(n_13812),
.A2(n_2536),
.A3(n_2534),
.B(n_2535),
.Y(n_13921)
);

AOI21xp33_ASAP7_75t_L g13922 ( 
.A1(n_13833),
.A2(n_2536),
.B(n_2538),
.Y(n_13922)
);

INVx1_ASAP7_75t_L g13923 ( 
.A(n_13762),
.Y(n_13923)
);

AOI21xp5_ASAP7_75t_L g13924 ( 
.A1(n_13826),
.A2(n_2539),
.B(n_2540),
.Y(n_13924)
);

INVx1_ASAP7_75t_L g13925 ( 
.A(n_13781),
.Y(n_13925)
);

AOI221x1_ASAP7_75t_L g13926 ( 
.A1(n_13802),
.A2(n_2542),
.B1(n_2539),
.B2(n_2541),
.C(n_2544),
.Y(n_13926)
);

AOI221xp5_ASAP7_75t_L g13927 ( 
.A1(n_13804),
.A2(n_13803),
.B1(n_13838),
.B2(n_13821),
.C(n_13782),
.Y(n_13927)
);

OAI22xp33_ASAP7_75t_L g13928 ( 
.A1(n_13766),
.A2(n_2544),
.B1(n_2545),
.B2(n_2542),
.Y(n_13928)
);

OAI211xp5_ASAP7_75t_L g13929 ( 
.A1(n_13855),
.A2(n_2546),
.B(n_2541),
.C(n_2545),
.Y(n_13929)
);

AOI221xp5_ASAP7_75t_L g13930 ( 
.A1(n_13787),
.A2(n_2548),
.B1(n_2546),
.B2(n_2547),
.C(n_2549),
.Y(n_13930)
);

OAI221xp5_ASAP7_75t_L g13931 ( 
.A1(n_13845),
.A2(n_2552),
.B1(n_2548),
.B2(n_2550),
.C(n_2553),
.Y(n_13931)
);

OAI22xp5_ASAP7_75t_L g13932 ( 
.A1(n_13784),
.A2(n_2555),
.B1(n_2552),
.B2(n_2554),
.Y(n_13932)
);

AOI211xp5_ASAP7_75t_L g13933 ( 
.A1(n_13837),
.A2(n_2556),
.B(n_2554),
.C(n_2555),
.Y(n_13933)
);

OAI31xp33_ASAP7_75t_L g13934 ( 
.A1(n_13811),
.A2(n_2559),
.A3(n_2557),
.B(n_2558),
.Y(n_13934)
);

INVx2_ASAP7_75t_L g13935 ( 
.A(n_13754),
.Y(n_13935)
);

AOI221x1_ASAP7_75t_L g13936 ( 
.A1(n_13752),
.A2(n_2559),
.B1(n_2557),
.B2(n_2558),
.C(n_2560),
.Y(n_13936)
);

OR2x2_ASAP7_75t_L g13937 ( 
.A(n_13774),
.B(n_2560),
.Y(n_13937)
);

OAI21xp33_ASAP7_75t_SL g13938 ( 
.A1(n_13813),
.A2(n_2561),
.B(n_2562),
.Y(n_13938)
);

NAND2xp5_ASAP7_75t_L g13939 ( 
.A(n_13799),
.B(n_2562),
.Y(n_13939)
);

INVxp67_ASAP7_75t_L g13940 ( 
.A(n_13744),
.Y(n_13940)
);

AO22x1_ASAP7_75t_L g13941 ( 
.A1(n_13851),
.A2(n_2564),
.B1(n_2561),
.B2(n_2563),
.Y(n_13941)
);

AOI22xp5_ASAP7_75t_L g13942 ( 
.A1(n_13795),
.A2(n_2566),
.B1(n_2564),
.B2(n_2565),
.Y(n_13942)
);

OAI211xp5_ASAP7_75t_L g13943 ( 
.A1(n_13738),
.A2(n_2568),
.B(n_2565),
.C(n_2567),
.Y(n_13943)
);

OAI221xp5_ASAP7_75t_SL g13944 ( 
.A1(n_13825),
.A2(n_2570),
.B1(n_2567),
.B2(n_2568),
.C(n_2571),
.Y(n_13944)
);

AND2x2_ASAP7_75t_L g13945 ( 
.A(n_13793),
.B(n_2570),
.Y(n_13945)
);

NOR3xp33_ASAP7_75t_L g13946 ( 
.A(n_13801),
.B(n_2573),
.C(n_2572),
.Y(n_13946)
);

O2A1O1Ixp5_ASAP7_75t_L g13947 ( 
.A1(n_13817),
.A2(n_2574),
.B(n_2571),
.C(n_2572),
.Y(n_13947)
);

OAI221xp5_ASAP7_75t_L g13948 ( 
.A1(n_13827),
.A2(n_2576),
.B1(n_2574),
.B2(n_2575),
.C(n_2577),
.Y(n_13948)
);

OAI22xp5_ASAP7_75t_L g13949 ( 
.A1(n_13800),
.A2(n_13810),
.B1(n_13739),
.B2(n_13751),
.Y(n_13949)
);

OAI32xp33_ASAP7_75t_L g13950 ( 
.A1(n_13834),
.A2(n_2577),
.A3(n_2575),
.B1(n_2576),
.B2(n_2578),
.Y(n_13950)
);

NOR2xp33_ASAP7_75t_L g13951 ( 
.A(n_13858),
.B(n_2579),
.Y(n_13951)
);

INVx1_ASAP7_75t_L g13952 ( 
.A(n_13818),
.Y(n_13952)
);

OAI221xp5_ASAP7_75t_L g13953 ( 
.A1(n_13835),
.A2(n_2582),
.B1(n_2580),
.B2(n_2581),
.C(n_2583),
.Y(n_13953)
);

OAI22xp5_ASAP7_75t_L g13954 ( 
.A1(n_13770),
.A2(n_2582),
.B1(n_2580),
.B2(n_2581),
.Y(n_13954)
);

AOI221xp5_ASAP7_75t_L g13955 ( 
.A1(n_13808),
.A2(n_2585),
.B1(n_2583),
.B2(n_2584),
.C(n_2586),
.Y(n_13955)
);

AND3x1_ASAP7_75t_L g13956 ( 
.A(n_13737),
.B(n_2584),
.C(n_2585),
.Y(n_13956)
);

AOI31xp33_ASAP7_75t_L g13957 ( 
.A1(n_13859),
.A2(n_2588),
.A3(n_2586),
.B(n_2587),
.Y(n_13957)
);

NAND2xp33_ASAP7_75t_L g13958 ( 
.A(n_13859),
.B(n_2587),
.Y(n_13958)
);

OAI222xp33_ASAP7_75t_L g13959 ( 
.A1(n_13736),
.A2(n_2615),
.B1(n_2598),
.B2(n_2624),
.C1(n_2606),
.C2(n_2589),
.Y(n_13959)
);

AOI221xp5_ASAP7_75t_L g13960 ( 
.A1(n_13786),
.A2(n_2591),
.B1(n_2589),
.B2(n_2590),
.C(n_2592),
.Y(n_13960)
);

OAI22xp5_ASAP7_75t_L g13961 ( 
.A1(n_13736),
.A2(n_2594),
.B1(n_2590),
.B2(n_2592),
.Y(n_13961)
);

AOI21xp5_ASAP7_75t_L g13962 ( 
.A1(n_13763),
.A2(n_2594),
.B(n_2595),
.Y(n_13962)
);

NOR4xp25_ASAP7_75t_SL g13963 ( 
.A(n_13839),
.B(n_2597),
.C(n_2595),
.D(n_2596),
.Y(n_13963)
);

OAI31xp33_ASAP7_75t_L g13964 ( 
.A1(n_13839),
.A2(n_2599),
.A3(n_2596),
.B(n_2598),
.Y(n_13964)
);

AOI221xp5_ASAP7_75t_L g13965 ( 
.A1(n_13786),
.A2(n_2601),
.B1(n_2599),
.B2(n_2600),
.C(n_2602),
.Y(n_13965)
);

OAI21xp5_ASAP7_75t_L g13966 ( 
.A1(n_13736),
.A2(n_2600),
.B(n_2601),
.Y(n_13966)
);

OAI221xp5_ASAP7_75t_L g13967 ( 
.A1(n_13736),
.A2(n_2604),
.B1(n_2602),
.B2(n_2603),
.C(n_2605),
.Y(n_13967)
);

XOR2xp5_ASAP7_75t_L g13968 ( 
.A(n_13736),
.B(n_3451),
.Y(n_13968)
);

INVx1_ASAP7_75t_L g13969 ( 
.A(n_13791),
.Y(n_13969)
);

AOI221x1_ASAP7_75t_L g13970 ( 
.A1(n_13737),
.A2(n_2608),
.B1(n_2606),
.B2(n_2607),
.C(n_2609),
.Y(n_13970)
);

NAND2xp5_ASAP7_75t_L g13971 ( 
.A(n_13750),
.B(n_2608),
.Y(n_13971)
);

OAI31xp33_ASAP7_75t_L g13972 ( 
.A1(n_13839),
.A2(n_2610),
.A3(n_2607),
.B(n_2609),
.Y(n_13972)
);

INVx3_ASAP7_75t_L g13973 ( 
.A(n_13750),
.Y(n_13973)
);

INVx1_ASAP7_75t_L g13974 ( 
.A(n_13915),
.Y(n_13974)
);

AOI22xp5_ASAP7_75t_L g13975 ( 
.A1(n_13973),
.A2(n_2620),
.B1(n_2628),
.B2(n_2610),
.Y(n_13975)
);

NAND3xp33_ASAP7_75t_SL g13976 ( 
.A(n_13963),
.B(n_2611),
.C(n_2613),
.Y(n_13976)
);

O2A1O1Ixp5_ASAP7_75t_L g13977 ( 
.A1(n_13909),
.A2(n_2615),
.B(n_2611),
.C(n_2614),
.Y(n_13977)
);

O2A1O1Ixp33_ASAP7_75t_L g13978 ( 
.A1(n_13958),
.A2(n_2619),
.B(n_2616),
.C(n_2617),
.Y(n_13978)
);

AOI22xp5_ASAP7_75t_L g13979 ( 
.A1(n_13973),
.A2(n_13895),
.B1(n_13900),
.B2(n_13951),
.Y(n_13979)
);

AOI211xp5_ASAP7_75t_L g13980 ( 
.A1(n_13876),
.A2(n_2621),
.B(n_2617),
.C(n_2620),
.Y(n_13980)
);

NAND3xp33_ASAP7_75t_SL g13981 ( 
.A(n_13964),
.B(n_2621),
.C(n_2622),
.Y(n_13981)
);

NOR2xp33_ASAP7_75t_L g13982 ( 
.A(n_13917),
.B(n_2622),
.Y(n_13982)
);

OAI211xp5_ASAP7_75t_L g13983 ( 
.A1(n_13938),
.A2(n_2625),
.B(n_2623),
.C(n_2624),
.Y(n_13983)
);

OAI21xp5_ASAP7_75t_SL g13984 ( 
.A1(n_13907),
.A2(n_2626),
.B(n_2625),
.Y(n_13984)
);

NAND2xp5_ASAP7_75t_L g13985 ( 
.A(n_13941),
.B(n_2623),
.Y(n_13985)
);

AOI22xp5_ASAP7_75t_L g13986 ( 
.A1(n_13968),
.A2(n_2634),
.B1(n_2643),
.B2(n_2626),
.Y(n_13986)
);

NOR2xp33_ASAP7_75t_L g13987 ( 
.A(n_13904),
.B(n_2627),
.Y(n_13987)
);

AOI222xp33_ASAP7_75t_L g13988 ( 
.A1(n_13866),
.A2(n_2629),
.B1(n_2631),
.B2(n_2627),
.C1(n_2628),
.C2(n_2630),
.Y(n_13988)
);

OAI21xp33_ASAP7_75t_L g13989 ( 
.A1(n_13878),
.A2(n_2629),
.B(n_2630),
.Y(n_13989)
);

AOI222xp33_ASAP7_75t_L g13990 ( 
.A1(n_13971),
.A2(n_2633),
.B1(n_2636),
.B2(n_2631),
.C1(n_2632),
.C2(n_2635),
.Y(n_13990)
);

AOI221x1_ASAP7_75t_L g13991 ( 
.A1(n_13877),
.A2(n_13966),
.B1(n_13962),
.B2(n_13901),
.C(n_13879),
.Y(n_13991)
);

AOI211x1_ASAP7_75t_L g13992 ( 
.A1(n_13873),
.A2(n_2638),
.B(n_2632),
.C(n_2637),
.Y(n_13992)
);

INVx1_ASAP7_75t_L g13993 ( 
.A(n_13865),
.Y(n_13993)
);

OAI211xp5_ASAP7_75t_L g13994 ( 
.A1(n_13884),
.A2(n_2640),
.B(n_2637),
.C(n_2639),
.Y(n_13994)
);

AOI211xp5_ASAP7_75t_L g13995 ( 
.A1(n_13928),
.A2(n_13950),
.B(n_13943),
.C(n_13929),
.Y(n_13995)
);

AOI21xp5_ASAP7_75t_L g13996 ( 
.A1(n_13870),
.A2(n_2649),
.B(n_2639),
.Y(n_13996)
);

NAND3xp33_ASAP7_75t_L g13997 ( 
.A(n_13908),
.B(n_2641),
.C(n_2643),
.Y(n_13997)
);

AOI21xp5_ASAP7_75t_L g13998 ( 
.A1(n_13914),
.A2(n_2651),
.B(n_2641),
.Y(n_13998)
);

NAND2xp5_ASAP7_75t_L g13999 ( 
.A(n_13945),
.B(n_2644),
.Y(n_13999)
);

OAI211xp5_ASAP7_75t_L g14000 ( 
.A1(n_13972),
.A2(n_2646),
.B(n_2644),
.C(n_2645),
.Y(n_14000)
);

NAND2xp5_ASAP7_75t_L g14001 ( 
.A(n_13891),
.B(n_2645),
.Y(n_14001)
);

AOI211x1_ASAP7_75t_L g14002 ( 
.A1(n_13913),
.A2(n_2648),
.B(n_2646),
.C(n_2647),
.Y(n_14002)
);

INVx1_ASAP7_75t_SL g14003 ( 
.A(n_13890),
.Y(n_14003)
);

INVx1_ASAP7_75t_L g14004 ( 
.A(n_13903),
.Y(n_14004)
);

O2A1O1Ixp33_ASAP7_75t_SL g14005 ( 
.A1(n_13906),
.A2(n_2649),
.B(n_2647),
.C(n_2648),
.Y(n_14005)
);

AOI21xp5_ASAP7_75t_L g14006 ( 
.A1(n_13897),
.A2(n_13899),
.B(n_13924),
.Y(n_14006)
);

INVx2_ASAP7_75t_SL g14007 ( 
.A(n_13937),
.Y(n_14007)
);

AOI21xp5_ASAP7_75t_L g14008 ( 
.A1(n_13918),
.A2(n_2659),
.B(n_2650),
.Y(n_14008)
);

OAI221xp5_ASAP7_75t_L g14009 ( 
.A1(n_13919),
.A2(n_2668),
.B1(n_2677),
.B2(n_2660),
.C(n_2651),
.Y(n_14009)
);

AOI22xp33_ASAP7_75t_L g14010 ( 
.A1(n_13886),
.A2(n_2654),
.B1(n_2652),
.B2(n_2653),
.Y(n_14010)
);

AOI22xp5_ASAP7_75t_L g14011 ( 
.A1(n_13892),
.A2(n_2662),
.B1(n_2672),
.B2(n_2652),
.Y(n_14011)
);

INVx1_ASAP7_75t_L g14012 ( 
.A(n_13898),
.Y(n_14012)
);

OR2x2_ASAP7_75t_L g14013 ( 
.A(n_13868),
.B(n_13880),
.Y(n_14013)
);

NAND2xp5_ASAP7_75t_L g14014 ( 
.A(n_13957),
.B(n_2653),
.Y(n_14014)
);

AOI22xp5_ASAP7_75t_L g14015 ( 
.A1(n_13956),
.A2(n_2664),
.B1(n_2675),
.B2(n_2654),
.Y(n_14015)
);

NOR2xp33_ASAP7_75t_L g14016 ( 
.A(n_13921),
.B(n_2655),
.Y(n_14016)
);

INVx1_ASAP7_75t_L g14017 ( 
.A(n_13905),
.Y(n_14017)
);

INVx1_ASAP7_75t_L g14018 ( 
.A(n_13872),
.Y(n_14018)
);

NAND3xp33_ASAP7_75t_L g14019 ( 
.A(n_13916),
.B(n_2655),
.C(n_2656),
.Y(n_14019)
);

AOI21xp5_ASAP7_75t_L g14020 ( 
.A1(n_13867),
.A2(n_2667),
.B(n_2656),
.Y(n_14020)
);

NAND2xp5_ASAP7_75t_SL g14021 ( 
.A(n_13887),
.B(n_2658),
.Y(n_14021)
);

NAND3xp33_ASAP7_75t_L g14022 ( 
.A(n_13912),
.B(n_2658),
.C(n_2659),
.Y(n_14022)
);

AOI21xp5_ASAP7_75t_L g14023 ( 
.A1(n_13939),
.A2(n_2673),
.B(n_2661),
.Y(n_14023)
);

AOI211xp5_ASAP7_75t_L g14024 ( 
.A1(n_13922),
.A2(n_13931),
.B(n_13875),
.C(n_13949),
.Y(n_14024)
);

AOI21xp5_ASAP7_75t_L g14025 ( 
.A1(n_13940),
.A2(n_2673),
.B(n_2661),
.Y(n_14025)
);

A2O1A1Ixp33_ASAP7_75t_L g14026 ( 
.A1(n_13947),
.A2(n_13934),
.B(n_13965),
.C(n_13960),
.Y(n_14026)
);

AOI211xp5_ASAP7_75t_L g14027 ( 
.A1(n_13910),
.A2(n_2665),
.B(n_2662),
.C(n_2663),
.Y(n_14027)
);

AOI21xp5_ASAP7_75t_L g14028 ( 
.A1(n_13967),
.A2(n_13953),
.B(n_13948),
.Y(n_14028)
);

AND2x2_ASAP7_75t_L g14029 ( 
.A(n_13894),
.B(n_2663),
.Y(n_14029)
);

AOI21xp5_ASAP7_75t_L g14030 ( 
.A1(n_13954),
.A2(n_2677),
.B(n_2665),
.Y(n_14030)
);

AOI221xp5_ASAP7_75t_L g14031 ( 
.A1(n_13927),
.A2(n_2669),
.B1(n_2674),
.B2(n_2667),
.C(n_2670),
.Y(n_14031)
);

AOI22xp5_ASAP7_75t_L g14032 ( 
.A1(n_13969),
.A2(n_13871),
.B1(n_13911),
.B2(n_13952),
.Y(n_14032)
);

AOI322xp5_ASAP7_75t_L g14033 ( 
.A1(n_13883),
.A2(n_2678),
.A3(n_2676),
.B1(n_2674),
.B2(n_2666),
.C1(n_2669),
.C2(n_2675),
.Y(n_14033)
);

OAI22xp5_ASAP7_75t_L g14034 ( 
.A1(n_13933),
.A2(n_2679),
.B1(n_2666),
.B2(n_2676),
.Y(n_14034)
);

OAI211xp5_ASAP7_75t_L g14035 ( 
.A1(n_13970),
.A2(n_2681),
.B(n_2679),
.C(n_2680),
.Y(n_14035)
);

OAI22xp5_ASAP7_75t_L g14036 ( 
.A1(n_13869),
.A2(n_2683),
.B1(n_2681),
.B2(n_2682),
.Y(n_14036)
);

NOR4xp25_ASAP7_75t_L g14037 ( 
.A(n_13888),
.B(n_2685),
.C(n_2683),
.D(n_2684),
.Y(n_14037)
);

OAI21xp33_ASAP7_75t_SL g14038 ( 
.A1(n_13902),
.A2(n_2692),
.B(n_2684),
.Y(n_14038)
);

AOI211x1_ASAP7_75t_L g14039 ( 
.A1(n_13959),
.A2(n_2687),
.B(n_2685),
.C(n_2686),
.Y(n_14039)
);

NAND4xp25_ASAP7_75t_L g14040 ( 
.A(n_13926),
.B(n_2695),
.C(n_2704),
.D(n_2687),
.Y(n_14040)
);

NAND2xp33_ASAP7_75t_L g14041 ( 
.A(n_13946),
.B(n_2688),
.Y(n_14041)
);

AOI22xp5_ASAP7_75t_L g14042 ( 
.A1(n_13874),
.A2(n_2698),
.B1(n_2709),
.B2(n_2689),
.Y(n_14042)
);

OAI22xp33_ASAP7_75t_L g14043 ( 
.A1(n_13936),
.A2(n_2691),
.B1(n_2689),
.B2(n_2690),
.Y(n_14043)
);

AND2x2_ASAP7_75t_L g14044 ( 
.A(n_13893),
.B(n_13935),
.Y(n_14044)
);

NAND3xp33_ASAP7_75t_SL g14045 ( 
.A(n_13955),
.B(n_2690),
.C(n_2692),
.Y(n_14045)
);

AOI211xp5_ASAP7_75t_L g14046 ( 
.A1(n_13882),
.A2(n_2695),
.B(n_2693),
.C(n_2694),
.Y(n_14046)
);

AOI221xp5_ASAP7_75t_L g14047 ( 
.A1(n_13881),
.A2(n_2698),
.B1(n_2700),
.B2(n_2696),
.C(n_2699),
.Y(n_14047)
);

AOI221xp5_ASAP7_75t_L g14048 ( 
.A1(n_13961),
.A2(n_2700),
.B1(n_2702),
.B2(n_2696),
.C(n_2701),
.Y(n_14048)
);

AOI222xp33_ASAP7_75t_L g14049 ( 
.A1(n_13923),
.A2(n_13925),
.B1(n_13930),
.B2(n_13932),
.C1(n_13920),
.C2(n_13944),
.Y(n_14049)
);

AOI321xp33_ASAP7_75t_L g14050 ( 
.A1(n_13885),
.A2(n_2703),
.A3(n_2708),
.B1(n_2694),
.B2(n_2701),
.C(n_2706),
.Y(n_14050)
);

AOI221xp5_ASAP7_75t_L g14051 ( 
.A1(n_13942),
.A2(n_2709),
.B1(n_2711),
.B2(n_2706),
.C(n_2710),
.Y(n_14051)
);

A2O1A1Ixp33_ASAP7_75t_L g14052 ( 
.A1(n_13889),
.A2(n_2712),
.B(n_2703),
.C(n_2711),
.Y(n_14052)
);

NAND2xp5_ASAP7_75t_L g14053 ( 
.A(n_13896),
.B(n_2712),
.Y(n_14053)
);

OAI221xp5_ASAP7_75t_SL g14054 ( 
.A1(n_13878),
.A2(n_2715),
.B1(n_2713),
.B2(n_2714),
.C(n_2716),
.Y(n_14054)
);

AOI22xp5_ASAP7_75t_L g14055 ( 
.A1(n_13973),
.A2(n_2721),
.B1(n_2730),
.B2(n_2713),
.Y(n_14055)
);

NAND2xp5_ASAP7_75t_L g14056 ( 
.A(n_13941),
.B(n_2714),
.Y(n_14056)
);

HB1xp67_ASAP7_75t_L g14057 ( 
.A(n_13973),
.Y(n_14057)
);

OAI221xp5_ASAP7_75t_L g14058 ( 
.A1(n_13964),
.A2(n_2732),
.B1(n_2740),
.B2(n_2723),
.C(n_2715),
.Y(n_14058)
);

OAI221xp5_ASAP7_75t_L g14059 ( 
.A1(n_13964),
.A2(n_2733),
.B1(n_2741),
.B2(n_2724),
.C(n_2716),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13915),
.Y(n_14060)
);

INVxp67_ASAP7_75t_L g14061 ( 
.A(n_13905),
.Y(n_14061)
);

NAND2xp33_ASAP7_75t_L g14062 ( 
.A(n_13887),
.B(n_2717),
.Y(n_14062)
);

AND2x2_ASAP7_75t_L g14063 ( 
.A(n_13973),
.B(n_2717),
.Y(n_14063)
);

OAI22xp33_ASAP7_75t_L g14064 ( 
.A1(n_13908),
.A2(n_2720),
.B1(n_2718),
.B2(n_2719),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_L g14065 ( 
.A(n_14063),
.B(n_2718),
.Y(n_14065)
);

NOR2xp33_ASAP7_75t_R g14066 ( 
.A(n_13976),
.B(n_3461),
.Y(n_14066)
);

NAND2xp5_ASAP7_75t_L g14067 ( 
.A(n_14057),
.B(n_14064),
.Y(n_14067)
);

NOR4xp25_ASAP7_75t_L g14068 ( 
.A(n_13989),
.B(n_3462),
.C(n_2722),
.D(n_2719),
.Y(n_14068)
);

NOR3xp33_ASAP7_75t_L g14069 ( 
.A(n_14054),
.B(n_2721),
.C(n_2722),
.Y(n_14069)
);

AOI211x1_ASAP7_75t_SL g14070 ( 
.A1(n_13997),
.A2(n_2725),
.B(n_2723),
.C(n_2724),
.Y(n_14070)
);

OAI21xp5_ASAP7_75t_SL g14071 ( 
.A1(n_13979),
.A2(n_2725),
.B(n_2726),
.Y(n_14071)
);

NOR3xp33_ASAP7_75t_L g14072 ( 
.A(n_14038),
.B(n_2726),
.C(n_2727),
.Y(n_14072)
);

OAI22xp33_ASAP7_75t_L g14073 ( 
.A1(n_14011),
.A2(n_2731),
.B1(n_2728),
.B2(n_2730),
.Y(n_14073)
);

OAI211xp5_ASAP7_75t_L g14074 ( 
.A1(n_13980),
.A2(n_2734),
.B(n_2731),
.C(n_2732),
.Y(n_14074)
);

NAND3xp33_ASAP7_75t_SL g14075 ( 
.A(n_14046),
.B(n_2734),
.C(n_2735),
.Y(n_14075)
);

AOI21xp5_ASAP7_75t_L g14076 ( 
.A1(n_14041),
.A2(n_2735),
.B(n_2736),
.Y(n_14076)
);

NOR4xp25_ASAP7_75t_L g14077 ( 
.A(n_13981),
.B(n_3459),
.C(n_2738),
.D(n_2736),
.Y(n_14077)
);

NOR2xp33_ASAP7_75t_L g14078 ( 
.A(n_14000),
.B(n_2737),
.Y(n_14078)
);

AOI211xp5_ASAP7_75t_L g14079 ( 
.A1(n_14043),
.A2(n_2739),
.B(n_2737),
.C(n_2738),
.Y(n_14079)
);

AOI21xp5_ASAP7_75t_L g14080 ( 
.A1(n_14062),
.A2(n_2740),
.B(n_2741),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_14037),
.B(n_2742),
.Y(n_14081)
);

NOR3xp33_ASAP7_75t_L g14082 ( 
.A(n_14009),
.B(n_2743),
.C(n_2744),
.Y(n_14082)
);

NOR3xp33_ASAP7_75t_SL g14083 ( 
.A(n_14045),
.B(n_2743),
.C(n_2744),
.Y(n_14083)
);

AOI21xp5_ASAP7_75t_L g14084 ( 
.A1(n_14021),
.A2(n_14008),
.B(n_13998),
.Y(n_14084)
);

NAND3xp33_ASAP7_75t_SL g14085 ( 
.A(n_14015),
.B(n_2745),
.C(n_2746),
.Y(n_14085)
);

AOI221xp5_ASAP7_75t_L g14086 ( 
.A1(n_13992),
.A2(n_2749),
.B1(n_2745),
.B2(n_2747),
.C(n_2750),
.Y(n_14086)
);

OAI22xp5_ASAP7_75t_L g14087 ( 
.A1(n_14032),
.A2(n_2758),
.B1(n_2766),
.B2(n_2747),
.Y(n_14087)
);

OAI221xp5_ASAP7_75t_L g14088 ( 
.A1(n_13984),
.A2(n_3458),
.B1(n_3459),
.B2(n_3457),
.C(n_3456),
.Y(n_14088)
);

AOI222xp33_ASAP7_75t_L g14089 ( 
.A1(n_14018),
.A2(n_2753),
.B1(n_2755),
.B2(n_2750),
.C1(n_2751),
.C2(n_2754),
.Y(n_14089)
);

AOI22xp33_ASAP7_75t_L g14090 ( 
.A1(n_13987),
.A2(n_2757),
.B1(n_2754),
.B2(n_2756),
.Y(n_14090)
);

NAND4xp25_ASAP7_75t_L g14091 ( 
.A(n_14024),
.B(n_2758),
.C(n_2756),
.D(n_2757),
.Y(n_14091)
);

AOI22xp5_ASAP7_75t_L g14092 ( 
.A1(n_13982),
.A2(n_2761),
.B1(n_2759),
.B2(n_2760),
.Y(n_14092)
);

XOR2xp5_ASAP7_75t_L g14093 ( 
.A(n_14040),
.B(n_3450),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13985),
.Y(n_14094)
);

NAND2xp5_ASAP7_75t_L g14095 ( 
.A(n_14029),
.B(n_2759),
.Y(n_14095)
);

AOI221x1_ASAP7_75t_L g14096 ( 
.A1(n_14020),
.A2(n_2763),
.B1(n_2760),
.B2(n_2762),
.C(n_2764),
.Y(n_14096)
);

NAND3xp33_ASAP7_75t_SL g14097 ( 
.A(n_14047),
.B(n_2765),
.C(n_2766),
.Y(n_14097)
);

AOI221xp5_ASAP7_75t_L g14098 ( 
.A1(n_14005),
.A2(n_2768),
.B1(n_2765),
.B2(n_2767),
.C(n_2769),
.Y(n_14098)
);

NOR2xp33_ASAP7_75t_L g14099 ( 
.A(n_13983),
.B(n_2768),
.Y(n_14099)
);

OAI22xp5_ASAP7_75t_L g14100 ( 
.A1(n_14042),
.A2(n_2778),
.B1(n_2786),
.B2(n_2769),
.Y(n_14100)
);

AOI31xp33_ASAP7_75t_L g14101 ( 
.A1(n_14016),
.A2(n_2773),
.A3(n_2771),
.B(n_2772),
.Y(n_14101)
);

NOR2xp33_ASAP7_75t_L g14102 ( 
.A(n_14058),
.B(n_2772),
.Y(n_14102)
);

OAI221xp5_ASAP7_75t_L g14103 ( 
.A1(n_14035),
.A2(n_3449),
.B1(n_3450),
.B2(n_3448),
.C(n_3447),
.Y(n_14103)
);

OAI21xp33_ASAP7_75t_SL g14104 ( 
.A1(n_14056),
.A2(n_2774),
.B(n_2775),
.Y(n_14104)
);

OAI211xp5_ASAP7_75t_L g14105 ( 
.A1(n_13978),
.A2(n_2777),
.B(n_2774),
.C(n_2776),
.Y(n_14105)
);

OAI21xp5_ASAP7_75t_SL g14106 ( 
.A1(n_13994),
.A2(n_2777),
.B(n_2778),
.Y(n_14106)
);

NOR2x1_ASAP7_75t_L g14107 ( 
.A(n_13999),
.B(n_2780),
.Y(n_14107)
);

OAI211xp5_ASAP7_75t_SL g14108 ( 
.A1(n_14049),
.A2(n_2788),
.B(n_2797),
.C(n_2779),
.Y(n_14108)
);

INVx1_ASAP7_75t_SL g14109 ( 
.A(n_14014),
.Y(n_14109)
);

AOI221xp5_ASAP7_75t_L g14110 ( 
.A1(n_14039),
.A2(n_14002),
.B1(n_13977),
.B2(n_14019),
.C(n_14034),
.Y(n_14110)
);

AOI221xp5_ASAP7_75t_SL g14111 ( 
.A1(n_14028),
.A2(n_2782),
.B1(n_2779),
.B2(n_2781),
.C(n_2783),
.Y(n_14111)
);

NAND2xp5_ASAP7_75t_L g14112 ( 
.A(n_13988),
.B(n_2781),
.Y(n_14112)
);

OAI211xp5_ASAP7_75t_SL g14113 ( 
.A1(n_13995),
.A2(n_2793),
.B(n_2802),
.C(n_2783),
.Y(n_14113)
);

OAI221xp5_ASAP7_75t_L g14114 ( 
.A1(n_14059),
.A2(n_3465),
.B1(n_3464),
.B2(n_2786),
.C(n_2784),
.Y(n_14114)
);

AOI221xp5_ASAP7_75t_L g14115 ( 
.A1(n_14022),
.A2(n_2787),
.B1(n_2784),
.B2(n_2785),
.C(n_2789),
.Y(n_14115)
);

AOI21xp33_ASAP7_75t_L g14116 ( 
.A1(n_14001),
.A2(n_2785),
.B(n_2787),
.Y(n_14116)
);

NAND2xp5_ASAP7_75t_L g14117 ( 
.A(n_13990),
.B(n_2789),
.Y(n_14117)
);

OAI211xp5_ASAP7_75t_L g14118 ( 
.A1(n_13991),
.A2(n_2793),
.B(n_2790),
.C(n_2792),
.Y(n_14118)
);

AOI21xp5_ASAP7_75t_L g14119 ( 
.A1(n_13996),
.A2(n_2790),
.B(n_2792),
.Y(n_14119)
);

NAND2xp5_ASAP7_75t_L g14120 ( 
.A(n_14027),
.B(n_2794),
.Y(n_14120)
);

NAND2xp5_ASAP7_75t_L g14121 ( 
.A(n_14025),
.B(n_2794),
.Y(n_14121)
);

INVx1_ASAP7_75t_L g14122 ( 
.A(n_14044),
.Y(n_14122)
);

AOI22xp5_ASAP7_75t_L g14123 ( 
.A1(n_14003),
.A2(n_2798),
.B1(n_2795),
.B2(n_2796),
.Y(n_14123)
);

NAND2xp33_ASAP7_75t_SL g14124 ( 
.A(n_14007),
.B(n_2795),
.Y(n_14124)
);

OAI21xp33_ASAP7_75t_L g14125 ( 
.A1(n_13974),
.A2(n_2798),
.B(n_2799),
.Y(n_14125)
);

AOI221xp5_ASAP7_75t_L g14126 ( 
.A1(n_14030),
.A2(n_14026),
.B1(n_13993),
.B2(n_14006),
.C(n_14060),
.Y(n_14126)
);

NOR3xp33_ASAP7_75t_L g14127 ( 
.A(n_14061),
.B(n_2799),
.C(n_2800),
.Y(n_14127)
);

NAND2xp5_ASAP7_75t_L g14128 ( 
.A(n_13986),
.B(n_2800),
.Y(n_14128)
);

INVx1_ASAP7_75t_L g14129 ( 
.A(n_14053),
.Y(n_14129)
);

OAI221xp5_ASAP7_75t_L g14130 ( 
.A1(n_14050),
.A2(n_3464),
.B1(n_3460),
.B2(n_3458),
.C(n_2803),
.Y(n_14130)
);

OAI221xp5_ASAP7_75t_L g14131 ( 
.A1(n_14052),
.A2(n_2803),
.B1(n_2801),
.B2(n_2802),
.C(n_2804),
.Y(n_14131)
);

NAND2xp5_ASAP7_75t_L g14132 ( 
.A(n_14031),
.B(n_2801),
.Y(n_14132)
);

AOI22xp5_ASAP7_75t_L g14133 ( 
.A1(n_14017),
.A2(n_2806),
.B1(n_2804),
.B2(n_2805),
.Y(n_14133)
);

NOR2xp33_ASAP7_75t_L g14134 ( 
.A(n_14023),
.B(n_2805),
.Y(n_14134)
);

NOR2xp33_ASAP7_75t_L g14135 ( 
.A(n_14130),
.B(n_14013),
.Y(n_14135)
);

NAND3xp33_ASAP7_75t_L g14136 ( 
.A(n_14079),
.B(n_14048),
.C(n_14051),
.Y(n_14136)
);

NAND4xp25_ASAP7_75t_SL g14137 ( 
.A(n_14086),
.B(n_14004),
.C(n_14012),
.D(n_13975),
.Y(n_14137)
);

AND2x2_ASAP7_75t_L g14138 ( 
.A(n_14122),
.B(n_14055),
.Y(n_14138)
);

AOI22xp33_ASAP7_75t_L g14139 ( 
.A1(n_14072),
.A2(n_14036),
.B1(n_14010),
.B2(n_14033),
.Y(n_14139)
);

AOI211xp5_ASAP7_75t_L g14140 ( 
.A1(n_14118),
.A2(n_2808),
.B(n_2806),
.C(n_2807),
.Y(n_14140)
);

AND2x2_ASAP7_75t_L g14141 ( 
.A(n_14083),
.B(n_2809),
.Y(n_14141)
);

AND2x2_ASAP7_75t_L g14142 ( 
.A(n_14069),
.B(n_2810),
.Y(n_14142)
);

AOI22xp33_ASAP7_75t_L g14143 ( 
.A1(n_14082),
.A2(n_2812),
.B1(n_2810),
.B2(n_2811),
.Y(n_14143)
);

NAND3xp33_ASAP7_75t_SL g14144 ( 
.A(n_14066),
.B(n_14070),
.C(n_14098),
.Y(n_14144)
);

NAND2xp5_ASAP7_75t_L g14145 ( 
.A(n_14101),
.B(n_2811),
.Y(n_14145)
);

INVx1_ASAP7_75t_L g14146 ( 
.A(n_14081),
.Y(n_14146)
);

NOR4xp25_ASAP7_75t_L g14147 ( 
.A(n_14071),
.B(n_2814),
.C(n_2812),
.D(n_2813),
.Y(n_14147)
);

AOI311xp33_ASAP7_75t_L g14148 ( 
.A1(n_14084),
.A2(n_14126),
.A3(n_14110),
.B(n_14094),
.C(n_14067),
.Y(n_14148)
);

NOR2x1_ASAP7_75t_L g14149 ( 
.A(n_14107),
.B(n_2813),
.Y(n_14149)
);

AND2x2_ASAP7_75t_L g14150 ( 
.A(n_14077),
.B(n_2814),
.Y(n_14150)
);

NAND2xp5_ASAP7_75t_L g14151 ( 
.A(n_14111),
.B(n_14127),
.Y(n_14151)
);

NOR3xp33_ASAP7_75t_L g14152 ( 
.A(n_14116),
.B(n_3456),
.C(n_2815),
.Y(n_14152)
);

INVx1_ASAP7_75t_L g14153 ( 
.A(n_14065),
.Y(n_14153)
);

NAND2xp5_ASAP7_75t_L g14154 ( 
.A(n_14125),
.B(n_2816),
.Y(n_14154)
);

NOR2xp33_ASAP7_75t_L g14155 ( 
.A(n_14108),
.B(n_14113),
.Y(n_14155)
);

NAND3xp33_ASAP7_75t_SL g14156 ( 
.A(n_14090),
.B(n_2816),
.C(n_2817),
.Y(n_14156)
);

NAND3xp33_ASAP7_75t_SL g14157 ( 
.A(n_14068),
.B(n_2817),
.C(n_2818),
.Y(n_14157)
);

NAND3xp33_ASAP7_75t_SL g14158 ( 
.A(n_14080),
.B(n_2819),
.C(n_2820),
.Y(n_14158)
);

NOR2x1_ASAP7_75t_L g14159 ( 
.A(n_14091),
.B(n_2819),
.Y(n_14159)
);

AND4x1_ASAP7_75t_L g14160 ( 
.A(n_14099),
.B(n_2829),
.C(n_2837),
.D(n_2821),
.Y(n_14160)
);

INVx1_ASAP7_75t_L g14161 ( 
.A(n_14093),
.Y(n_14161)
);

INVx1_ASAP7_75t_L g14162 ( 
.A(n_14095),
.Y(n_14162)
);

NAND3xp33_ASAP7_75t_SL g14163 ( 
.A(n_14115),
.B(n_2821),
.C(n_2822),
.Y(n_14163)
);

INVx1_ASAP7_75t_L g14164 ( 
.A(n_14121),
.Y(n_14164)
);

INVx1_ASAP7_75t_SL g14165 ( 
.A(n_14124),
.Y(n_14165)
);

INVx1_ASAP7_75t_L g14166 ( 
.A(n_14120),
.Y(n_14166)
);

INVx1_ASAP7_75t_L g14167 ( 
.A(n_14078),
.Y(n_14167)
);

NAND4xp25_ASAP7_75t_L g14168 ( 
.A(n_14102),
.B(n_2824),
.C(n_2822),
.D(n_2823),
.Y(n_14168)
);

NOR3xp33_ASAP7_75t_L g14169 ( 
.A(n_14104),
.B(n_3451),
.C(n_3449),
.Y(n_14169)
);

INVx1_ASAP7_75t_L g14170 ( 
.A(n_14103),
.Y(n_14170)
);

NAND2xp5_ASAP7_75t_SL g14171 ( 
.A(n_14073),
.B(n_2823),
.Y(n_14171)
);

NAND2x1_ASAP7_75t_L g14172 ( 
.A(n_14134),
.B(n_2824),
.Y(n_14172)
);

NAND2xp5_ASAP7_75t_L g14173 ( 
.A(n_14087),
.B(n_2825),
.Y(n_14173)
);

AOI221xp5_ASAP7_75t_L g14174 ( 
.A1(n_14075),
.A2(n_2827),
.B1(n_2825),
.B2(n_2826),
.C(n_2828),
.Y(n_14174)
);

NAND2xp5_ASAP7_75t_L g14175 ( 
.A(n_14096),
.B(n_2827),
.Y(n_14175)
);

NOR3xp33_ASAP7_75t_L g14176 ( 
.A(n_14112),
.B(n_2828),
.C(n_2829),
.Y(n_14176)
);

HB1xp67_ASAP7_75t_L g14177 ( 
.A(n_14100),
.Y(n_14177)
);

AOI311xp33_ASAP7_75t_L g14178 ( 
.A1(n_14129),
.A2(n_2832),
.A3(n_2830),
.B(n_2831),
.C(n_2833),
.Y(n_14178)
);

NAND2xp5_ASAP7_75t_L g14179 ( 
.A(n_14106),
.B(n_2830),
.Y(n_14179)
);

NOR2xp33_ASAP7_75t_L g14180 ( 
.A(n_14088),
.B(n_2831),
.Y(n_14180)
);

NAND2xp5_ASAP7_75t_L g14181 ( 
.A(n_14076),
.B(n_2832),
.Y(n_14181)
);

INVx1_ASAP7_75t_L g14182 ( 
.A(n_14117),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_14092),
.B(n_2833),
.Y(n_14183)
);

NAND2xp5_ASAP7_75t_L g14184 ( 
.A(n_14119),
.B(n_14089),
.Y(n_14184)
);

INVx1_ASAP7_75t_L g14185 ( 
.A(n_14128),
.Y(n_14185)
);

AOI211xp5_ASAP7_75t_L g14186 ( 
.A1(n_14074),
.A2(n_2836),
.B(n_2834),
.C(n_2835),
.Y(n_14186)
);

INVx2_ASAP7_75t_SL g14187 ( 
.A(n_14109),
.Y(n_14187)
);

INVx1_ASAP7_75t_L g14188 ( 
.A(n_14132),
.Y(n_14188)
);

NAND4xp25_ASAP7_75t_L g14189 ( 
.A(n_14097),
.B(n_2836),
.C(n_2834),
.D(n_2835),
.Y(n_14189)
);

NOR3xp33_ASAP7_75t_L g14190 ( 
.A(n_14114),
.B(n_14085),
.C(n_14105),
.Y(n_14190)
);

INVx1_ASAP7_75t_L g14191 ( 
.A(n_14131),
.Y(n_14191)
);

AOI221xp5_ASAP7_75t_L g14192 ( 
.A1(n_14123),
.A2(n_2840),
.B1(n_2838),
.B2(n_2839),
.C(n_2841),
.Y(n_14192)
);

NAND2xp33_ASAP7_75t_SL g14193 ( 
.A(n_14133),
.B(n_3447),
.Y(n_14193)
);

NOR2xp33_ASAP7_75t_L g14194 ( 
.A(n_14130),
.B(n_2839),
.Y(n_14194)
);

NAND3xp33_ASAP7_75t_L g14195 ( 
.A(n_14079),
.B(n_2840),
.C(n_2841),
.Y(n_14195)
);

AOI21xp5_ASAP7_75t_L g14196 ( 
.A1(n_14067),
.A2(n_2842),
.B(n_2843),
.Y(n_14196)
);

AND2x2_ASAP7_75t_L g14197 ( 
.A(n_14122),
.B(n_2842),
.Y(n_14197)
);

INVx2_ASAP7_75t_L g14198 ( 
.A(n_14122),
.Y(n_14198)
);

INVx1_ASAP7_75t_L g14199 ( 
.A(n_14081),
.Y(n_14199)
);

NAND2xp5_ASAP7_75t_L g14200 ( 
.A(n_14101),
.B(n_2843),
.Y(n_14200)
);

NOR3xp33_ASAP7_75t_L g14201 ( 
.A(n_14122),
.B(n_2844),
.C(n_2845),
.Y(n_14201)
);

AOI222xp33_ASAP7_75t_L g14202 ( 
.A1(n_14075),
.A2(n_2846),
.B1(n_2848),
.B2(n_2849),
.C1(n_2845),
.C2(n_2847),
.Y(n_14202)
);

NAND2xp33_ASAP7_75t_L g14203 ( 
.A(n_14072),
.B(n_2844),
.Y(n_14203)
);

NAND2xp5_ASAP7_75t_L g14204 ( 
.A(n_14101),
.B(n_2846),
.Y(n_14204)
);

OAI211xp5_ASAP7_75t_L g14205 ( 
.A1(n_14118),
.A2(n_3442),
.B(n_3443),
.C(n_3441),
.Y(n_14205)
);

AOI211xp5_ASAP7_75t_L g14206 ( 
.A1(n_14118),
.A2(n_2850),
.B(n_2847),
.C(n_2849),
.Y(n_14206)
);

NAND3xp33_ASAP7_75t_SL g14207 ( 
.A(n_14066),
.B(n_2851),
.C(n_2852),
.Y(n_14207)
);

OAI211xp5_ASAP7_75t_L g14208 ( 
.A1(n_14118),
.A2(n_3446),
.B(n_3448),
.C(n_3445),
.Y(n_14208)
);

AND2x2_ASAP7_75t_L g14209 ( 
.A(n_14122),
.B(n_2851),
.Y(n_14209)
);

INVx1_ASAP7_75t_L g14210 ( 
.A(n_14081),
.Y(n_14210)
);

NAND2xp5_ASAP7_75t_L g14211 ( 
.A(n_14101),
.B(n_2852),
.Y(n_14211)
);

NOR3xp33_ASAP7_75t_L g14212 ( 
.A(n_14137),
.B(n_2853),
.C(n_2854),
.Y(n_14212)
);

AOI221xp5_ASAP7_75t_L g14213 ( 
.A1(n_14147),
.A2(n_2855),
.B1(n_2853),
.B2(n_2854),
.C(n_2856),
.Y(n_14213)
);

NOR2x1_ASAP7_75t_L g14214 ( 
.A(n_14149),
.B(n_2856),
.Y(n_14214)
);

NAND4xp75_ASAP7_75t_L g14215 ( 
.A(n_14196),
.B(n_2859),
.C(n_2857),
.D(n_2858),
.Y(n_14215)
);

INVx1_ASAP7_75t_L g14216 ( 
.A(n_14175),
.Y(n_14216)
);

NAND3xp33_ASAP7_75t_L g14217 ( 
.A(n_14160),
.B(n_2857),
.C(n_2858),
.Y(n_14217)
);

NOR3xp33_ASAP7_75t_L g14218 ( 
.A(n_14198),
.B(n_2859),
.C(n_2860),
.Y(n_14218)
);

NOR2xp33_ASAP7_75t_SL g14219 ( 
.A(n_14165),
.B(n_2860),
.Y(n_14219)
);

NOR2xp33_ASAP7_75t_L g14220 ( 
.A(n_14168),
.B(n_2861),
.Y(n_14220)
);

AND4x1_ASAP7_75t_L g14221 ( 
.A(n_14148),
.B(n_2864),
.C(n_2862),
.D(n_2863),
.Y(n_14221)
);

NAND4xp75_ASAP7_75t_L g14222 ( 
.A(n_14138),
.B(n_2864),
.C(n_2862),
.D(n_2863),
.Y(n_14222)
);

O2A1O1Ixp33_ASAP7_75t_L g14223 ( 
.A1(n_14145),
.A2(n_2867),
.B(n_2868),
.C(n_2866),
.Y(n_14223)
);

NAND2xp5_ASAP7_75t_L g14224 ( 
.A(n_14201),
.B(n_2865),
.Y(n_14224)
);

NAND5xp2_ASAP7_75t_L g14225 ( 
.A(n_14155),
.B(n_14139),
.C(n_14135),
.D(n_14190),
.E(n_14170),
.Y(n_14225)
);

OAI211xp5_ASAP7_75t_L g14226 ( 
.A1(n_14202),
.A2(n_3455),
.B(n_3442),
.C(n_2867),
.Y(n_14226)
);

NAND3xp33_ASAP7_75t_L g14227 ( 
.A(n_14176),
.B(n_2865),
.C(n_2866),
.Y(n_14227)
);

OAI221xp5_ASAP7_75t_L g14228 ( 
.A1(n_14143),
.A2(n_2870),
.B1(n_2868),
.B2(n_2869),
.C(n_2871),
.Y(n_14228)
);

NAND2xp5_ASAP7_75t_L g14229 ( 
.A(n_14140),
.B(n_14206),
.Y(n_14229)
);

AOI222xp33_ASAP7_75t_L g14230 ( 
.A1(n_14157),
.A2(n_2872),
.B1(n_2874),
.B2(n_2869),
.C1(n_2870),
.C2(n_2873),
.Y(n_14230)
);

OAI211xp5_ASAP7_75t_SL g14231 ( 
.A1(n_14203),
.A2(n_2874),
.B(n_2872),
.C(n_2873),
.Y(n_14231)
);

NOR3x1_ASAP7_75t_L g14232 ( 
.A(n_14207),
.B(n_2875),
.C(n_2876),
.Y(n_14232)
);

AOI211xp5_ASAP7_75t_L g14233 ( 
.A1(n_14205),
.A2(n_2878),
.B(n_2875),
.C(n_2877),
.Y(n_14233)
);

AOI21xp33_ASAP7_75t_SL g14234 ( 
.A1(n_14169),
.A2(n_2879),
.B(n_2878),
.Y(n_14234)
);

NOR2x1_ASAP7_75t_L g14235 ( 
.A(n_14200),
.B(n_2877),
.Y(n_14235)
);

NOR3xp33_ASAP7_75t_L g14236 ( 
.A(n_14187),
.B(n_2879),
.C(n_2880),
.Y(n_14236)
);

NAND3xp33_ASAP7_75t_L g14237 ( 
.A(n_14152),
.B(n_2880),
.C(n_2881),
.Y(n_14237)
);

NOR2x1_ASAP7_75t_L g14238 ( 
.A(n_14204),
.B(n_2882),
.Y(n_14238)
);

NAND2xp5_ASAP7_75t_L g14239 ( 
.A(n_14150),
.B(n_2882),
.Y(n_14239)
);

AOI211x1_ASAP7_75t_L g14240 ( 
.A1(n_14208),
.A2(n_2885),
.B(n_2883),
.C(n_2884),
.Y(n_14240)
);

NOR2x1_ASAP7_75t_L g14241 ( 
.A(n_14211),
.B(n_2884),
.Y(n_14241)
);

NOR4xp25_ASAP7_75t_L g14242 ( 
.A(n_14144),
.B(n_2888),
.C(n_2885),
.D(n_2886),
.Y(n_14242)
);

NAND4xp75_ASAP7_75t_L g14243 ( 
.A(n_14159),
.B(n_2889),
.C(n_2886),
.D(n_2888),
.Y(n_14243)
);

AND2x2_ASAP7_75t_L g14244 ( 
.A(n_14141),
.B(n_2889),
.Y(n_14244)
);

NOR2xp33_ASAP7_75t_L g14245 ( 
.A(n_14189),
.B(n_2890),
.Y(n_14245)
);

OAI221xp5_ASAP7_75t_L g14246 ( 
.A1(n_14174),
.A2(n_2892),
.B1(n_2890),
.B2(n_2891),
.C(n_2893),
.Y(n_14246)
);

A2O1A1Ixp33_ASAP7_75t_L g14247 ( 
.A1(n_14194),
.A2(n_2895),
.B(n_2892),
.C(n_2894),
.Y(n_14247)
);

NOR2x1_ASAP7_75t_L g14248 ( 
.A(n_14172),
.B(n_2896),
.Y(n_14248)
);

O2A1O1Ixp33_ASAP7_75t_L g14249 ( 
.A1(n_14179),
.A2(n_2898),
.B(n_2899),
.C(n_2897),
.Y(n_14249)
);

NAND2xp5_ASAP7_75t_L g14250 ( 
.A(n_14186),
.B(n_2896),
.Y(n_14250)
);

NOR2x1_ASAP7_75t_L g14251 ( 
.A(n_14158),
.B(n_2898),
.Y(n_14251)
);

O2A1O1Ixp5_ASAP7_75t_L g14252 ( 
.A1(n_14171),
.A2(n_2902),
.B(n_2900),
.C(n_2901),
.Y(n_14252)
);

NAND3xp33_ASAP7_75t_SL g14253 ( 
.A(n_14181),
.B(n_2901),
.C(n_2902),
.Y(n_14253)
);

NAND2xp5_ASAP7_75t_L g14254 ( 
.A(n_14142),
.B(n_2903),
.Y(n_14254)
);

OAI221xp5_ASAP7_75t_L g14255 ( 
.A1(n_14192),
.A2(n_2905),
.B1(n_2903),
.B2(n_2904),
.C(n_2906),
.Y(n_14255)
);

NAND2xp5_ASAP7_75t_L g14256 ( 
.A(n_14183),
.B(n_2907),
.Y(n_14256)
);

NOR3xp33_ASAP7_75t_L g14257 ( 
.A(n_14146),
.B(n_2907),
.C(n_2908),
.Y(n_14257)
);

NAND2xp5_ASAP7_75t_L g14258 ( 
.A(n_14180),
.B(n_14197),
.Y(n_14258)
);

NOR2xp33_ASAP7_75t_L g14259 ( 
.A(n_14156),
.B(n_2908),
.Y(n_14259)
);

AND4x1_ASAP7_75t_L g14260 ( 
.A(n_14178),
.B(n_2911),
.C(n_2909),
.D(n_2910),
.Y(n_14260)
);

OAI211xp5_ASAP7_75t_L g14261 ( 
.A1(n_14154),
.A2(n_3452),
.B(n_3435),
.C(n_2911),
.Y(n_14261)
);

NAND3xp33_ASAP7_75t_L g14262 ( 
.A(n_14195),
.B(n_2909),
.C(n_2910),
.Y(n_14262)
);

AOI221xp5_ASAP7_75t_L g14263 ( 
.A1(n_14193),
.A2(n_2914),
.B1(n_2912),
.B2(n_2913),
.C(n_2915),
.Y(n_14263)
);

NAND2xp5_ASAP7_75t_L g14264 ( 
.A(n_14209),
.B(n_2913),
.Y(n_14264)
);

NOR3xp33_ASAP7_75t_L g14265 ( 
.A(n_14199),
.B(n_2914),
.C(n_2915),
.Y(n_14265)
);

NAND2xp5_ASAP7_75t_SL g14266 ( 
.A(n_14173),
.B(n_2916),
.Y(n_14266)
);

AOI21xp5_ASAP7_75t_L g14267 ( 
.A1(n_14184),
.A2(n_2917),
.B(n_2919),
.Y(n_14267)
);

NOR3xp33_ASAP7_75t_L g14268 ( 
.A(n_14210),
.B(n_2919),
.C(n_2920),
.Y(n_14268)
);

NAND3xp33_ASAP7_75t_L g14269 ( 
.A(n_14177),
.B(n_14191),
.C(n_14167),
.Y(n_14269)
);

INVx1_ASAP7_75t_SL g14270 ( 
.A(n_14222),
.Y(n_14270)
);

XNOR2xp5_ASAP7_75t_L g14271 ( 
.A(n_14260),
.B(n_14136),
.Y(n_14271)
);

NOR2x1p5_ASAP7_75t_L g14272 ( 
.A(n_14243),
.B(n_14151),
.Y(n_14272)
);

INVx2_ASAP7_75t_SL g14273 ( 
.A(n_14248),
.Y(n_14273)
);

AND2x2_ASAP7_75t_L g14274 ( 
.A(n_14244),
.B(n_14153),
.Y(n_14274)
);

INVx1_ASAP7_75t_L g14275 ( 
.A(n_14214),
.Y(n_14275)
);

OR2x2_ASAP7_75t_L g14276 ( 
.A(n_14242),
.B(n_14163),
.Y(n_14276)
);

NAND2xp5_ASAP7_75t_L g14277 ( 
.A(n_14212),
.B(n_14162),
.Y(n_14277)
);

INVx1_ASAP7_75t_SL g14278 ( 
.A(n_14215),
.Y(n_14278)
);

INVx1_ASAP7_75t_L g14279 ( 
.A(n_14264),
.Y(n_14279)
);

AND2x2_ASAP7_75t_L g14280 ( 
.A(n_14245),
.B(n_14161),
.Y(n_14280)
);

NAND2xp5_ASAP7_75t_L g14281 ( 
.A(n_14236),
.B(n_14230),
.Y(n_14281)
);

INVx1_ASAP7_75t_L g14282 ( 
.A(n_14239),
.Y(n_14282)
);

XOR2x2_ASAP7_75t_L g14283 ( 
.A(n_14217),
.B(n_14251),
.Y(n_14283)
);

NAND2xp5_ASAP7_75t_L g14284 ( 
.A(n_14257),
.B(n_14164),
.Y(n_14284)
);

OR2x2_ASAP7_75t_L g14285 ( 
.A(n_14253),
.B(n_14182),
.Y(n_14285)
);

AND2x4_ASAP7_75t_L g14286 ( 
.A(n_14269),
.B(n_14185),
.Y(n_14286)
);

NOR2x1_ASAP7_75t_SL g14287 ( 
.A(n_14261),
.B(n_14188),
.Y(n_14287)
);

INVx1_ASAP7_75t_SL g14288 ( 
.A(n_14235),
.Y(n_14288)
);

INVx1_ASAP7_75t_L g14289 ( 
.A(n_14238),
.Y(n_14289)
);

AND2x4_ASAP7_75t_L g14290 ( 
.A(n_14241),
.B(n_14166),
.Y(n_14290)
);

OR2x2_ASAP7_75t_L g14291 ( 
.A(n_14254),
.B(n_2920),
.Y(n_14291)
);

INVx1_ASAP7_75t_L g14292 ( 
.A(n_14240),
.Y(n_14292)
);

NOR2x1p5_ASAP7_75t_L g14293 ( 
.A(n_14224),
.B(n_2923),
.Y(n_14293)
);

AND2x4_ASAP7_75t_L g14294 ( 
.A(n_14216),
.B(n_2923),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_14256),
.Y(n_14295)
);

NAND2xp5_ASAP7_75t_L g14296 ( 
.A(n_14265),
.B(n_2924),
.Y(n_14296)
);

INVx1_ASAP7_75t_L g14297 ( 
.A(n_14221),
.Y(n_14297)
);

NAND2xp5_ASAP7_75t_L g14298 ( 
.A(n_14268),
.B(n_2924),
.Y(n_14298)
);

OR2x2_ASAP7_75t_L g14299 ( 
.A(n_14250),
.B(n_14227),
.Y(n_14299)
);

NAND2xp5_ASAP7_75t_L g14300 ( 
.A(n_14218),
.B(n_3429),
.Y(n_14300)
);

INVx1_ASAP7_75t_L g14301 ( 
.A(n_14219),
.Y(n_14301)
);

AND2x2_ASAP7_75t_L g14302 ( 
.A(n_14220),
.B(n_2925),
.Y(n_14302)
);

OR2x2_ASAP7_75t_L g14303 ( 
.A(n_14247),
.B(n_14262),
.Y(n_14303)
);

OAI21xp5_ASAP7_75t_SL g14304 ( 
.A1(n_14231),
.A2(n_2928),
.B(n_2927),
.Y(n_14304)
);

INVx3_ASAP7_75t_L g14305 ( 
.A(n_14258),
.Y(n_14305)
);

NOR2xp33_ASAP7_75t_L g14306 ( 
.A(n_14234),
.B(n_2926),
.Y(n_14306)
);

INVx1_ASAP7_75t_L g14307 ( 
.A(n_14252),
.Y(n_14307)
);

INVx1_ASAP7_75t_L g14308 ( 
.A(n_14223),
.Y(n_14308)
);

NAND2xp5_ASAP7_75t_L g14309 ( 
.A(n_14213),
.B(n_14267),
.Y(n_14309)
);

HB1xp67_ASAP7_75t_L g14310 ( 
.A(n_14232),
.Y(n_14310)
);

NOR3xp33_ASAP7_75t_L g14311 ( 
.A(n_14225),
.B(n_2926),
.C(n_2927),
.Y(n_14311)
);

OR2x2_ASAP7_75t_L g14312 ( 
.A(n_14237),
.B(n_2929),
.Y(n_14312)
);

INVx1_ASAP7_75t_L g14313 ( 
.A(n_14226),
.Y(n_14313)
);

INVx1_ASAP7_75t_L g14314 ( 
.A(n_14249),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_14266),
.Y(n_14315)
);

INVx1_ASAP7_75t_L g14316 ( 
.A(n_14259),
.Y(n_14316)
);

INVx1_ASAP7_75t_L g14317 ( 
.A(n_14233),
.Y(n_14317)
);

INVx1_ASAP7_75t_L g14318 ( 
.A(n_14229),
.Y(n_14318)
);

INVx1_ASAP7_75t_L g14319 ( 
.A(n_14246),
.Y(n_14319)
);

XOR2x2_ASAP7_75t_L g14320 ( 
.A(n_14263),
.B(n_2929),
.Y(n_14320)
);

INVxp67_ASAP7_75t_L g14321 ( 
.A(n_14228),
.Y(n_14321)
);

INVx1_ASAP7_75t_L g14322 ( 
.A(n_14255),
.Y(n_14322)
);

NAND2x1_ASAP7_75t_L g14323 ( 
.A(n_14248),
.B(n_2930),
.Y(n_14323)
);

INVx2_ASAP7_75t_L g14324 ( 
.A(n_14222),
.Y(n_14324)
);

NAND2xp5_ASAP7_75t_L g14325 ( 
.A(n_14212),
.B(n_3438),
.Y(n_14325)
);

NAND3xp33_ASAP7_75t_L g14326 ( 
.A(n_14212),
.B(n_2930),
.C(n_2931),
.Y(n_14326)
);

NAND2xp5_ASAP7_75t_L g14327 ( 
.A(n_14212),
.B(n_3439),
.Y(n_14327)
);

XOR2xp5_ASAP7_75t_L g14328 ( 
.A(n_14243),
.B(n_2931),
.Y(n_14328)
);

NOR2xp33_ASAP7_75t_L g14329 ( 
.A(n_14231),
.B(n_2932),
.Y(n_14329)
);

INVx2_ASAP7_75t_SL g14330 ( 
.A(n_14248),
.Y(n_14330)
);

NAND4xp25_ASAP7_75t_L g14331 ( 
.A(n_14311),
.B(n_2935),
.C(n_2933),
.D(n_2934),
.Y(n_14331)
);

INVx2_ASAP7_75t_L g14332 ( 
.A(n_14294),
.Y(n_14332)
);

NOR2xp67_ASAP7_75t_L g14333 ( 
.A(n_14326),
.B(n_2935),
.Y(n_14333)
);

NOR3xp33_ASAP7_75t_L g14334 ( 
.A(n_14273),
.B(n_2934),
.C(n_2936),
.Y(n_14334)
);

HB1xp67_ASAP7_75t_L g14335 ( 
.A(n_14323),
.Y(n_14335)
);

NAND4xp75_ASAP7_75t_L g14336 ( 
.A(n_14302),
.B(n_2938),
.C(n_2936),
.D(n_2937),
.Y(n_14336)
);

NAND4xp25_ASAP7_75t_L g14337 ( 
.A(n_14329),
.B(n_2940),
.C(n_2937),
.D(n_2938),
.Y(n_14337)
);

OA211x2_ASAP7_75t_L g14338 ( 
.A1(n_14306),
.A2(n_2943),
.B(n_2941),
.C(n_2942),
.Y(n_14338)
);

AND5x1_ASAP7_75t_L g14339 ( 
.A(n_14320),
.B(n_2945),
.C(n_2941),
.D(n_2943),
.E(n_2946),
.Y(n_14339)
);

INVxp67_ASAP7_75t_SL g14340 ( 
.A(n_14291),
.Y(n_14340)
);

NOR4xp25_ASAP7_75t_L g14341 ( 
.A(n_14270),
.B(n_3446),
.C(n_3434),
.D(n_2947),
.Y(n_14341)
);

NAND2x1p5_ASAP7_75t_L g14342 ( 
.A(n_14330),
.B(n_2945),
.Y(n_14342)
);

NAND3xp33_ASAP7_75t_L g14343 ( 
.A(n_14297),
.B(n_14271),
.C(n_14292),
.Y(n_14343)
);

AND2x2_ASAP7_75t_L g14344 ( 
.A(n_14293),
.B(n_2946),
.Y(n_14344)
);

NOR2xp67_ASAP7_75t_L g14345 ( 
.A(n_14276),
.B(n_2948),
.Y(n_14345)
);

NOR2xp33_ASAP7_75t_L g14346 ( 
.A(n_14304),
.B(n_14325),
.Y(n_14346)
);

NAND4xp25_ASAP7_75t_SL g14347 ( 
.A(n_14327),
.B(n_2950),
.C(n_2947),
.D(n_2949),
.Y(n_14347)
);

NOR3xp33_ASAP7_75t_SL g14348 ( 
.A(n_14277),
.B(n_2949),
.C(n_2951),
.Y(n_14348)
);

OR2x2_ASAP7_75t_L g14349 ( 
.A(n_14300),
.B(n_2952),
.Y(n_14349)
);

AOI211xp5_ASAP7_75t_L g14350 ( 
.A1(n_14296),
.A2(n_2955),
.B(n_2953),
.C(n_2954),
.Y(n_14350)
);

NOR2x1_ASAP7_75t_L g14351 ( 
.A(n_14275),
.B(n_2955),
.Y(n_14351)
);

NOR2x1_ASAP7_75t_SL g14352 ( 
.A(n_14312),
.B(n_2956),
.Y(n_14352)
);

INVx1_ASAP7_75t_L g14353 ( 
.A(n_14328),
.Y(n_14353)
);

NAND4xp75_ASAP7_75t_L g14354 ( 
.A(n_14313),
.B(n_2958),
.C(n_2953),
.D(n_2957),
.Y(n_14354)
);

NOR4xp75_ASAP7_75t_L g14355 ( 
.A(n_14284),
.B(n_2959),
.C(n_2957),
.D(n_2958),
.Y(n_14355)
);

NOR2x1p5_ASAP7_75t_L g14356 ( 
.A(n_14298),
.B(n_2959),
.Y(n_14356)
);

INVx1_ASAP7_75t_L g14357 ( 
.A(n_14310),
.Y(n_14357)
);

NOR3xp33_ASAP7_75t_L g14358 ( 
.A(n_14305),
.B(n_2960),
.C(n_2961),
.Y(n_14358)
);

NOR2xp33_ASAP7_75t_L g14359 ( 
.A(n_14278),
.B(n_3431),
.Y(n_14359)
);

INVx2_ASAP7_75t_SL g14360 ( 
.A(n_14272),
.Y(n_14360)
);

AND2x4_ASAP7_75t_L g14361 ( 
.A(n_14289),
.B(n_2960),
.Y(n_14361)
);

AOI22xp5_ASAP7_75t_L g14362 ( 
.A1(n_14286),
.A2(n_2963),
.B1(n_2961),
.B2(n_2962),
.Y(n_14362)
);

INVx1_ASAP7_75t_L g14363 ( 
.A(n_14283),
.Y(n_14363)
);

AND2x4_ASAP7_75t_L g14364 ( 
.A(n_14324),
.B(n_2962),
.Y(n_14364)
);

NOR2x1_ASAP7_75t_L g14365 ( 
.A(n_14290),
.B(n_2964),
.Y(n_14365)
);

NAND2xp5_ASAP7_75t_L g14366 ( 
.A(n_14288),
.B(n_2965),
.Y(n_14366)
);

NAND2xp5_ASAP7_75t_L g14367 ( 
.A(n_14307),
.B(n_2966),
.Y(n_14367)
);

NOR3xp33_ASAP7_75t_L g14368 ( 
.A(n_14301),
.B(n_2963),
.C(n_2967),
.Y(n_14368)
);

NAND4xp25_ASAP7_75t_L g14369 ( 
.A(n_14281),
.B(n_2969),
.C(n_2967),
.D(n_2968),
.Y(n_14369)
);

AND2x4_ASAP7_75t_L g14370 ( 
.A(n_14274),
.B(n_2968),
.Y(n_14370)
);

NOR3xp33_ASAP7_75t_L g14371 ( 
.A(n_14318),
.B(n_2969),
.C(n_2970),
.Y(n_14371)
);

NOR2xp33_ASAP7_75t_L g14372 ( 
.A(n_14308),
.B(n_3453),
.Y(n_14372)
);

INVx2_ASAP7_75t_SL g14373 ( 
.A(n_14285),
.Y(n_14373)
);

NAND3xp33_ASAP7_75t_SL g14374 ( 
.A(n_14314),
.B(n_14317),
.C(n_14299),
.Y(n_14374)
);

NOR4xp75_ASAP7_75t_L g14375 ( 
.A(n_14309),
.B(n_2972),
.C(n_2970),
.D(n_2971),
.Y(n_14375)
);

OAI21xp33_ASAP7_75t_L g14376 ( 
.A1(n_14279),
.A2(n_2972),
.B(n_2973),
.Y(n_14376)
);

AND2x2_ASAP7_75t_L g14377 ( 
.A(n_14287),
.B(n_2973),
.Y(n_14377)
);

NAND3xp33_ASAP7_75t_L g14378 ( 
.A(n_14321),
.B(n_2974),
.C(n_2975),
.Y(n_14378)
);

INVx1_ASAP7_75t_L g14379 ( 
.A(n_14303),
.Y(n_14379)
);

NAND3xp33_ASAP7_75t_L g14380 ( 
.A(n_14319),
.B(n_2974),
.C(n_2976),
.Y(n_14380)
);

NOR4xp75_ASAP7_75t_L g14381 ( 
.A(n_14280),
.B(n_2978),
.C(n_2976),
.D(n_2977),
.Y(n_14381)
);

NOR3xp33_ASAP7_75t_L g14382 ( 
.A(n_14315),
.B(n_2978),
.C(n_2980),
.Y(n_14382)
);

AND2x2_ASAP7_75t_L g14383 ( 
.A(n_14322),
.B(n_14316),
.Y(n_14383)
);

NOR2x1_ASAP7_75t_L g14384 ( 
.A(n_14282),
.B(n_2981),
.Y(n_14384)
);

NOR3xp33_ASAP7_75t_SL g14385 ( 
.A(n_14295),
.B(n_2980),
.C(n_2981),
.Y(n_14385)
);

NAND3xp33_ASAP7_75t_SL g14386 ( 
.A(n_14311),
.B(n_2982),
.C(n_2983),
.Y(n_14386)
);

INVx1_ASAP7_75t_L g14387 ( 
.A(n_14323),
.Y(n_14387)
);

NOR3xp33_ASAP7_75t_L g14388 ( 
.A(n_14311),
.B(n_2982),
.C(n_2983),
.Y(n_14388)
);

NAND2xp5_ASAP7_75t_L g14389 ( 
.A(n_14311),
.B(n_2985),
.Y(n_14389)
);

NOR3x1_ASAP7_75t_L g14390 ( 
.A(n_14323),
.B(n_2984),
.C(n_2986),
.Y(n_14390)
);

NAND3xp33_ASAP7_75t_SL g14391 ( 
.A(n_14311),
.B(n_2984),
.C(n_2988),
.Y(n_14391)
);

AOI211x1_ASAP7_75t_L g14392 ( 
.A1(n_14297),
.A2(n_2990),
.B(n_2988),
.C(n_2989),
.Y(n_14392)
);

AOI211xp5_ASAP7_75t_L g14393 ( 
.A1(n_14326),
.A2(n_2991),
.B(n_2989),
.C(n_2990),
.Y(n_14393)
);

NAND2xp5_ASAP7_75t_L g14394 ( 
.A(n_14311),
.B(n_2992),
.Y(n_14394)
);

NAND2xp5_ASAP7_75t_SL g14395 ( 
.A(n_14311),
.B(n_2991),
.Y(n_14395)
);

NOR2x1_ASAP7_75t_L g14396 ( 
.A(n_14323),
.B(n_2993),
.Y(n_14396)
);

NOR2x1_ASAP7_75t_L g14397 ( 
.A(n_14323),
.B(n_2993),
.Y(n_14397)
);

AOI22xp5_ASAP7_75t_L g14398 ( 
.A1(n_14388),
.A2(n_2995),
.B1(n_2992),
.B2(n_2994),
.Y(n_14398)
);

INVx1_ASAP7_75t_L g14399 ( 
.A(n_14377),
.Y(n_14399)
);

INVx1_ASAP7_75t_L g14400 ( 
.A(n_14365),
.Y(n_14400)
);

INVx1_ASAP7_75t_L g14401 ( 
.A(n_14351),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_14384),
.Y(n_14402)
);

INVx1_ASAP7_75t_SL g14403 ( 
.A(n_14366),
.Y(n_14403)
);

AND2x4_ASAP7_75t_L g14404 ( 
.A(n_14396),
.B(n_14397),
.Y(n_14404)
);

OAI21xp5_ASAP7_75t_L g14405 ( 
.A1(n_14343),
.A2(n_2994),
.B(n_2995),
.Y(n_14405)
);

BUFx3_ASAP7_75t_L g14406 ( 
.A(n_14367),
.Y(n_14406)
);

INVx2_ASAP7_75t_L g14407 ( 
.A(n_14342),
.Y(n_14407)
);

OAI22xp33_ASAP7_75t_L g14408 ( 
.A1(n_14331),
.A2(n_2998),
.B1(n_2996),
.B2(n_2997),
.Y(n_14408)
);

NOR2xp33_ASAP7_75t_SL g14409 ( 
.A(n_14359),
.B(n_2998),
.Y(n_14409)
);

NOR2x1_ASAP7_75t_L g14410 ( 
.A(n_14336),
.B(n_3440),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_14344),
.Y(n_14411)
);

AOI22xp33_ASAP7_75t_L g14412 ( 
.A1(n_14386),
.A2(n_3001),
.B1(n_2999),
.B2(n_3000),
.Y(n_14412)
);

NOR2x1_ASAP7_75t_L g14413 ( 
.A(n_14354),
.B(n_3443),
.Y(n_14413)
);

NOR2x2_ASAP7_75t_L g14414 ( 
.A(n_14332),
.B(n_3000),
.Y(n_14414)
);

AOI22xp5_ASAP7_75t_L g14415 ( 
.A1(n_14373),
.A2(n_14360),
.B1(n_14357),
.B2(n_14391),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_14345),
.Y(n_14416)
);

AOI22xp5_ASAP7_75t_L g14417 ( 
.A1(n_14363),
.A2(n_3003),
.B1(n_3001),
.B2(n_3002),
.Y(n_14417)
);

AOI31xp33_ASAP7_75t_L g14418 ( 
.A1(n_14335),
.A2(n_3004),
.A3(n_3002),
.B(n_3003),
.Y(n_14418)
);

INVx1_ASAP7_75t_L g14419 ( 
.A(n_14338),
.Y(n_14419)
);

NAND2xp5_ASAP7_75t_SL g14420 ( 
.A(n_14341),
.B(n_3004),
.Y(n_14420)
);

NOR2x1_ASAP7_75t_L g14421 ( 
.A(n_14387),
.B(n_3005),
.Y(n_14421)
);

CKINVDCx20_ASAP7_75t_R g14422 ( 
.A(n_14353),
.Y(n_14422)
);

INVx1_ASAP7_75t_L g14423 ( 
.A(n_14375),
.Y(n_14423)
);

INVx1_ASAP7_75t_L g14424 ( 
.A(n_14349),
.Y(n_14424)
);

INVx1_ASAP7_75t_L g14425 ( 
.A(n_14355),
.Y(n_14425)
);

NAND2xp5_ASAP7_75t_L g14426 ( 
.A(n_14372),
.B(n_14350),
.Y(n_14426)
);

NAND2xp5_ASAP7_75t_L g14427 ( 
.A(n_14385),
.B(n_3005),
.Y(n_14427)
);

NAND3xp33_ASAP7_75t_SL g14428 ( 
.A(n_14393),
.B(n_3006),
.C(n_3007),
.Y(n_14428)
);

NAND3x1_ASAP7_75t_L g14429 ( 
.A(n_14381),
.B(n_3006),
.C(n_3008),
.Y(n_14429)
);

AOI22xp5_ASAP7_75t_L g14430 ( 
.A1(n_14379),
.A2(n_3010),
.B1(n_3008),
.B2(n_3009),
.Y(n_14430)
);

AOI22xp5_ASAP7_75t_L g14431 ( 
.A1(n_14337),
.A2(n_3011),
.B1(n_3009),
.B2(n_3010),
.Y(n_14431)
);

HB1xp67_ASAP7_75t_L g14432 ( 
.A(n_14390),
.Y(n_14432)
);

INVx1_ASAP7_75t_L g14433 ( 
.A(n_14389),
.Y(n_14433)
);

INVx2_ASAP7_75t_L g14434 ( 
.A(n_14370),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_14394),
.Y(n_14435)
);

INVx1_ASAP7_75t_L g14436 ( 
.A(n_14352),
.Y(n_14436)
);

INVx1_ASAP7_75t_L g14437 ( 
.A(n_14348),
.Y(n_14437)
);

INVxp67_ASAP7_75t_SL g14438 ( 
.A(n_14356),
.Y(n_14438)
);

INVx1_ASAP7_75t_L g14439 ( 
.A(n_14392),
.Y(n_14439)
);

NOR2x1_ASAP7_75t_L g14440 ( 
.A(n_14347),
.B(n_14380),
.Y(n_14440)
);

AOI22xp5_ASAP7_75t_L g14441 ( 
.A1(n_14374),
.A2(n_3014),
.B1(n_3011),
.B2(n_3012),
.Y(n_14441)
);

OAI22xp5_ASAP7_75t_L g14442 ( 
.A1(n_14378),
.A2(n_3016),
.B1(n_3014),
.B2(n_3015),
.Y(n_14442)
);

INVx1_ASAP7_75t_L g14443 ( 
.A(n_14395),
.Y(n_14443)
);

NAND2xp5_ASAP7_75t_SL g14444 ( 
.A(n_14333),
.B(n_14334),
.Y(n_14444)
);

NOR2xp67_ASAP7_75t_L g14445 ( 
.A(n_14369),
.B(n_3439),
.Y(n_14445)
);

INVx1_ASAP7_75t_L g14446 ( 
.A(n_14376),
.Y(n_14446)
);

INVx1_ASAP7_75t_L g14447 ( 
.A(n_14340),
.Y(n_14447)
);

INVx1_ASAP7_75t_L g14448 ( 
.A(n_14421),
.Y(n_14448)
);

NOR3xp33_ASAP7_75t_L g14449 ( 
.A(n_14447),
.B(n_14383),
.C(n_14346),
.Y(n_14449)
);

NOR3xp33_ASAP7_75t_L g14450 ( 
.A(n_14399),
.B(n_14368),
.C(n_14371),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_14427),
.Y(n_14451)
);

NOR2x1_ASAP7_75t_L g14452 ( 
.A(n_14404),
.B(n_14370),
.Y(n_14452)
);

AND2x4_ASAP7_75t_L g14453 ( 
.A(n_14404),
.B(n_14339),
.Y(n_14453)
);

NOR4xp25_ASAP7_75t_L g14454 ( 
.A(n_14400),
.B(n_14358),
.C(n_14382),
.D(n_14362),
.Y(n_14454)
);

NOR3xp33_ASAP7_75t_L g14455 ( 
.A(n_14416),
.B(n_14364),
.C(n_14361),
.Y(n_14455)
);

XNOR2xp5_ASAP7_75t_L g14456 ( 
.A(n_14429),
.B(n_14364),
.Y(n_14456)
);

NOR3x2_ASAP7_75t_L g14457 ( 
.A(n_14414),
.B(n_14361),
.C(n_3023),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_14410),
.Y(n_14458)
);

AND4x1_ASAP7_75t_L g14459 ( 
.A(n_14415),
.B(n_3017),
.C(n_3018),
.D(n_3016),
.Y(n_14459)
);

NAND4xp25_ASAP7_75t_SL g14460 ( 
.A(n_14412),
.B(n_14431),
.C(n_14398),
.D(n_14413),
.Y(n_14460)
);

AOI22xp5_ASAP7_75t_L g14461 ( 
.A1(n_14422),
.A2(n_14409),
.B1(n_14445),
.B2(n_14425),
.Y(n_14461)
);

NOR2x1p5_ASAP7_75t_L g14462 ( 
.A(n_14419),
.B(n_3015),
.Y(n_14462)
);

NAND2xp5_ASAP7_75t_L g14463 ( 
.A(n_14408),
.B(n_3019),
.Y(n_14463)
);

OAI221xp5_ASAP7_75t_L g14464 ( 
.A1(n_14405),
.A2(n_3022),
.B1(n_3020),
.B2(n_3021),
.C(n_3024),
.Y(n_14464)
);

NOR3xp33_ASAP7_75t_L g14465 ( 
.A(n_14436),
.B(n_14434),
.C(n_14401),
.Y(n_14465)
);

HB1xp67_ASAP7_75t_L g14466 ( 
.A(n_14442),
.Y(n_14466)
);

AND3x4_ASAP7_75t_L g14467 ( 
.A(n_14440),
.B(n_3030),
.C(n_3020),
.Y(n_14467)
);

AOI22xp5_ASAP7_75t_L g14468 ( 
.A1(n_14423),
.A2(n_3025),
.B1(n_3021),
.B2(n_3024),
.Y(n_14468)
);

AOI221xp5_ASAP7_75t_L g14469 ( 
.A1(n_14428),
.A2(n_3027),
.B1(n_3025),
.B2(n_3026),
.C(n_3028),
.Y(n_14469)
);

NAND2xp5_ASAP7_75t_L g14470 ( 
.A(n_14441),
.B(n_3026),
.Y(n_14470)
);

AOI21xp33_ASAP7_75t_L g14471 ( 
.A1(n_14402),
.A2(n_3435),
.B(n_3434),
.Y(n_14471)
);

NAND2x1p5_ASAP7_75t_L g14472 ( 
.A(n_14407),
.B(n_3027),
.Y(n_14472)
);

NOR2x1_ASAP7_75t_L g14473 ( 
.A(n_14420),
.B(n_3029),
.Y(n_14473)
);

NAND4xp25_ASAP7_75t_L g14474 ( 
.A(n_14437),
.B(n_3032),
.C(n_3029),
.D(n_3030),
.Y(n_14474)
);

NAND4xp25_ASAP7_75t_L g14475 ( 
.A(n_14403),
.B(n_14439),
.C(n_14426),
.D(n_14446),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_14432),
.Y(n_14476)
);

NAND2xp5_ASAP7_75t_L g14477 ( 
.A(n_14417),
.B(n_3033),
.Y(n_14477)
);

AND2x2_ASAP7_75t_L g14478 ( 
.A(n_14438),
.B(n_3033),
.Y(n_14478)
);

OAI221xp5_ASAP7_75t_L g14479 ( 
.A1(n_14443),
.A2(n_3036),
.B1(n_3034),
.B2(n_3035),
.C(n_3037),
.Y(n_14479)
);

NAND2xp5_ASAP7_75t_L g14480 ( 
.A(n_14411),
.B(n_3034),
.Y(n_14480)
);

NAND4xp75_ASAP7_75t_L g14481 ( 
.A(n_14444),
.B(n_3039),
.C(n_3035),
.D(n_3038),
.Y(n_14481)
);

NAND3xp33_ASAP7_75t_SL g14482 ( 
.A(n_14424),
.B(n_3039),
.C(n_3040),
.Y(n_14482)
);

OAI322xp33_ASAP7_75t_L g14483 ( 
.A1(n_14433),
.A2(n_3429),
.A3(n_3427),
.B1(n_3431),
.B2(n_3437),
.C1(n_3428),
.C2(n_3426),
.Y(n_14483)
);

NAND4xp75_ASAP7_75t_L g14484 ( 
.A(n_14435),
.B(n_3042),
.C(n_3040),
.D(n_3041),
.Y(n_14484)
);

HB1xp67_ASAP7_75t_L g14485 ( 
.A(n_14406),
.Y(n_14485)
);

NOR3xp33_ASAP7_75t_L g14486 ( 
.A(n_14475),
.B(n_14418),
.C(n_14430),
.Y(n_14486)
);

INVx1_ASAP7_75t_L g14487 ( 
.A(n_14457),
.Y(n_14487)
);

OR3x2_ASAP7_75t_L g14488 ( 
.A(n_14476),
.B(n_3041),
.C(n_3042),
.Y(n_14488)
);

OR2x2_ASAP7_75t_L g14489 ( 
.A(n_14482),
.B(n_3043),
.Y(n_14489)
);

AOI221x1_ASAP7_75t_L g14490 ( 
.A1(n_14465),
.A2(n_3045),
.B1(n_3043),
.B2(n_3044),
.C(n_3046),
.Y(n_14490)
);

NAND2xp5_ASAP7_75t_L g14491 ( 
.A(n_14462),
.B(n_3044),
.Y(n_14491)
);

NAND4xp75_ASAP7_75t_L g14492 ( 
.A(n_14452),
.B(n_14473),
.C(n_14461),
.D(n_14458),
.Y(n_14492)
);

OR2x2_ASAP7_75t_L g14493 ( 
.A(n_14463),
.B(n_3045),
.Y(n_14493)
);

NOR3xp33_ASAP7_75t_L g14494 ( 
.A(n_14449),
.B(n_3047),
.C(n_3048),
.Y(n_14494)
);

AOI21xp5_ASAP7_75t_L g14495 ( 
.A1(n_14448),
.A2(n_14453),
.B(n_14456),
.Y(n_14495)
);

OR2x2_ASAP7_75t_L g14496 ( 
.A(n_14470),
.B(n_14477),
.Y(n_14496)
);

OAI21xp33_ASAP7_75t_SL g14497 ( 
.A1(n_14469),
.A2(n_3048),
.B(n_3049),
.Y(n_14497)
);

INVx1_ASAP7_75t_SL g14498 ( 
.A(n_14472),
.Y(n_14498)
);

NOR3xp33_ASAP7_75t_L g14499 ( 
.A(n_14455),
.B(n_14485),
.C(n_14451),
.Y(n_14499)
);

OAI322xp33_ASAP7_75t_L g14500 ( 
.A1(n_14466),
.A2(n_3073),
.A3(n_3057),
.B1(n_3081),
.B2(n_3092),
.C1(n_3065),
.C2(n_3049),
.Y(n_14500)
);

NOR3xp33_ASAP7_75t_L g14501 ( 
.A(n_14450),
.B(n_3050),
.C(n_3051),
.Y(n_14501)
);

AO22x2_ASAP7_75t_L g14502 ( 
.A1(n_14453),
.A2(n_3053),
.B1(n_3054),
.B2(n_3052),
.Y(n_14502)
);

OAI22xp5_ASAP7_75t_L g14503 ( 
.A1(n_14464),
.A2(n_3055),
.B1(n_3050),
.B2(n_3052),
.Y(n_14503)
);

AND2x4_ASAP7_75t_L g14504 ( 
.A(n_14459),
.B(n_3055),
.Y(n_14504)
);

HB1xp67_ASAP7_75t_L g14505 ( 
.A(n_14467),
.Y(n_14505)
);

NAND2xp5_ASAP7_75t_L g14506 ( 
.A(n_14454),
.B(n_3056),
.Y(n_14506)
);

AOI22xp5_ASAP7_75t_L g14507 ( 
.A1(n_14460),
.A2(n_14481),
.B1(n_14484),
.B2(n_14474),
.Y(n_14507)
);

OAI322xp33_ASAP7_75t_L g14508 ( 
.A1(n_14468),
.A2(n_3080),
.A3(n_3064),
.B1(n_3090),
.B2(n_3099),
.C1(n_3072),
.C2(n_3056),
.Y(n_14508)
);

NOR3xp33_ASAP7_75t_L g14509 ( 
.A(n_14471),
.B(n_3057),
.C(n_3058),
.Y(n_14509)
);

AND2x2_ASAP7_75t_L g14510 ( 
.A(n_14478),
.B(n_3059),
.Y(n_14510)
);

NOR3xp33_ASAP7_75t_L g14511 ( 
.A(n_14479),
.B(n_3059),
.C(n_3060),
.Y(n_14511)
);

AOI21xp33_ASAP7_75t_L g14512 ( 
.A1(n_14480),
.A2(n_3060),
.B(n_3061),
.Y(n_14512)
);

NOR3xp33_ASAP7_75t_L g14513 ( 
.A(n_14483),
.B(n_3061),
.C(n_3062),
.Y(n_14513)
);

A2O1A1Ixp33_ASAP7_75t_L g14514 ( 
.A1(n_14469),
.A2(n_3066),
.B(n_3063),
.C(n_3065),
.Y(n_14514)
);

NAND3xp33_ASAP7_75t_L g14515 ( 
.A(n_14465),
.B(n_3063),
.C(n_3066),
.Y(n_14515)
);

OR2x2_ASAP7_75t_L g14516 ( 
.A(n_14482),
.B(n_3067),
.Y(n_14516)
);

XNOR2xp5_ASAP7_75t_L g14517 ( 
.A(n_14457),
.B(n_3067),
.Y(n_14517)
);

NAND4xp75_ASAP7_75t_L g14518 ( 
.A(n_14452),
.B(n_3070),
.C(n_3068),
.D(n_3069),
.Y(n_14518)
);

NOR2xp33_ASAP7_75t_L g14519 ( 
.A(n_14463),
.B(n_3068),
.Y(n_14519)
);

AOI221xp5_ASAP7_75t_L g14520 ( 
.A1(n_14454),
.A2(n_3073),
.B1(n_3070),
.B2(n_3071),
.C(n_3074),
.Y(n_14520)
);

NOR2x1_ASAP7_75t_L g14521 ( 
.A(n_14452),
.B(n_3071),
.Y(n_14521)
);

AOI22xp5_ASAP7_75t_L g14522 ( 
.A1(n_14465),
.A2(n_3076),
.B1(n_3077),
.B2(n_3075),
.Y(n_14522)
);

OAI221xp5_ASAP7_75t_L g14523 ( 
.A1(n_14469),
.A2(n_3076),
.B1(n_3074),
.B2(n_3075),
.C(n_3077),
.Y(n_14523)
);

A2O1A1Ixp33_ASAP7_75t_L g14524 ( 
.A1(n_14469),
.A2(n_3080),
.B(n_3078),
.C(n_3079),
.Y(n_14524)
);

AND2x4_ASAP7_75t_L g14525 ( 
.A(n_14486),
.B(n_3079),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_14521),
.Y(n_14526)
);

OAI22xp5_ASAP7_75t_L g14527 ( 
.A1(n_14488),
.A2(n_3084),
.B1(n_3081),
.B2(n_3083),
.Y(n_14527)
);

AND3x2_ASAP7_75t_L g14528 ( 
.A(n_14505),
.B(n_3083),
.C(n_3085),
.Y(n_14528)
);

HB1xp67_ASAP7_75t_L g14529 ( 
.A(n_14510),
.Y(n_14529)
);

NOR2xp33_ASAP7_75t_L g14530 ( 
.A(n_14506),
.B(n_3086),
.Y(n_14530)
);

INVx1_ASAP7_75t_L g14531 ( 
.A(n_14517),
.Y(n_14531)
);

XOR2xp5_ASAP7_75t_L g14532 ( 
.A(n_14492),
.B(n_3088),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_14493),
.Y(n_14533)
);

AOI22x1_ASAP7_75t_L g14534 ( 
.A1(n_14495),
.A2(n_3092),
.B1(n_3089),
.B2(n_3090),
.Y(n_14534)
);

BUFx2_ASAP7_75t_L g14535 ( 
.A(n_14504),
.Y(n_14535)
);

XNOR2xp5_ASAP7_75t_L g14536 ( 
.A(n_14507),
.B(n_3089),
.Y(n_14536)
);

O2A1O1Ixp33_ASAP7_75t_L g14537 ( 
.A1(n_14499),
.A2(n_3095),
.B(n_3093),
.C(n_3094),
.Y(n_14537)
);

NAND2xp5_ASAP7_75t_L g14538 ( 
.A(n_14504),
.B(n_3094),
.Y(n_14538)
);

AND2x4_ASAP7_75t_L g14539 ( 
.A(n_14509),
.B(n_14498),
.Y(n_14539)
);

AOI22xp5_ASAP7_75t_L g14540 ( 
.A1(n_14519),
.A2(n_3103),
.B1(n_3111),
.B2(n_3093),
.Y(n_14540)
);

INVx1_ASAP7_75t_L g14541 ( 
.A(n_14491),
.Y(n_14541)
);

AND3x2_ASAP7_75t_L g14542 ( 
.A(n_14494),
.B(n_3096),
.C(n_3097),
.Y(n_14542)
);

AND3x1_ASAP7_75t_L g14543 ( 
.A(n_14511),
.B(n_3097),
.C(n_3098),
.Y(n_14543)
);

AND2x4_ASAP7_75t_L g14544 ( 
.A(n_14487),
.B(n_3098),
.Y(n_14544)
);

AOI21xp5_ASAP7_75t_SL g14545 ( 
.A1(n_14489),
.A2(n_3099),
.B(n_3100),
.Y(n_14545)
);

AO21x2_ASAP7_75t_L g14546 ( 
.A1(n_14513),
.A2(n_3100),
.B(n_3101),
.Y(n_14546)
);

NOR2xp67_ASAP7_75t_L g14547 ( 
.A(n_14516),
.B(n_3101),
.Y(n_14547)
);

XNOR2x1_ASAP7_75t_SL g14548 ( 
.A(n_14497),
.B(n_3102),
.Y(n_14548)
);

XNOR2xp5_ASAP7_75t_L g14549 ( 
.A(n_14515),
.B(n_3102),
.Y(n_14549)
);

INVx2_ASAP7_75t_L g14550 ( 
.A(n_14518),
.Y(n_14550)
);

OR3x2_ASAP7_75t_L g14551 ( 
.A(n_14496),
.B(n_3106),
.C(n_3105),
.Y(n_14551)
);

NAND2xp5_ASAP7_75t_L g14552 ( 
.A(n_14514),
.B(n_3105),
.Y(n_14552)
);

NOR2x1_ASAP7_75t_L g14553 ( 
.A(n_14508),
.B(n_3104),
.Y(n_14553)
);

INVx2_ASAP7_75t_L g14554 ( 
.A(n_14502),
.Y(n_14554)
);

NAND2x1p5_ASAP7_75t_L g14555 ( 
.A(n_14522),
.B(n_3104),
.Y(n_14555)
);

NAND3xp33_ASAP7_75t_L g14556 ( 
.A(n_14524),
.B(n_3106),
.C(n_3107),
.Y(n_14556)
);

AOI21xp33_ASAP7_75t_SL g14557 ( 
.A1(n_14503),
.A2(n_3107),
.B(n_3108),
.Y(n_14557)
);

OAI22xp5_ASAP7_75t_L g14558 ( 
.A1(n_14523),
.A2(n_3110),
.B1(n_3108),
.B2(n_3109),
.Y(n_14558)
);

NAND2xp5_ASAP7_75t_L g14559 ( 
.A(n_14501),
.B(n_14512),
.Y(n_14559)
);

INVx2_ASAP7_75t_L g14560 ( 
.A(n_14502),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_14490),
.Y(n_14561)
);

OR2x2_ASAP7_75t_L g14562 ( 
.A(n_14520),
.B(n_3109),
.Y(n_14562)
);

NAND3x1_ASAP7_75t_L g14563 ( 
.A(n_14500),
.B(n_3112),
.C(n_3111),
.Y(n_14563)
);

AOI221xp5_ASAP7_75t_L g14564 ( 
.A1(n_14557),
.A2(n_14558),
.B1(n_14543),
.B2(n_14545),
.C(n_14530),
.Y(n_14564)
);

AOI322xp5_ASAP7_75t_L g14565 ( 
.A1(n_14553),
.A2(n_3116),
.A3(n_3115),
.B1(n_3113),
.B2(n_3110),
.C1(n_3112),
.C2(n_3114),
.Y(n_14565)
);

INVx1_ASAP7_75t_L g14566 ( 
.A(n_14532),
.Y(n_14566)
);

AOI321xp33_ASAP7_75t_L g14567 ( 
.A1(n_14550),
.A2(n_3116),
.A3(n_3118),
.B1(n_3114),
.B2(n_3115),
.C(n_3117),
.Y(n_14567)
);

AOI22xp33_ASAP7_75t_SL g14568 ( 
.A1(n_14538),
.A2(n_3120),
.B1(n_3117),
.B2(n_3118),
.Y(n_14568)
);

NOR3xp33_ASAP7_75t_L g14569 ( 
.A(n_14526),
.B(n_3120),
.C(n_3121),
.Y(n_14569)
);

INVx1_ASAP7_75t_L g14570 ( 
.A(n_14536),
.Y(n_14570)
);

AOI322xp5_ASAP7_75t_L g14571 ( 
.A1(n_14561),
.A2(n_3127),
.A3(n_3125),
.B1(n_3123),
.B2(n_3121),
.C1(n_3122),
.C2(n_3124),
.Y(n_14571)
);

OAI211xp5_ASAP7_75t_L g14572 ( 
.A1(n_14547),
.A2(n_3125),
.B(n_3122),
.C(n_3123),
.Y(n_14572)
);

AOI22xp5_ASAP7_75t_L g14573 ( 
.A1(n_14527),
.A2(n_3130),
.B1(n_3127),
.B2(n_3129),
.Y(n_14573)
);

NAND2xp5_ASAP7_75t_L g14574 ( 
.A(n_14542),
.B(n_14525),
.Y(n_14574)
);

INVx1_ASAP7_75t_L g14575 ( 
.A(n_14549),
.Y(n_14575)
);

INVx2_ASAP7_75t_L g14576 ( 
.A(n_14528),
.Y(n_14576)
);

AOI221xp5_ASAP7_75t_L g14577 ( 
.A1(n_14556),
.A2(n_3131),
.B1(n_3129),
.B2(n_3130),
.C(n_3132),
.Y(n_14577)
);

OAI322xp33_ASAP7_75t_L g14578 ( 
.A1(n_14562),
.A2(n_3138),
.A3(n_3137),
.B1(n_3135),
.B2(n_3131),
.C1(n_3134),
.C2(n_3136),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_14551),
.Y(n_14579)
);

NOR2x1_ASAP7_75t_L g14580 ( 
.A(n_14554),
.B(n_3134),
.Y(n_14580)
);

AOI221xp5_ASAP7_75t_L g14581 ( 
.A1(n_14552),
.A2(n_3137),
.B1(n_3135),
.B2(n_3136),
.C(n_3139),
.Y(n_14581)
);

AOI322xp5_ASAP7_75t_L g14582 ( 
.A1(n_14529),
.A2(n_3144),
.A3(n_3143),
.B1(n_3141),
.B2(n_3139),
.C1(n_3140),
.C2(n_3142),
.Y(n_14582)
);

NAND2xp5_ASAP7_75t_L g14583 ( 
.A(n_14546),
.B(n_3142),
.Y(n_14583)
);

AOI322xp5_ASAP7_75t_L g14584 ( 
.A1(n_14531),
.A2(n_14539),
.A3(n_14535),
.B1(n_14560),
.B2(n_14541),
.C1(n_14533),
.C2(n_14559),
.Y(n_14584)
);

OAI221xp5_ASAP7_75t_L g14585 ( 
.A1(n_14534),
.A2(n_14555),
.B1(n_14537),
.B2(n_14540),
.C(n_14548),
.Y(n_14585)
);

INVx1_ASAP7_75t_L g14586 ( 
.A(n_14563),
.Y(n_14586)
);

INVx2_ASAP7_75t_SL g14587 ( 
.A(n_14544),
.Y(n_14587)
);

INVxp67_ASAP7_75t_SL g14588 ( 
.A(n_14547),
.Y(n_14588)
);

INVxp67_ASAP7_75t_SL g14589 ( 
.A(n_14547),
.Y(n_14589)
);

AOI322xp5_ASAP7_75t_L g14590 ( 
.A1(n_14530),
.A2(n_3149),
.A3(n_3148),
.B1(n_3146),
.B2(n_3143),
.C1(n_3145),
.C2(n_3147),
.Y(n_14590)
);

OAI221xp5_ASAP7_75t_L g14591 ( 
.A1(n_14532),
.A2(n_3147),
.B1(n_3145),
.B2(n_3146),
.C(n_3148),
.Y(n_14591)
);

AOI32xp33_ASAP7_75t_L g14592 ( 
.A1(n_14543),
.A2(n_3151),
.A3(n_3149),
.B1(n_3150),
.B2(n_3152),
.Y(n_14592)
);

OAI221xp5_ASAP7_75t_L g14593 ( 
.A1(n_14532),
.A2(n_3152),
.B1(n_3150),
.B2(n_3151),
.C(n_3153),
.Y(n_14593)
);

NOR2xp33_ASAP7_75t_L g14594 ( 
.A(n_14530),
.B(n_3153),
.Y(n_14594)
);

OAI211xp5_ASAP7_75t_L g14595 ( 
.A1(n_14532),
.A2(n_3156),
.B(n_3154),
.C(n_3155),
.Y(n_14595)
);

OAI322xp33_ASAP7_75t_L g14596 ( 
.A1(n_14530),
.A2(n_3160),
.A3(n_3159),
.B1(n_3157),
.B2(n_3154),
.C1(n_3155),
.C2(n_3158),
.Y(n_14596)
);

NOR3x1_ASAP7_75t_L g14597 ( 
.A(n_14585),
.B(n_3159),
.C(n_3158),
.Y(n_14597)
);

BUFx2_ASAP7_75t_L g14598 ( 
.A(n_14580),
.Y(n_14598)
);

NOR2xp33_ASAP7_75t_L g14599 ( 
.A(n_14576),
.B(n_3427),
.Y(n_14599)
);

AO22x2_ASAP7_75t_L g14600 ( 
.A1(n_14586),
.A2(n_3167),
.B1(n_3176),
.B2(n_3157),
.Y(n_14600)
);

OAI22x1_ASAP7_75t_L g14601 ( 
.A1(n_14588),
.A2(n_3162),
.B1(n_3160),
.B2(n_3161),
.Y(n_14601)
);

AOI22xp5_ASAP7_75t_L g14602 ( 
.A1(n_14595),
.A2(n_3163),
.B1(n_3161),
.B2(n_3162),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_14583),
.Y(n_14603)
);

AO22x2_ASAP7_75t_L g14604 ( 
.A1(n_14587),
.A2(n_14589),
.B1(n_14566),
.B2(n_14570),
.Y(n_14604)
);

XNOR2x1_ASAP7_75t_SL g14605 ( 
.A(n_14579),
.B(n_3163),
.Y(n_14605)
);

O2A1O1Ixp33_ASAP7_75t_R g14606 ( 
.A1(n_14574),
.A2(n_3166),
.B(n_3164),
.C(n_3165),
.Y(n_14606)
);

OAI22xp5_ASAP7_75t_SL g14607 ( 
.A1(n_14575),
.A2(n_3174),
.B1(n_3184),
.B2(n_3164),
.Y(n_14607)
);

INVx1_ASAP7_75t_L g14608 ( 
.A(n_14594),
.Y(n_14608)
);

OAI211xp5_ASAP7_75t_L g14609 ( 
.A1(n_14584),
.A2(n_3168),
.B(n_3165),
.C(n_3166),
.Y(n_14609)
);

XNOR2xp5_ASAP7_75t_L g14610 ( 
.A(n_14564),
.B(n_3168),
.Y(n_14610)
);

AOI22xp5_ASAP7_75t_L g14611 ( 
.A1(n_14573),
.A2(n_3172),
.B1(n_3169),
.B2(n_3170),
.Y(n_14611)
);

OR2x2_ASAP7_75t_L g14612 ( 
.A(n_14591),
.B(n_3169),
.Y(n_14612)
);

INVx1_ASAP7_75t_L g14613 ( 
.A(n_14572),
.Y(n_14613)
);

NOR3xp33_ASAP7_75t_L g14614 ( 
.A(n_14593),
.B(n_3170),
.C(n_3173),
.Y(n_14614)
);

OAI22xp5_ASAP7_75t_SL g14615 ( 
.A1(n_14568),
.A2(n_3182),
.B1(n_3191),
.B2(n_3173),
.Y(n_14615)
);

NAND2xp5_ASAP7_75t_L g14616 ( 
.A(n_14592),
.B(n_3425),
.Y(n_14616)
);

NAND2x1_ASAP7_75t_L g14617 ( 
.A(n_14569),
.B(n_3174),
.Y(n_14617)
);

INVx1_ASAP7_75t_SL g14618 ( 
.A(n_14565),
.Y(n_14618)
);

NAND4xp25_ASAP7_75t_L g14619 ( 
.A(n_14577),
.B(n_3177),
.C(n_3175),
.D(n_3176),
.Y(n_14619)
);

BUFx2_ASAP7_75t_L g14620 ( 
.A(n_14581),
.Y(n_14620)
);

AO22x2_ASAP7_75t_L g14621 ( 
.A1(n_14613),
.A2(n_14618),
.B1(n_14603),
.B2(n_14608),
.Y(n_14621)
);

INVx2_ASAP7_75t_L g14622 ( 
.A(n_14597),
.Y(n_14622)
);

INVx1_ASAP7_75t_L g14623 ( 
.A(n_14605),
.Y(n_14623)
);

XNOR2x1_ASAP7_75t_L g14624 ( 
.A(n_14604),
.B(n_14578),
.Y(n_14624)
);

INVx1_ASAP7_75t_L g14625 ( 
.A(n_14610),
.Y(n_14625)
);

NAND2xp5_ASAP7_75t_L g14626 ( 
.A(n_14614),
.B(n_14590),
.Y(n_14626)
);

OAI22xp5_ASAP7_75t_L g14627 ( 
.A1(n_14602),
.A2(n_14567),
.B1(n_14596),
.B2(n_14582),
.Y(n_14627)
);

INVx2_ASAP7_75t_L g14628 ( 
.A(n_14601),
.Y(n_14628)
);

OAI22xp5_ASAP7_75t_SL g14629 ( 
.A1(n_14617),
.A2(n_14571),
.B1(n_3178),
.B2(n_3175),
.Y(n_14629)
);

NAND2x1p5_ASAP7_75t_L g14630 ( 
.A(n_14598),
.B(n_3177),
.Y(n_14630)
);

INVx4_ASAP7_75t_L g14631 ( 
.A(n_14604),
.Y(n_14631)
);

AOI22xp5_ASAP7_75t_L g14632 ( 
.A1(n_14615),
.A2(n_3180),
.B1(n_3178),
.B2(n_3179),
.Y(n_14632)
);

AO22x2_ASAP7_75t_L g14633 ( 
.A1(n_14609),
.A2(n_3452),
.B1(n_3454),
.B2(n_3444),
.Y(n_14633)
);

INVx2_ASAP7_75t_L g14634 ( 
.A(n_14612),
.Y(n_14634)
);

NAND2xp5_ASAP7_75t_L g14635 ( 
.A(n_14619),
.B(n_3179),
.Y(n_14635)
);

INVx1_ASAP7_75t_L g14636 ( 
.A(n_14616),
.Y(n_14636)
);

OAI22xp5_ASAP7_75t_SL g14637 ( 
.A1(n_14620),
.A2(n_3184),
.B1(n_3180),
.B2(n_3182),
.Y(n_14637)
);

OAI22xp5_ASAP7_75t_L g14638 ( 
.A1(n_14632),
.A2(n_14611),
.B1(n_14606),
.B2(n_14607),
.Y(n_14638)
);

INVx1_ASAP7_75t_L g14639 ( 
.A(n_14629),
.Y(n_14639)
);

XOR2x1_ASAP7_75t_L g14640 ( 
.A(n_14624),
.B(n_14600),
.Y(n_14640)
);

OAI22x1_ASAP7_75t_L g14641 ( 
.A1(n_14631),
.A2(n_14628),
.B1(n_14622),
.B2(n_14623),
.Y(n_14641)
);

OAI22x1_ASAP7_75t_L g14642 ( 
.A1(n_14625),
.A2(n_14599),
.B1(n_14600),
.B2(n_3187),
.Y(n_14642)
);

AOI22xp5_ASAP7_75t_L g14643 ( 
.A1(n_14633),
.A2(n_3195),
.B1(n_3203),
.B2(n_3185),
.Y(n_14643)
);

XNOR2xp5_ASAP7_75t_L g14644 ( 
.A(n_14621),
.B(n_14627),
.Y(n_14644)
);

INVx1_ASAP7_75t_L g14645 ( 
.A(n_14635),
.Y(n_14645)
);

INVxp67_ASAP7_75t_L g14646 ( 
.A(n_14626),
.Y(n_14646)
);

NAND2xp5_ASAP7_75t_L g14647 ( 
.A(n_14634),
.B(n_3185),
.Y(n_14647)
);

INVx1_ASAP7_75t_L g14648 ( 
.A(n_14636),
.Y(n_14648)
);

XOR2xp5_ASAP7_75t_L g14649 ( 
.A(n_14630),
.B(n_3186),
.Y(n_14649)
);

AND2x2_ASAP7_75t_L g14650 ( 
.A(n_14637),
.B(n_3187),
.Y(n_14650)
);

HB1xp67_ASAP7_75t_L g14651 ( 
.A(n_14649),
.Y(n_14651)
);

AOI22xp5_ASAP7_75t_L g14652 ( 
.A1(n_14641),
.A2(n_3189),
.B1(n_3190),
.B2(n_3188),
.Y(n_14652)
);

INVx2_ASAP7_75t_SL g14653 ( 
.A(n_14650),
.Y(n_14653)
);

NAND2xp5_ASAP7_75t_L g14654 ( 
.A(n_14642),
.B(n_3188),
.Y(n_14654)
);

AOI22xp5_ASAP7_75t_SL g14655 ( 
.A1(n_14644),
.A2(n_3192),
.B1(n_3186),
.B2(n_3189),
.Y(n_14655)
);

INVx2_ASAP7_75t_L g14656 ( 
.A(n_14643),
.Y(n_14656)
);

AOI21xp5_ASAP7_75t_L g14657 ( 
.A1(n_14646),
.A2(n_3192),
.B(n_3193),
.Y(n_14657)
);

AOI21xp33_ASAP7_75t_SL g14658 ( 
.A1(n_14648),
.A2(n_3438),
.B(n_3437),
.Y(n_14658)
);

OAI22xp5_ASAP7_75t_SL g14659 ( 
.A1(n_14639),
.A2(n_3198),
.B1(n_3196),
.B2(n_3197),
.Y(n_14659)
);

HB1xp67_ASAP7_75t_L g14660 ( 
.A(n_14640),
.Y(n_14660)
);

AOI221x1_ASAP7_75t_L g14661 ( 
.A1(n_14645),
.A2(n_14638),
.B1(n_14647),
.B2(n_3199),
.C(n_3197),
.Y(n_14661)
);

OAI22xp5_ASAP7_75t_L g14662 ( 
.A1(n_14643),
.A2(n_3200),
.B1(n_3198),
.B2(n_3199),
.Y(n_14662)
);

INVx1_ASAP7_75t_L g14663 ( 
.A(n_14654),
.Y(n_14663)
);

INVx1_ASAP7_75t_L g14664 ( 
.A(n_14660),
.Y(n_14664)
);

AND2x4_ASAP7_75t_L g14665 ( 
.A(n_14656),
.B(n_3200),
.Y(n_14665)
);

AOI22xp33_ASAP7_75t_L g14666 ( 
.A1(n_14653),
.A2(n_3203),
.B1(n_3201),
.B2(n_3202),
.Y(n_14666)
);

AOI22xp5_ASAP7_75t_L g14667 ( 
.A1(n_14662),
.A2(n_3204),
.B1(n_3201),
.B2(n_3202),
.Y(n_14667)
);

OAI21x1_ASAP7_75t_SL g14668 ( 
.A1(n_14657),
.A2(n_3204),
.B(n_3205),
.Y(n_14668)
);

INVx1_ASAP7_75t_L g14669 ( 
.A(n_14651),
.Y(n_14669)
);

AOI22xp33_ASAP7_75t_L g14670 ( 
.A1(n_14652),
.A2(n_3208),
.B1(n_3205),
.B2(n_3206),
.Y(n_14670)
);

AOI22xp5_ASAP7_75t_L g14671 ( 
.A1(n_14664),
.A2(n_14659),
.B1(n_14661),
.B2(n_14655),
.Y(n_14671)
);

INVx1_ASAP7_75t_L g14672 ( 
.A(n_14669),
.Y(n_14672)
);

INVx1_ASAP7_75t_L g14673 ( 
.A(n_14663),
.Y(n_14673)
);

INVx1_ASAP7_75t_L g14674 ( 
.A(n_14668),
.Y(n_14674)
);

INVx1_ASAP7_75t_L g14675 ( 
.A(n_14667),
.Y(n_14675)
);

INVx1_ASAP7_75t_L g14676 ( 
.A(n_14672),
.Y(n_14676)
);

NAND2xp5_ASAP7_75t_L g14677 ( 
.A(n_14674),
.B(n_14670),
.Y(n_14677)
);

AOI21xp33_ASAP7_75t_L g14678 ( 
.A1(n_14673),
.A2(n_14658),
.B(n_14666),
.Y(n_14678)
);

NAND2xp5_ASAP7_75t_L g14679 ( 
.A(n_14671),
.B(n_14665),
.Y(n_14679)
);

AO22x2_ASAP7_75t_L g14680 ( 
.A1(n_14676),
.A2(n_14675),
.B1(n_3422),
.B2(n_3423),
.Y(n_14680)
);

OA22x2_ASAP7_75t_L g14681 ( 
.A1(n_14677),
.A2(n_3209),
.B1(n_3206),
.B2(n_3208),
.Y(n_14681)
);

AOI22xp5_ASAP7_75t_L g14682 ( 
.A1(n_14679),
.A2(n_3211),
.B1(n_3209),
.B2(n_3210),
.Y(n_14682)
);

XNOR2xp5_ASAP7_75t_L g14683 ( 
.A(n_14680),
.B(n_14678),
.Y(n_14683)
);

OA21x2_ASAP7_75t_L g14684 ( 
.A1(n_14682),
.A2(n_3212),
.B(n_3213),
.Y(n_14684)
);

OR2x6_ASAP7_75t_L g14685 ( 
.A(n_14681),
.B(n_3213),
.Y(n_14685)
);

INVx2_ASAP7_75t_SL g14686 ( 
.A(n_14683),
.Y(n_14686)
);

INVx1_ASAP7_75t_L g14687 ( 
.A(n_14685),
.Y(n_14687)
);

NAND2xp5_ASAP7_75t_L g14688 ( 
.A(n_14686),
.B(n_14684),
.Y(n_14688)
);

AOI22xp33_ASAP7_75t_SL g14689 ( 
.A1(n_14688),
.A2(n_14687),
.B1(n_3217),
.B2(n_3214),
.Y(n_14689)
);

AOI22xp5_ASAP7_75t_L g14690 ( 
.A1(n_14689),
.A2(n_3217),
.B1(n_3214),
.B2(n_3215),
.Y(n_14690)
);

AOI211xp5_ASAP7_75t_L g14691 ( 
.A1(n_14690),
.A2(n_3219),
.B(n_3215),
.C(n_3218),
.Y(n_14691)
);


endmodule