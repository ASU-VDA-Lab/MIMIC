module fake_jpeg_21257_n_310 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_25),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_19),
.B(n_17),
.C(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_25),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_40),
.B1(n_24),
.B2(n_37),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_44),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_45),
.B(n_43),
.C(n_15),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_65),
.B(n_67),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_45),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_75),
.CI(n_49),
.CON(n_87),
.SN(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_24),
.B1(n_36),
.B2(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_36),
.B1(n_41),
.B2(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_83),
.B1(n_42),
.B2(n_30),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_95),
.B(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_58),
.B1(n_56),
.B2(n_59),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_52),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_93),
.B(n_72),
.C(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_42),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_69),
.B1(n_76),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_66),
.B1(n_95),
.B2(n_71),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_108),
.B(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_72),
.B1(n_75),
.B2(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_75),
.C(n_70),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_61),
.B1(n_70),
.B2(n_39),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_61),
.B1(n_48),
.B2(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_61),
.B1(n_41),
.B2(n_36),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_32),
.C(n_33),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_20),
.B(n_13),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_20),
.B(n_13),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_92),
.B(n_78),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_94),
.B1(n_87),
.B2(n_42),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_42),
.B1(n_31),
.B2(n_28),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_119),
.B1(n_80),
.B2(n_83),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_32),
.C(n_33),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_87),
.Y(n_135)
);

OR2x4_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_15),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_76),
.B1(n_69),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_140),
.B1(n_138),
.B2(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_92),
.B(n_87),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_134),
.B(n_147),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_84),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_141),
.B(n_144),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_90),
.B1(n_86),
.B2(n_89),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_145),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_99),
.B1(n_105),
.B2(n_106),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_143),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_99),
.B1(n_110),
.B2(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_91),
.B(n_71),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_91),
.A3(n_71),
.B1(n_29),
.B2(n_35),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_109),
.B(n_116),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_157),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_158),
.B1(n_170),
.B2(n_175),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_147),
.B(n_141),
.Y(n_189)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_112),
.B1(n_108),
.B2(n_15),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_29),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_162),
.C(n_168),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_139),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_176),
.B1(n_123),
.B2(n_128),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_35),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_14),
.B1(n_17),
.B2(n_2),
.Y(n_170)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_14),
.B1(n_17),
.B2(n_2),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_71),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_131),
.C(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_151),
.B1(n_152),
.B2(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_195),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_23),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_144),
.B(n_120),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_125),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_195),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_10),
.B(n_9),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_209),
.B1(n_213),
.B2(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_177),
.C(n_168),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_211),
.C(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_163),
.B1(n_158),
.B2(n_150),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_159),
.C(n_162),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_184),
.B1(n_176),
.B2(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_187),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_150),
.B1(n_34),
.B2(n_46),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_46),
.C(n_16),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_46),
.C(n_16),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_219),
.C(n_192),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_46),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_223),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_16),
.C(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_178),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_233),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_181),
.B(n_196),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_236),
.B(n_200),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_181),
.B(n_188),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_191),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_238),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_206),
.B1(n_201),
.B2(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_179),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_211),
.C(n_203),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_223),
.C(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_213),
.B1(n_199),
.B2(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_214),
.C(n_212),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_217),
.C(n_185),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_257),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_194),
.B(n_10),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_9),
.B(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_235),
.B1(n_234),
.B2(n_236),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_226),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_252),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_0),
.B(n_2),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_12),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_272),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_16),
.C(n_23),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_258),
.B1(n_246),
.B2(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_278),
.Y(n_288)
);

AOI321xp33_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_264),
.A3(n_266),
.B1(n_269),
.B2(n_267),
.C(n_262),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_4),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_282),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_265),
.B(n_263),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_16),
.CI(n_12),
.CON(n_283),
.SN(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_0),
.B(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_16),
.C(n_23),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_291),
.C(n_294),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_293),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.C(n_283),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_276),
.B(n_4),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_5),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_5),
.B(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_292),
.C(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_300),
.B(n_288),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_297),
.B(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_305),
.C(n_286),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_5),
.B(n_6),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_7),
.B1(n_8),
.B2(n_280),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_7),
.C(n_8),
.Y(n_310)
);


endmodule