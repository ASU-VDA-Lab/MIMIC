module fake_netlist_5_476_n_2096 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2096);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2096;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_10),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_118),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_10),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_98),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_90),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_74),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_64),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_95),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_29),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_62),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_14),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_120),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_1),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_77),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_46),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_93),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_91),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_133),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_45),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_196),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_81),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_107),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_24),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_153),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_97),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_202),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_155),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_179),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_96),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_166),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_22),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_177),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_189),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_171),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_78),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_40),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_192),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_102),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_154),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_161),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_0),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_127),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_101),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_162),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_203),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_168),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_67),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_175),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_72),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_191),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_63),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_187),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_53),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_130),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_19),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_25),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_138),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_57),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_47),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_56),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_23),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_50),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_125),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_18),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_35),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_68),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_82),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_43),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_86),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_198),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_122),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_150),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_104),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_47),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_12),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_182),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_49),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_20),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_65),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_114),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_126),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_84),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_49),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_25),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_50),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_178),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_190),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_170),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_21),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_72),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_115),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_52),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_92),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_169),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_15),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_135),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_143),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_134),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_129),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_1),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_100),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_144),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_43),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_52),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_74),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_12),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_42),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_128),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_111),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_22),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_16),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_163),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_99),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_67),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_123),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_41),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_57),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_146),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_83),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_11),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_141),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_5),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_39),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_31),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_108),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_56),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_44),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_27),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_145),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_59),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_76),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_31),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_139),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_131),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_181),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_37),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_27),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_29),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_46),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_149),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_105),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_113),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_35),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_156),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_68),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_4),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_119),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_61),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_160),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_110),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_79),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_20),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_152),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_180),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_252),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_214),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_216),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_254),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_224),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_209),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_207),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_252),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_217),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_252),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_252),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_238),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_252),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_234),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_252),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_280),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_237),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_351),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_306),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_247),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_309),
.B(n_3),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_252),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_218),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_278),
.B(n_3),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_252),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_252),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_255),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_251),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_309),
.B(n_4),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_260),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_262),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_263),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_359),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_264),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_329),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_265),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g456 ( 
.A(n_218),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_272),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_274),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_276),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_284),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_344),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_344),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_212),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_344),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_344),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_317),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_286),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_344),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_317),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_255),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_211),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_298),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_357),
.B(n_5),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_339),
.B(n_6),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_212),
.B(n_6),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_298),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_288),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_289),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_349),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_292),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_207),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_324),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_293),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_349),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_295),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_361),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_223),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_361),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_207),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_297),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_230),
.B(n_7),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_299),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_321),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_223),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_258),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_230),
.B(n_7),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_326),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_207),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_327),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_207),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_339),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_258),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_259),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_244),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_259),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_220),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_331),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_336),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_266),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_453),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_486),
.A2(n_281),
.B(n_266),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_478),
.B(n_324),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_465),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_357),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_466),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_422),
.B(n_387),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_467),
.B(n_503),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_440),
.B(n_267),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_419),
.B(n_369),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_267),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_479),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_468),
.B(n_323),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_469),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_369),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_419),
.B(n_323),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_469),
.B(n_382),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_472),
.B(n_382),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_472),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_420),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_423),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_228),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_424),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

BUFx8_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_426),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_426),
.B(n_228),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_495),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_495),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_428),
.B(n_270),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_495),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_439),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_474),
.B(n_411),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_505),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_505),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_441),
.B(n_270),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_441),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_445),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_507),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_507),
.A2(n_282),
.B(n_281),
.Y(n_580)
);

CKINVDCx8_ASAP7_75t_R g581 ( 
.A(n_432),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_432),
.B(n_400),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_447),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_447),
.A2(n_308),
.B(n_282),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_467),
.B(n_240),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_437),
.B(n_253),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_448),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_474),
.B(n_337),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g593 ( 
.A1(n_451),
.A2(n_310),
.B(n_308),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_487),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_487),
.B(n_411),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_511),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_459),
.B(n_341),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_586),
.B(n_454),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_574),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_528),
.B(n_454),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_475),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_523),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_537),
.B(n_413),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_523),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_527),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_594),
.B(n_415),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_594),
.B(n_417),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_528),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_588),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_530),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_521),
.B(n_283),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_582),
.A2(n_416),
.B1(n_430),
.B2(n_427),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_532),
.B(n_433),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_594),
.B(n_442),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_574),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_532),
.B(n_444),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_581),
.Y(n_630)
);

CKINVDCx6p67_ASAP7_75t_R g631 ( 
.A(n_582),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_520),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_520),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_537),
.A2(n_414),
.B1(n_443),
.B2(n_434),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_588),
.B(n_446),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_580),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_591),
.B(n_449),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_517),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_533),
.C(n_585),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_518),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_588),
.B(n_452),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_585),
.A2(n_457),
.B1(n_458),
.B2(n_455),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_591),
.B(n_460),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_552),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_528),
.A2(n_328),
.B1(n_443),
.B2(n_434),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_539),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_588),
.B(n_533),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_598),
.B(n_463),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_525),
.B(n_482),
.C(n_471),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_568),
.B(n_387),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_517),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_581),
.B(n_483),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_539),
.A2(n_488),
.B1(n_490),
.B2(n_485),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_476),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_517),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_517),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_521),
.A2(n_477),
.B1(n_330),
.B2(n_333),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_581),
.B(n_496),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_596),
.B(n_210),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_596),
.B(n_477),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_521),
.A2(n_330),
.B1(n_333),
.B2(n_310),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_581),
.B(n_498),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_555),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_580),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_552),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_580),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_521),
.A2(n_338),
.B1(n_360),
.B2(n_334),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_518),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_552),
.B(n_208),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_580),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_568),
.A2(n_558),
.B1(n_573),
.B2(n_562),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_518),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_543),
.B(n_283),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_584),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_598),
.A2(n_513),
.B1(n_504),
.B2(n_506),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_584),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_543),
.A2(n_514),
.B1(n_515),
.B2(n_499),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_529),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_529),
.Y(n_686)
);

AO21x2_ASAP7_75t_L g687 ( 
.A1(n_587),
.A2(n_213),
.B(n_210),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_589),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_592),
.B(n_462),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_568),
.B(n_476),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_529),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_592),
.B(n_462),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_543),
.B(n_456),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_517),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_544),
.B(n_290),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_531),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_584),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_555),
.B(n_220),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_568),
.B(n_213),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_555),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_555),
.B(n_220),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_555),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_584),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_589),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_584),
.B(n_593),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_549),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_592),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_592),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_531),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_531),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_555),
.A2(n_421),
.B1(n_425),
.B2(n_418),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_589),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_592),
.A2(n_429),
.B1(n_461),
.B2(n_450),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_549),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_597),
.B(n_431),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_592),
.B(n_436),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_530),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_592),
.B(n_464),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_534),
.B(n_464),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_593),
.Y(n_726)
);

NOR2x1p5_ASAP7_75t_L g727 ( 
.A(n_541),
.B(n_312),
.Y(n_727)
);

XNOR2x2_ASAP7_75t_L g728 ( 
.A(n_541),
.B(n_334),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_558),
.A2(n_395),
.B1(n_362),
.B2(n_360),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_563),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_563),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_593),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_563),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_583),
.B(n_492),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_550),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_597),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_597),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_593),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_550),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_550),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_545),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_583),
.B(n_271),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_534),
.B(n_303),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_534),
.A2(n_379),
.B1(n_221),
.B2(n_222),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_534),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_534),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_550),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_583),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_546),
.B(n_481),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_534),
.A2(n_378),
.B1(n_375),
.B2(n_355),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_681),
.B(n_558),
.Y(n_753)
);

AND2x6_ASAP7_75t_SL g754 ( 
.A(n_605),
.B(n_338),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_607),
.B(n_583),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_618),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_708),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_681),
.A2(n_305),
.B1(n_354),
.B2(n_290),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_747),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_640),
.A2(n_558),
.B1(n_573),
.B2(n_562),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_708),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_628),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_743),
.B(n_583),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_638),
.A2(n_558),
.B1(n_573),
.B2(n_562),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_746),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_583),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_708),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_734),
.B(n_595),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_663),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_626),
.B(n_629),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_649),
.B(n_595),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_603),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_693),
.B(n_501),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_681),
.B(n_558),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_746),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_706),
.B(n_562),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_690),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_721),
.B(n_595),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_648),
.A2(n_562),
.B1(n_573),
.B2(n_544),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_713),
.B(n_225),
.C(n_215),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_603),
.Y(n_782)
);

INVxp33_ASAP7_75t_L g783 ( 
.A(n_647),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_501),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_706),
.B(n_725),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_730),
.B(n_362),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_739),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_655),
.Y(n_789)
);

BUFx6f_ASAP7_75t_SL g790 ( 
.A(n_744),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_655),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_750),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_706),
.B(n_562),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_677),
.B(n_573),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_739),
.A2(n_595),
.B(n_573),
.C(n_544),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_750),
.B(n_502),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_600),
.B(n_502),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_617),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_683),
.B(n_530),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_599),
.B(n_742),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_648),
.A2(n_544),
.B1(n_546),
.B2(n_343),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_730),
.B(n_364),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_657),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_688),
.B(n_595),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_643),
.B(n_342),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_682),
.B(n_347),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_684),
.B(n_348),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_707),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_683),
.A2(n_374),
.B1(n_384),
.B2(n_364),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_716),
.Y(n_811)
);

OR2x2_ASAP7_75t_SL g812 ( 
.A(n_698),
.B(n_374),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_699),
.B(n_530),
.Y(n_813)
);

O2A1O1Ixp5_ASAP7_75t_L g814 ( 
.A1(n_718),
.A2(n_544),
.B(n_546),
.C(n_595),
.Y(n_814)
);

AO221x1_ASAP7_75t_L g815 ( 
.A1(n_646),
.A2(n_208),
.B1(n_227),
.B2(n_385),
.C(n_384),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_699),
.B(n_530),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_723),
.B(n_530),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_604),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_723),
.B(n_530),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_726),
.B(n_736),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_726),
.B(n_736),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_619),
.B(n_530),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_732),
.B(n_604),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_608),
.B(n_548),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_749),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_608),
.B(n_548),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_620),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_623),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_620),
.B(n_548),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_712),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_622),
.B(n_548),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_622),
.A2(n_395),
.B1(n_405),
.B2(n_385),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_548),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_632),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_634),
.B(n_548),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_634),
.B(n_548),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_727),
.B(n_509),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_650),
.B(n_545),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_637),
.B(n_548),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_742),
.B(n_509),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_648),
.A2(n_544),
.B1(n_546),
.B2(n_353),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_613),
.B(n_232),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_667),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_667),
.B(n_548),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_630),
.B(n_510),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_669),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_648),
.A2(n_546),
.B1(n_356),
.B2(n_366),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_669),
.B(n_551),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_673),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_663),
.A2(n_625),
.B1(n_631),
.B2(n_744),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_673),
.B(n_551),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_676),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_663),
.A2(n_546),
.B1(n_370),
.B2(n_372),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_676),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_654),
.B(n_751),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_731),
.B(n_510),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_680),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_680),
.B(n_551),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_701),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_610),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_701),
.B(n_551),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_701),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_235),
.C(n_233),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_662),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_662),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_616),
.B(n_627),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_662),
.B(n_551),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_633),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_636),
.B(n_551),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_687),
.A2(n_405),
.B1(n_409),
.B2(n_226),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_642),
.B(n_551),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_630),
.B(n_512),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_738),
.B(n_512),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_689),
.B(n_551),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_692),
.B(n_551),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_717),
.B(n_631),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_633),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_663),
.A2(n_350),
.B1(n_376),
.B2(n_388),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_687),
.A2(n_409),
.B1(n_226),
.B2(n_301),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_712),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_624),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_744),
.A2(n_305),
.B1(n_354),
.B2(n_386),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_641),
.Y(n_885)
);

AND2x6_ASAP7_75t_SL g886 ( 
.A(n_744),
.B(n_516),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_624),
.B(n_553),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_641),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_624),
.B(n_553),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_660),
.B(n_653),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_656),
.Y(n_891)
);

INVxp33_ASAP7_75t_L g892 ( 
.A(n_714),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_535),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_687),
.A2(n_302),
.B1(n_250),
.B2(n_408),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_733),
.B(n_516),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_624),
.B(n_553),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_738),
.B(n_219),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_624),
.A2(n_397),
.B1(n_398),
.B2(n_410),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_745),
.B(n_651),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_611),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_724),
.B(n_553),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_623),
.B(n_553),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_656),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_728),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_671),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_671),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_728),
.A2(n_257),
.B1(n_219),
.B2(n_261),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_737),
.Y(n_908)
);

OAI22x1_ASAP7_75t_L g909 ( 
.A1(n_715),
.A2(n_320),
.B1(n_277),
.B2(n_275),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_624),
.B(n_553),
.Y(n_910)
);

AND2x2_ASAP7_75t_SL g911 ( 
.A(n_666),
.B(n_358),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_675),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_679),
.B(n_553),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_623),
.B(n_553),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_720),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_661),
.B(n_236),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_665),
.B(n_481),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_666),
.B(n_484),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_679),
.B(n_553),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_651),
.B(n_239),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_L g921 ( 
.A1(n_664),
.A2(n_315),
.B1(n_352),
.B2(n_304),
.C(n_294),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_675),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_756),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_776),
.Y(n_924)
);

AND2x2_ASAP7_75t_SL g925 ( 
.A(n_911),
.B(n_702),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_765),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_794),
.A2(n_821),
.B(n_775),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_895),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_774),
.B(n_679),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_771),
.B(n_679),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_791),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_791),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_861),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_819),
.B(n_835),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_758),
.A2(n_704),
.B(n_241),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_819),
.B(n_679),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_794),
.A2(n_711),
.B(n_658),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_814),
.A2(n_795),
.B(n_824),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_847),
.B(n_702),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_835),
.B(n_679),
.Y(n_940)
);

AOI21xp33_ASAP7_75t_L g941 ( 
.A1(n_843),
.A2(n_737),
.B(n_705),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_864),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_753),
.A2(n_711),
.B(n_658),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_874),
.B(n_705),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_851),
.B(n_614),
.Y(n_945)
);

O2A1O1Ixp5_ASAP7_75t_L g946 ( 
.A1(n_871),
.A2(n_639),
.B(n_652),
.C(n_614),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_755),
.A2(n_767),
.B1(n_854),
.B2(n_851),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_770),
.B(n_231),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_762),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_868),
.A2(n_697),
.B1(n_639),
.B2(n_652),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_841),
.B(n_670),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_854),
.B(n_614),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_858),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_776),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_824),
.A2(n_686),
.B(n_685),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_776),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_875),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_797),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_776),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_856),
.B(n_639),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_783),
.B(n_229),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_866),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_752),
.B(n_729),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_856),
.B(n_652),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_752),
.B(n_399),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_859),
.B(n_659),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_859),
.B(n_828),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_862),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_844),
.B(n_659),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_845),
.B(n_659),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_916),
.A2(n_250),
.B(n_246),
.C(n_256),
.Y(n_971)
);

AO21x1_ASAP7_75t_L g972 ( 
.A1(n_772),
.A2(n_241),
.B(n_231),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_800),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_753),
.A2(n_658),
.B(n_621),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_867),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_848),
.B(n_695),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_787),
.B(n_695),
.Y(n_977)
);

AOI33xp33_ASAP7_75t_L g978 ( 
.A1(n_907),
.A2(n_500),
.A3(n_494),
.B1(n_493),
.B2(n_491),
.B3(n_489),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_787),
.B(n_695),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_792),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_892),
.B(n_621),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_822),
.A2(n_827),
.B(n_777),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_798),
.B(n_697),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_868),
.B(n_401),
.Y(n_984)
);

OR2x2_ASAP7_75t_SL g985 ( 
.A(n_899),
.B(n_246),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_770),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_803),
.B(n_697),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_822),
.A2(n_748),
.B(n_686),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_809),
.B(n_697),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_786),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_775),
.A2(n_703),
.B(n_621),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_883),
.A2(n_358),
.B1(n_386),
.B2(n_392),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_786),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_862),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_900),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_808),
.B(n_703),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_900),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_777),
.A2(n_703),
.B(n_678),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_811),
.B(n_697),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_778),
.B(n_697),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_793),
.A2(n_678),
.B(n_685),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_788),
.B(n_748),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_827),
.A2(n_694),
.B(n_691),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_796),
.B(n_691),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_796),
.B(n_741),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_883),
.B(n_645),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_793),
.A2(n_696),
.B(n_694),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_808),
.B(n_696),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_916),
.A2(n_256),
.B(n_257),
.C(n_261),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_852),
.B(n_404),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_786),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_808),
.B(n_741),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_785),
.A2(n_710),
.B(n_709),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_808),
.B(n_709),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_789),
.B(n_838),
.Y(n_1015)
);

OAI22x1_ASAP7_75t_L g1016 ( 
.A1(n_904),
.A2(n_322),
.B1(n_242),
.B2(n_243),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_799),
.A2(n_817),
.B(n_813),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_790),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_826),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_815),
.A2(n_392),
.B1(n_273),
.B2(n_279),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_918),
.B(n_740),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_785),
.A2(n_719),
.B(n_710),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_825),
.A2(n_735),
.B(n_719),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_830),
.A2(n_740),
.B(n_735),
.Y(n_1024)
);

AO22x1_ASAP7_75t_L g1025 ( 
.A1(n_843),
.A2(n_318),
.B1(n_291),
.B2(n_287),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_832),
.A2(n_612),
.B(n_611),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_894),
.A2(n_273),
.B1(n_407),
.B2(n_391),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_917),
.B(n_601),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_406),
.B1(n_674),
.B2(n_623),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_784),
.B(n_601),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_799),
.A2(n_606),
.B(n_602),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_870),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_773),
.B(n_245),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_831),
.Y(n_1034)
);

AO21x1_ASAP7_75t_L g1035 ( 
.A1(n_871),
.A2(n_279),
.B(n_269),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_834),
.A2(n_615),
.B(n_612),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_757),
.B(n_602),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_836),
.A2(n_615),
.B(n_609),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_831),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_766),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_812),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_911),
.B(n_674),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_757),
.B(n_606),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_921),
.B(n_285),
.C(n_269),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_879),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_837),
.A2(n_609),
.B(n_672),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_759),
.B(n_674),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_873),
.A2(n_722),
.B(n_674),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_761),
.B(n_674),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_831),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_915),
.B(n_722),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_813),
.A2(n_566),
.B(n_559),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_817),
.A2(n_566),
.B(n_559),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_840),
.A2(n_672),
.B(n_566),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_831),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_820),
.A2(n_566),
.B(n_559),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_846),
.A2(n_570),
.B(n_559),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_761),
.B(n_722),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_873),
.A2(n_722),
.B(n_517),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_768),
.B(n_722),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_850),
.A2(n_668),
.B(n_645),
.Y(n_1061)
);

NOR2x2_ASAP7_75t_L g1062 ( 
.A(n_897),
.B(n_220),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_885),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_853),
.A2(n_860),
.B(n_818),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_890),
.A2(n_407),
.B(n_391),
.C(n_335),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_768),
.B(n_570),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_779),
.A2(n_820),
.B(n_863),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_782),
.B(n_248),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_770),
.B(n_908),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_769),
.B(n_570),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_880),
.B(n_668),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_760),
.A2(n_570),
.B(n_576),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_888),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_833),
.B(n_575),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_920),
.A2(n_780),
.B(n_857),
.C(n_764),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_894),
.A2(n_881),
.B1(n_801),
.B2(n_842),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_763),
.A2(n_590),
.B(n_575),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_L g1079 ( 
.A(n_800),
.B(n_865),
.C(n_878),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_891),
.Y(n_1080)
);

AND2x2_ASAP7_75t_SL g1081 ( 
.A(n_907),
.B(n_285),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_863),
.A2(n_576),
.B(n_575),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_833),
.B(n_575),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_920),
.B(n_249),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_810),
.B(n_576),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_806),
.A2(n_805),
.B(n_884),
.C(n_807),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_810),
.B(n_881),
.Y(n_1087)
);

OAI321xp33_ASAP7_75t_L g1088 ( 
.A1(n_872),
.A2(n_390),
.A3(n_408),
.B1(n_301),
.B2(n_302),
.C(n_325),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_872),
.A2(n_325),
.B1(n_335),
.B2(n_390),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_855),
.B(n_208),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_849),
.A2(n_590),
.B(n_576),
.C(n_577),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_869),
.A2(n_577),
.B1(n_590),
.B2(n_552),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_922),
.B(n_577),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_804),
.A2(n_590),
.B(n_577),
.C(n_536),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_905),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_906),
.Y(n_1097)
);

AND2x6_ASAP7_75t_L g1098 ( 
.A(n_887),
.B(n_208),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_869),
.A2(n_524),
.B(n_557),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_781),
.B(n_897),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_912),
.B(n_557),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_889),
.A2(n_524),
.B(n_557),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_897),
.B(n_268),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_902),
.A2(n_542),
.B(n_540),
.C(n_519),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_882),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_882),
.B(n_557),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_882),
.B(n_557),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_802),
.B(n_296),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_816),
.B(n_557),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_896),
.A2(n_524),
.B(n_557),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_910),
.A2(n_524),
.B(n_557),
.Y(n_1111)
);

AND2x6_ASAP7_75t_L g1112 ( 
.A(n_913),
.B(n_208),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_919),
.A2(n_552),
.B(n_535),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_893),
.A2(n_535),
.B(n_536),
.C(n_522),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1076),
.A2(n_898),
.B(n_823),
.C(n_901),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_973),
.B(n_1084),
.Y(n_1116)
);

AO32x1_ASAP7_75t_L g1117 ( 
.A1(n_1089),
.A2(n_484),
.A3(n_489),
.B1(n_491),
.B2(n_493),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1044),
.A2(n_802),
.B(n_876),
.C(n_877),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_927),
.A2(n_901),
.B(n_877),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1077),
.A2(n_876),
.B(n_914),
.C(n_902),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_961),
.B(n_307),
.C(n_300),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1081),
.A2(n_802),
.B1(n_909),
.B2(n_227),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_923),
.B(n_958),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_929),
.A2(n_829),
.B(n_914),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_928),
.B(n_886),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1015),
.B(n_519),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_953),
.B(n_754),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_927),
.A2(n_947),
.B(n_1064),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_949),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_926),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_1018),
.B(n_311),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_941),
.A2(n_519),
.B(n_542),
.C(n_540),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_935),
.A2(n_522),
.B(n_526),
.C(n_538),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1049),
.A2(n_668),
.B(n_645),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_980),
.B(n_522),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_925),
.B(n_313),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_981),
.B(n_526),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_956),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1050),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_933),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_982),
.A2(n_227),
.B1(n_314),
.B2(n_316),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_L g1142 ( 
.A(n_986),
.B(n_526),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_951),
.B(n_538),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_938),
.A2(n_524),
.B(n_557),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1067),
.A2(n_524),
.B(n_565),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_986),
.B(n_319),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1021),
.B(n_538),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1058),
.A2(n_1060),
.B(n_991),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_974),
.A2(n_668),
.B(n_645),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1030),
.B(n_540),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_942),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1041),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_962),
.B(n_542),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_975),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1019),
.B(n_547),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_L g1156 ( 
.A(n_1025),
.B(n_381),
.C(n_380),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_971),
.A2(n_547),
.B(n_579),
.C(n_572),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_931),
.B(n_547),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1079),
.B(n_332),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_932),
.B(n_565),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_957),
.B(n_340),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1028),
.B(n_565),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1009),
.A2(n_500),
.B(n_494),
.C(n_535),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1002),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_956),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1011),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_985),
.B(n_345),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1033),
.B(n_346),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_L g1169 ( 
.A1(n_972),
.A2(n_571),
.B(n_579),
.C(n_556),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_990),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_1040),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1103),
.B(n_363),
.C(n_367),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_954),
.B(n_956),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1067),
.B(n_565),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_974),
.A2(n_668),
.B(n_645),
.Y(n_1175)
);

HAxp5_ASAP7_75t_L g1176 ( 
.A(n_1062),
.B(n_368),
.CON(n_1176),
.SN(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1010),
.A2(n_536),
.B(n_535),
.C(n_572),
.Y(n_1177)
);

NAND2x1_ASAP7_75t_L g1178 ( 
.A(n_1050),
.B(n_535),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1073),
.A2(n_524),
.B(n_567),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_984),
.B(n_565),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1068),
.B(n_371),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_930),
.A2(n_579),
.B(n_556),
.C(n_572),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_954),
.B(n_377),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1042),
.A2(n_560),
.B(n_571),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_924),
.B(n_565),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_939),
.B(n_383),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_924),
.B(n_565),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_959),
.B(n_565),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1108),
.B(n_393),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1086),
.A2(n_394),
.B(n_396),
.C(n_403),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_993),
.B(n_536),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_968),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_944),
.B(n_8),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_1016),
.B(n_85),
.Y(n_1194)
);

CKINVDCx6p67_ASAP7_75t_R g1195 ( 
.A(n_1069),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_994),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_959),
.B(n_565),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_963),
.B(n_567),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1100),
.B(n_8),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_1090),
.A2(n_560),
.B(n_571),
.C(n_569),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1050),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1100),
.A2(n_227),
.B1(n_552),
.B2(n_536),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_965),
.B(n_569),
.C(n_560),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_948),
.B(n_536),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_991),
.A2(n_524),
.B(n_567),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1069),
.B(n_948),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1017),
.B(n_567),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1071),
.A2(n_524),
.B(n_567),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_948),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_995),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1031),
.A2(n_556),
.B(n_569),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_936),
.A2(n_567),
.B(n_578),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_997),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1032),
.A2(n_1096),
.B1(n_1074),
.B2(n_1095),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1020),
.A2(n_578),
.B(n_564),
.C(n_561),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1069),
.Y(n_1216)
);

AND2x2_ASAP7_75t_SL g1217 ( 
.A(n_978),
.B(n_9),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1063),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1080),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1065),
.A2(n_578),
.B(n_564),
.C(n_561),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1088),
.A2(n_578),
.B(n_564),
.C(n_561),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1039),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_940),
.A2(n_567),
.B(n_578),
.Y(n_1223)
);

CKINVDCx16_ASAP7_75t_R g1224 ( 
.A(n_1070),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1070),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1070),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1039),
.B(n_1105),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1034),
.B(n_157),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_967),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_992),
.A2(n_1047),
.B(n_1091),
.C(n_1005),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1039),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1078),
.A2(n_578),
.B(n_564),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1097),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1013),
.A2(n_552),
.B(n_561),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_R g1235 ( 
.A(n_1034),
.B(n_1055),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1045),
.A2(n_552),
.B1(n_561),
.B2(n_554),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1000),
.A2(n_552),
.B1(n_561),
.B2(n_554),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1004),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1093),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1055),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_937),
.A2(n_564),
.B(n_554),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_937),
.A2(n_564),
.B(n_554),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_934),
.A2(n_554),
.B(n_552),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1094),
.A2(n_554),
.B(n_11),
.C(n_13),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1013),
.A2(n_552),
.B(n_204),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1035),
.A2(n_552),
.B1(n_13),
.B2(n_17),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1066),
.A2(n_140),
.B(n_197),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1105),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1008),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_9),
.B(n_17),
.C(n_19),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1105),
.A2(n_200),
.B(n_193),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1029),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_R g1253 ( 
.A(n_1105),
.B(n_183),
.Y(n_1253)
);

OR2x6_ASAP7_75t_SL g1254 ( 
.A(n_983),
.B(n_21),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_950),
.A2(n_167),
.B1(n_165),
.B2(n_151),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1037),
.B(n_24),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1012),
.A2(n_147),
.B(n_137),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1014),
.A2(n_124),
.B(n_112),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1043),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1006),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1104),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1098),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_945),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_969),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_SL g1265 ( 
.A(n_987),
.B(n_26),
.C(n_28),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_943),
.A2(n_103),
.B(n_94),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_943),
.A2(n_88),
.B(n_87),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_952),
.B(n_30),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_989),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_970),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1098),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1054),
.A2(n_32),
.B(n_33),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_999),
.B(n_36),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1072),
.A2(n_38),
.B1(n_40),
.B2(n_48),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1140),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1116),
.A2(n_946),
.B(n_1054),
.C(n_1075),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1151),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1129),
.B(n_996),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_L g1279 ( 
.A1(n_1168),
.A2(n_1022),
.B(n_1048),
.C(n_1024),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1206),
.B(n_1106),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1128),
.A2(n_998),
.B(n_1107),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1170),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

OAI22x1_ASAP7_75t_L g1284 ( 
.A1(n_1199),
.A2(n_1085),
.B1(n_1083),
.B2(n_1053),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1128),
.A2(n_1022),
.B(n_1057),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1148),
.A2(n_998),
.B(n_1109),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1164),
.B(n_1057),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_L g1288 ( 
.A1(n_1181),
.A2(n_1024),
.B(n_1023),
.C(n_1007),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1218),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1190),
.A2(n_976),
.B(n_966),
.C(n_964),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1165),
.B(n_1092),
.Y(n_1292)
);

NOR4xp25_ASAP7_75t_L g1293 ( 
.A(n_1250),
.B(n_955),
.C(n_1003),
.D(n_988),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1133),
.A2(n_1023),
.B(n_1026),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1115),
.A2(n_1144),
.A3(n_1120),
.B(n_1174),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1152),
.Y(n_1297)
);

BUFx10_ASAP7_75t_L g1298 ( 
.A(n_1127),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1118),
.A2(n_1001),
.B(n_1046),
.C(n_1007),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1145),
.A2(n_1036),
.B(n_1026),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1145),
.A2(n_1036),
.B(n_1038),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1249),
.B(n_960),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1144),
.A2(n_1038),
.B(n_1046),
.Y(n_1303)
);

AOI211x1_ASAP7_75t_L g1304 ( 
.A1(n_1272),
.A2(n_1052),
.B(n_1056),
.C(n_1082),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1119),
.A2(n_977),
.B(n_979),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1124),
.A2(n_1001),
.B(n_1059),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1238),
.B(n_1082),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1154),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1219),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1259),
.B(n_1112),
.Y(n_1310)
);

AOI221xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1122),
.A2(n_1099),
.B1(n_1102),
.B2(n_1111),
.C(n_1110),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1131),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1233),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1124),
.A2(n_1162),
.B(n_1137),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1167),
.A2(n_1113),
.B1(n_1099),
.B2(n_1101),
.C(n_1061),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1159),
.A2(n_1112),
.B(n_1098),
.C(n_1006),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1172),
.A2(n_38),
.B(n_48),
.C(n_51),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1207),
.A2(n_1112),
.B(n_1098),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1252),
.A2(n_1112),
.B1(n_1098),
.B2(n_54),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1189),
.B(n_1112),
.Y(n_1321)
);

INVx3_ASAP7_75t_R g1322 ( 
.A(n_1206),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1179),
.A2(n_51),
.A3(n_53),
.B(n_55),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1230),
.A2(n_58),
.B(n_60),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1165),
.B(n_58),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1254),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1143),
.B(n_75),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1216),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1245),
.A2(n_61),
.B(n_62),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1272),
.A2(n_63),
.A3(n_64),
.B(n_65),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_SL g1331 ( 
.A1(n_1273),
.A2(n_66),
.B(n_69),
.C(n_70),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1191),
.B(n_66),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1224),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1261),
.A2(n_69),
.A3(n_70),
.B(n_71),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1229),
.A2(n_71),
.B(n_73),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1192),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1264),
.B(n_73),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_75),
.B(n_1242),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1121),
.C(n_1274),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_SL g1340 ( 
.A(n_1253),
.B(n_1231),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1240),
.B(n_1166),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1196),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1150),
.A2(n_1222),
.B(n_1180),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1209),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1186),
.A2(n_1194),
.B(n_1171),
.C(n_1270),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1266),
.A2(n_1267),
.A3(n_1232),
.B(n_1241),
.Y(n_1346)
);

AO32x2_ASAP7_75t_L g1347 ( 
.A1(n_1269),
.A2(n_1141),
.A3(n_1255),
.B1(n_1117),
.B2(n_1222),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1203),
.A2(n_1256),
.B(n_1244),
.C(n_1268),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1147),
.A2(n_1198),
.B(n_1208),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1208),
.A2(n_1239),
.B(n_1227),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1138),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1210),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1126),
.A2(n_1263),
.B(n_1149),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1213),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1195),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1158),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1135),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1204),
.B(n_1228),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1175),
.A2(n_1188),
.B(n_1187),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1242),
.A2(n_1223),
.A3(n_1212),
.B(n_1247),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1155),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1214),
.B(n_1217),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1169),
.A2(n_1212),
.B(n_1223),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1153),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1247),
.A2(n_1258),
.A3(n_1257),
.B(n_1160),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1156),
.A2(n_1257),
.B(n_1258),
.C(n_1132),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1184),
.A2(n_1197),
.B(n_1185),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1215),
.A2(n_1183),
.B(n_1173),
.C(n_1265),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1138),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1176),
.B(n_1161),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

AOI221xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1246),
.A2(n_1202),
.B1(n_1163),
.B2(n_1221),
.C(n_1243),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1146),
.B(n_1139),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1231),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1201),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1237),
.A2(n_1177),
.B(n_1182),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1139),
.A2(n_1117),
.B1(n_1251),
.B2(n_1178),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1248),
.A2(n_1165),
.B1(n_1260),
.B2(n_1231),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1201),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1134),
.A2(n_1117),
.B(n_1260),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1201),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1142),
.A2(n_1220),
.B(n_1236),
.C(n_1260),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1225),
.A2(n_1226),
.B(n_1200),
.C(n_1157),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1226),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1235),
.A2(n_1262),
.B(n_1271),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1116),
.B(n_847),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1140),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1116),
.B(n_774),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1116),
.A2(n_1076),
.B1(n_1087),
.B2(n_925),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1394)
);

NOR2x1_ASAP7_75t_SL g1395 ( 
.A(n_1222),
.B(n_1231),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1138),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1128),
.A2(n_972),
.A3(n_935),
.B(n_1035),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1116),
.A2(n_1084),
.B(n_1076),
.C(n_605),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1168),
.A2(n_605),
.B(n_1084),
.C(n_1181),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1116),
.A2(n_1084),
.B(n_1076),
.C(n_605),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1165),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1116),
.B(n_630),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1129),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1133),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1129),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1116),
.B(n_973),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1116),
.B(n_774),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_1148),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1218),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1116),
.B(n_630),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1115),
.A2(n_1076),
.B(n_1120),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1129),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1234),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1130),
.B(n_618),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1129),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1190),
.A2(n_1076),
.B(n_1087),
.C(n_700),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1116),
.B(n_973),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_SL g1426 ( 
.A(n_1231),
.B(n_666),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1252),
.A2(n_1044),
.B1(n_605),
.B2(n_1084),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1253),
.B(n_630),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1122),
.A2(n_1087),
.B1(n_1027),
.B2(n_1081),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_SL g1430 ( 
.A(n_1231),
.B(n_666),
.Y(n_1430)
);

AOI221x1_ASAP7_75t_L g1431 ( 
.A1(n_1128),
.A2(n_1084),
.B1(n_1190),
.B2(n_1077),
.C(n_1272),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1116),
.A2(n_1084),
.B(n_1076),
.C(n_605),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1128),
.A2(n_972),
.A3(n_935),
.B(n_1035),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1128),
.A2(n_972),
.A3(n_935),
.B(n_1035),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1116),
.B(n_774),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1140),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1076),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1274),
.A2(n_1077),
.B1(n_904),
.B2(n_1044),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1116),
.A2(n_1084),
.B(n_1076),
.C(n_605),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1401),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1427),
.A2(n_1399),
.B1(n_1400),
.B2(n_1439),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1297),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1415),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1429),
.A2(n_1417),
.B1(n_1393),
.B2(n_1438),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1429),
.B2(n_1417),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1407),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1275),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1422),
.Y(n_1448)
);

CKINVDCx6p67_ASAP7_75t_R g1449 ( 
.A(n_1333),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1407),
.Y(n_1450)
);

INVx6_ASAP7_75t_SL g1451 ( 
.A(n_1341),
.Y(n_1451)
);

BUFx4_ASAP7_75t_SL g1452 ( 
.A(n_1403),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1418),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1282),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1277),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1312),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1344),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1308),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1320),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1392),
.B(n_1411),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1309),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1298),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1298),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1380),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1383),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1326),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1421),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1328),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1435),
.B(n_1388),
.Y(n_1469)
);

CKINVDCx6p67_ASAP7_75t_R g1470 ( 
.A(n_1355),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1398),
.A2(n_1432),
.B1(n_1409),
.B2(n_1425),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1335),
.A2(n_1362),
.B1(n_1327),
.B2(n_1319),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1322),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1370),
.A2(n_1416),
.B1(n_1402),
.B2(n_1428),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1341),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1357),
.A2(n_1364),
.B1(n_1361),
.B2(n_1356),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1313),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1324),
.A2(n_1337),
.B1(n_1332),
.B2(n_1336),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1390),
.A2(n_1437),
.B1(n_1419),
.B2(n_1406),
.Y(n_1479)
);

INVx3_ASAP7_75t_SL g1480 ( 
.A(n_1376),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1290),
.Y(n_1481)
);

INVx6_ASAP7_75t_L g1482 ( 
.A(n_1380),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1391),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1436),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1342),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1339),
.A2(n_1317),
.B(n_1431),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1352),
.A2(n_1354),
.B1(n_1371),
.B2(n_1358),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1320),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1320),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1369),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1369),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1369),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1358),
.B(n_1280),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1287),
.A2(n_1394),
.B1(n_1423),
.B2(n_1410),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1405),
.A2(n_1280),
.B1(n_1302),
.B2(n_1284),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1382),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1338),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1307),
.A2(n_1321),
.B1(n_1315),
.B2(n_1325),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1351),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1360),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1375),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1283),
.A2(n_1373),
.B1(n_1377),
.B2(n_1292),
.Y(n_1502)
);

CKINVDCx11_ASAP7_75t_R g1503 ( 
.A(n_1375),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1345),
.A2(n_1366),
.B(n_1348),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1278),
.A2(n_1343),
.B(n_1384),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1377),
.A2(n_1424),
.B1(n_1329),
.B2(n_1379),
.Y(n_1506)
);

INVx4_ASAP7_75t_SL g1507 ( 
.A(n_1330),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1375),
.Y(n_1508)
);

CKINVDCx6p67_ASAP7_75t_R g1509 ( 
.A(n_1396),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1325),
.A2(n_1310),
.B1(n_1353),
.B2(n_1351),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_R g1511 ( 
.A1(n_1386),
.A2(n_1374),
.B1(n_1331),
.B2(n_1334),
.Y(n_1511)
);

BUFx8_ASAP7_75t_L g1512 ( 
.A(n_1396),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1396),
.Y(n_1513)
);

BUFx12f_ASAP7_75t_L g1514 ( 
.A(n_1340),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1515)
);

CKINVDCx14_ASAP7_75t_R g1516 ( 
.A(n_1387),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1395),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1314),
.A2(n_1426),
.B1(n_1430),
.B2(n_1349),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1330),
.Y(n_1519)
);

CKINVDCx6p67_ASAP7_75t_R g1520 ( 
.A(n_1334),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1350),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1363),
.A2(n_1404),
.B1(n_1303),
.B2(n_1285),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1363),
.Y(n_1523)
);

CKINVDCx6p67_ASAP7_75t_R g1524 ( 
.A(n_1323),
.Y(n_1524)
);

OAI21xp33_ASAP7_75t_L g1525 ( 
.A1(n_1276),
.A2(n_1293),
.B(n_1299),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1323),
.Y(n_1526)
);

INVx6_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1378),
.A2(n_1318),
.B1(n_1404),
.B2(n_1305),
.Y(n_1528)
);

CKINVDCx11_ASAP7_75t_R g1529 ( 
.A(n_1368),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1378),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1296),
.B(n_1311),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1311),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1303),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1381),
.Y(n_1534)
);

INVx6_ASAP7_75t_L g1535 ( 
.A(n_1316),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1367),
.Y(n_1536)
);

BUFx8_ASAP7_75t_L g1537 ( 
.A(n_1347),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1285),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1372),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1372),
.Y(n_1540)
);

BUFx10_ASAP7_75t_L g1541 ( 
.A(n_1291),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1296),
.B(n_1365),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1295),
.A2(n_1281),
.B1(n_1306),
.B2(n_1359),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1295),
.A2(n_1301),
.B1(n_1300),
.B2(n_1286),
.Y(n_1544)
);

INVx4_ASAP7_75t_SL g1545 ( 
.A(n_1397),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1279),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1414),
.A2(n_1347),
.B(n_1293),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1304),
.A2(n_1347),
.B1(n_1434),
.B2(n_1397),
.Y(n_1548)
);

CKINVDCx11_ASAP7_75t_R g1549 ( 
.A(n_1304),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1294),
.A2(n_1408),
.B1(n_1420),
.B2(n_1413),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1397),
.A2(n_1433),
.B1(n_1434),
.B2(n_1365),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1389),
.A2(n_1412),
.B1(n_1288),
.B2(n_1433),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1433),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1434),
.A2(n_1427),
.B1(n_1044),
.B2(n_1417),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1346),
.B(n_1388),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1346),
.A2(n_1429),
.B1(n_1417),
.B2(n_904),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1407),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1401),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1427),
.A2(n_1399),
.B(n_605),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1427),
.A2(n_904),
.B1(n_1411),
.B2(n_1392),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1320),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1401),
.Y(n_1565)
);

CKINVDCx11_ASAP7_75t_R g1566 ( 
.A(n_1297),
.Y(n_1566)
);

BUFx10_ASAP7_75t_L g1567 ( 
.A(n_1312),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1289),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1427),
.A2(n_1399),
.B1(n_1400),
.B2(n_1398),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1427),
.A2(n_1084),
.B1(n_605),
.B2(n_421),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1320),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1289),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1427),
.A2(n_1044),
.B1(n_1417),
.B2(n_1393),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1388),
.B(n_973),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1289),
.Y(n_1578)
);

INVx6_ASAP7_75t_L g1579 ( 
.A(n_1418),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1297),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1427),
.A2(n_1399),
.B1(n_1400),
.B2(n_1398),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1427),
.A2(n_1399),
.B1(n_1400),
.B2(n_1398),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1418),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1289),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1429),
.A2(n_1417),
.B1(n_904),
.B2(n_1077),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1427),
.A2(n_1084),
.B1(n_605),
.B2(n_421),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1289),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1526),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1547),
.A2(n_1525),
.B(n_1528),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1447),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1572),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1446),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1515),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1455),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1507),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1467),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1512),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1458),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1507),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1450),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1504),
.B(n_1519),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1507),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1460),
.B(n_1469),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1529),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1586),
.A2(n_1570),
.B1(n_1441),
.B2(n_1581),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1500),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1454),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1523),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1461),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1500),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1477),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_1531),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1557),
.Y(n_1614)
);

INVxp33_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1464),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1483),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1582),
.A2(n_1560),
.B1(n_1569),
.B2(n_1576),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1465),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1484),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1444),
.B(n_1445),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1444),
.B(n_1549),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1486),
.A2(n_1510),
.B(n_1542),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1464),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1485),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1538),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1536),
.B(n_1545),
.Y(n_1627)
);

AND2x2_ASAP7_75t_SL g1628 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1464),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1558),
.A2(n_1562),
.B(n_1576),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1532),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1534),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1457),
.Y(n_1633)
);

AOI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1471),
.A2(n_1563),
.B(n_1474),
.C(n_1480),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1520),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1497),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1497),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1544),
.A2(n_1550),
.B(n_1543),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1512),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1533),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1524),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1551),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1552),
.A2(n_1522),
.B(n_1546),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1550),
.A2(n_1522),
.B(n_1494),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1556),
.B(n_1554),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1482),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1488),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1482),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1562),
.A2(n_1569),
.B1(n_1571),
.B2(n_1573),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1587),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1481),
.B(n_1448),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1568),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1556),
.B(n_1554),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1548),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1571),
.A2(n_1573),
.B1(n_1585),
.B2(n_1476),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1482),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1575),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1585),
.A2(n_1539),
.B1(n_1540),
.B2(n_1563),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1476),
.B(n_1443),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1578),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1495),
.B(n_1530),
.Y(n_1661)
);

AO21x2_ASAP7_75t_L g1662 ( 
.A1(n_1510),
.A2(n_1505),
.B(n_1584),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1496),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1535),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1521),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1535),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1535),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1541),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1494),
.A2(n_1518),
.B(n_1495),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1440),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1671)
);

AO21x2_ASAP7_75t_L g1672 ( 
.A1(n_1541),
.A2(n_1479),
.B(n_1506),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1527),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1537),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1566),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1527),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1527),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1511),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1506),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1475),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1517),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1498),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1472),
.B(n_1487),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1502),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1478),
.A2(n_1518),
.B(n_1502),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1487),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1490),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1499),
.B(n_1463),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1452),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1516),
.A2(n_1559),
.B(n_1442),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1452),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1459),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1565),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1462),
.A2(n_1453),
.B(n_1503),
.C(n_1473),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1449),
.B(n_1491),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1514),
.B(n_1565),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1491),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1491),
.B(n_1508),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1609),
.B(n_1661),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1609),
.B(n_1513),
.Y(n_1701)
);

NOR2xp67_ASAP7_75t_SL g1702 ( 
.A(n_1605),
.B(n_1579),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1661),
.B(n_1508),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1628),
.A2(n_1579),
.B1(n_1583),
.B2(n_1451),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_SL g1705 ( 
.A1(n_1634),
.A2(n_1580),
.B(n_1451),
.C(n_1509),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1674),
.B(n_1508),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1649),
.A2(n_1466),
.B1(n_1489),
.B2(n_1508),
.C(n_1574),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1630),
.A2(n_1564),
.B1(n_1574),
.B2(n_1470),
.C(n_1583),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1628),
.A2(n_1583),
.B1(n_1579),
.B2(n_1456),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1679),
.B(n_1574),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1592),
.A2(n_1492),
.B1(n_1501),
.B2(n_1567),
.Y(n_1711)
);

INVx5_ASAP7_75t_SL g1712 ( 
.A(n_1697),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1675),
.Y(n_1713)
);

OR2x6_ASAP7_75t_L g1714 ( 
.A(n_1602),
.B(n_1564),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1679),
.B(n_1574),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1606),
.A2(n_1492),
.B1(n_1567),
.B2(n_1658),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1631),
.B(n_1492),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1618),
.A2(n_1628),
.B(n_1686),
.C(n_1655),
.Y(n_1718)
);

AO32x2_ASAP7_75t_L g1719 ( 
.A1(n_1594),
.A2(n_1613),
.A3(n_1670),
.B1(n_1654),
.B2(n_1623),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1632),
.B(n_1615),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_R g1721 ( 
.A(n_1691),
.B(n_1622),
.Y(n_1721)
);

AOI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1618),
.A2(n_1621),
.B1(n_1683),
.B2(n_1677),
.C(n_1622),
.Y(n_1722)
);

AO32x2_ASAP7_75t_L g1723 ( 
.A1(n_1594),
.A2(n_1613),
.A3(n_1670),
.B1(n_1654),
.B2(n_1623),
.Y(n_1723)
);

CKINVDCx16_ASAP7_75t_R g1724 ( 
.A(n_1605),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_SL g1725 ( 
.A1(n_1695),
.A2(n_1681),
.B(n_1668),
.C(n_1673),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1626),
.B(n_1591),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_SL g1727 ( 
.A(n_1602),
.B(n_1662),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1619),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1632),
.B(n_1665),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_R g1730 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1602),
.A2(n_1684),
.B1(n_1677),
.B2(n_1683),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1591),
.B(n_1595),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1650),
.B(n_1633),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1645),
.A2(n_1653),
.B1(n_1604),
.B2(n_1685),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1627),
.B(n_1641),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1599),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1610),
.B(n_1612),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_SL g1738 ( 
.A(n_1602),
.B(n_1662),
.Y(n_1738)
);

AO32x2_ASAP7_75t_L g1739 ( 
.A1(n_1670),
.A2(n_1623),
.A3(n_1590),
.B1(n_1629),
.B2(n_1648),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_SL g1740 ( 
.A1(n_1668),
.A2(n_1673),
.B(n_1678),
.C(n_1676),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1669),
.A2(n_1684),
.B(n_1685),
.C(n_1680),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1602),
.B(n_1691),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1691),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1638),
.A2(n_1644),
.B(n_1642),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1636),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1664),
.B(n_1666),
.Y(n_1746)
);

BUFx4f_ASAP7_75t_SL g1747 ( 
.A(n_1605),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1617),
.B(n_1620),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1625),
.B(n_1699),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_L g1750 ( 
.A(n_1605),
.B(n_1690),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_R g1751 ( 
.A(n_1643),
.B(n_1590),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1607),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1687),
.A2(n_1597),
.B1(n_1614),
.B2(n_1601),
.C(n_1593),
.Y(n_1753)
);

AO32x2_ASAP7_75t_L g1754 ( 
.A1(n_1590),
.A2(n_1629),
.A3(n_1616),
.B1(n_1624),
.B2(n_1646),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1589),
.Y(n_1755)
);

OAI21x1_ASAP7_75t_SL g1756 ( 
.A1(n_1659),
.A2(n_1635),
.B(n_1667),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1588),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1635),
.B(n_1589),
.Y(n_1758)
);

AO21x2_ASAP7_75t_L g1759 ( 
.A1(n_1596),
.A2(n_1600),
.B(n_1603),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1607),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1611),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1652),
.B(n_1657),
.Y(n_1762)
);

BUFx12f_ASAP7_75t_L g1763 ( 
.A(n_1690),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1667),
.A2(n_1678),
.B(n_1676),
.C(n_1687),
.Y(n_1764)
);

AND2x4_ASAP7_75t_SL g1765 ( 
.A(n_1605),
.B(n_1697),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1660),
.B(n_1693),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1660),
.B(n_1693),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1608),
.A2(n_1590),
.B(n_1663),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1714),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1757),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1736),
.Y(n_1771)
);

NOR2xp67_ASAP7_75t_L g1772 ( 
.A(n_1745),
.B(n_1637),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1754),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1643),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1722),
.A2(n_1716),
.B1(n_1734),
.B2(n_1753),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1744),
.B(n_1643),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1754),
.B(n_1643),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1748),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1719),
.B(n_1723),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1752),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1752),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1732),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1754),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1718),
.B(n_1668),
.Y(n_1784)
);

INVx5_ASAP7_75t_SL g1785 ( 
.A(n_1742),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1754),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1737),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1743),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1722),
.A2(n_1672),
.B1(n_1662),
.B2(n_1689),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1760),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1762),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1719),
.B(n_1723),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1760),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1742),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1761),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1761),
.Y(n_1796)
);

OAI221xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1753),
.A2(n_1689),
.B1(n_1639),
.B2(n_1598),
.C(n_1697),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1759),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1731),
.A2(n_1672),
.B1(n_1671),
.B2(n_1639),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1768),
.B(n_1726),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1735),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1709),
.A2(n_1672),
.B1(n_1720),
.B2(n_1707),
.Y(n_1803)
);

INVxp67_ASAP7_75t_SL g1804 ( 
.A(n_1751),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1766),
.Y(n_1805)
);

CKINVDCx14_ASAP7_75t_R g1806 ( 
.A(n_1713),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1741),
.B(n_1640),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1781),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1804),
.B(n_1728),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1772),
.Y(n_1811)
);

AND2x2_ASAP7_75t_SL g1812 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1802),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1794),
.B(n_1742),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1778),
.B(n_1733),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1807),
.B(n_1729),
.Y(n_1816)
);

AO31x2_ASAP7_75t_L g1817 ( 
.A1(n_1773),
.A2(n_1738),
.A3(n_1727),
.B(n_1588),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1770),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1777),
.A2(n_1747),
.B1(n_1765),
.B2(n_1712),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1805),
.B(n_1791),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1795),
.Y(n_1821)
);

NAND2x1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.B(n_1756),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1777),
.A2(n_1747),
.B1(n_1712),
.B2(n_1724),
.Y(n_1823)
);

AOI33xp33_ASAP7_75t_L g1824 ( 
.A1(n_1775),
.A2(n_1709),
.A3(n_1725),
.B1(n_1700),
.B2(n_1704),
.B3(n_1701),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1795),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1788),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1795),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1794),
.B(n_1758),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1771),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1796),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1749),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1805),
.B(n_1755),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1805),
.B(n_1739),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1796),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1791),
.B(n_1739),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1791),
.B(n_1739),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1806),
.A2(n_1692),
.B1(n_1763),
.B2(n_1704),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1781),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1790),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1790),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1800),
.A2(n_1707),
.B1(n_1708),
.B2(n_1714),
.Y(n_1841)
);

OAI31xp33_ASAP7_75t_L g1842 ( 
.A1(n_1797),
.A2(n_1705),
.A3(n_1764),
.B(n_1746),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1793),
.Y(n_1843)
);

AOI33xp33_ASAP7_75t_L g1844 ( 
.A1(n_1789),
.A2(n_1767),
.A3(n_1703),
.B1(n_1758),
.B2(n_1711),
.B3(n_1708),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1801),
.B(n_1640),
.Y(n_1845)
);

INVx4_ASAP7_75t_L g1846 ( 
.A(n_1769),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1789),
.B(n_1751),
.C(n_1730),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1739),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1797),
.B(n_1730),
.C(n_1721),
.Y(n_1849)
);

INVx4_ASAP7_75t_L g1850 ( 
.A(n_1769),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1793),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1784),
.A2(n_1746),
.B1(n_1715),
.B2(n_1710),
.C(n_1717),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1769),
.B(n_1714),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1769),
.B(n_1596),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1780),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1809),
.B(n_1794),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1814),
.B(n_1794),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1814),
.B(n_1788),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1845),
.B(n_1801),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1809),
.B(n_1785),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1821),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1825),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1813),
.B(n_1785),
.Y(n_1865)
);

AND2x4_ASAP7_75t_SL g1866 ( 
.A(n_1828),
.B(n_1769),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1825),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1837),
.B(n_1806),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1808),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1845),
.B(n_1801),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1810),
.B(n_1773),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1827),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1813),
.B(n_1785),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1818),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1816),
.B(n_1798),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1826),
.B(n_1785),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1814),
.B(n_1788),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1853),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1827),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1830),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1810),
.B(n_1773),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1855),
.B(n_1783),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1815),
.B(n_1798),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1826),
.B(n_1785),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1828),
.B(n_1785),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1855),
.B(n_1783),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1854),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1828),
.B(n_1785),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1839),
.B(n_1783),
.Y(n_1890)
);

AND2x4_ASAP7_75t_SL g1891 ( 
.A(n_1853),
.B(n_1769),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1838),
.Y(n_1892)
);

NAND2x1_ASAP7_75t_L g1893 ( 
.A(n_1854),
.B(n_1792),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1830),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1829),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1820),
.B(n_1802),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1834),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1839),
.B(n_1787),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1852),
.B(n_1782),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1831),
.B(n_1782),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1899),
.B(n_1884),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1882),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1862),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1875),
.B(n_1842),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1878),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1882),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1886),
.B(n_1889),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1887),
.Y(n_1908)
);

OAI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1868),
.A2(n_1812),
.B(n_1824),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1887),
.Y(n_1910)
);

INVxp67_ASAP7_75t_SL g1911 ( 
.A(n_1869),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1886),
.B(n_1848),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1889),
.B(n_1848),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1862),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1863),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1863),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1883),
.B(n_1844),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1893),
.A2(n_1784),
.B1(n_1871),
.B2(n_1881),
.Y(n_1918)
);

AND3x2_ASAP7_75t_L g1919 ( 
.A(n_1888),
.B(n_1885),
.C(n_1876),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1871),
.B(n_1840),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1864),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1881),
.B(n_1840),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1878),
.A2(n_1812),
.B1(n_1847),
.B2(n_1841),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1856),
.B(n_1833),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1878),
.A2(n_1721),
.B(n_1822),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1878),
.B(n_1692),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1866),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1856),
.B(n_1833),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1864),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1876),
.B(n_1835),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1892),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1859),
.B(n_1843),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1900),
.B(n_1832),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1857),
.A2(n_1803),
.B1(n_1800),
.B2(n_1823),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1885),
.B(n_1835),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1867),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1867),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1872),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1893),
.A2(n_1777),
.B(n_1792),
.C(n_1779),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1872),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1859),
.B(n_1832),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1866),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1860),
.B(n_1836),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1857),
.B(n_1651),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1890),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1861),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1860),
.B(n_1836),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1901),
.B(n_1896),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1903),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1917),
.B(n_1896),
.Y(n_1950)
);

NOR2x1p5_ASAP7_75t_L g1951 ( 
.A(n_1911),
.B(n_1598),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1903),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1914),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1945),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1914),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1945),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1919),
.Y(n_1958)
);

OR2x6_ASAP7_75t_L g1959 ( 
.A(n_1905),
.B(n_1888),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1915),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1927),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1915),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1945),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1916),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1920),
.B(n_1870),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1916),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1931),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1920),
.B(n_1870),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1921),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1904),
.B(n_1857),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1921),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1907),
.B(n_1858),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1912),
.B(n_1858),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1912),
.B(n_1858),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1923),
.B(n_1909),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1929),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_L g1977 ( 
.A(n_1909),
.B(n_1807),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1922),
.B(n_1890),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1923),
.B(n_1858),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1922),
.B(n_1898),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1913),
.B(n_1877),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1944),
.B(n_1905),
.Y(n_1982)
);

OAI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1918),
.A2(n_1777),
.B(n_1891),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1902),
.B(n_1898),
.Y(n_1984)
);

O2A1O1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1975),
.A2(n_1918),
.B(n_1934),
.C(n_1925),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1958),
.B(n_1926),
.Y(n_1986)
);

NAND3xp33_ASAP7_75t_SL g1987 ( 
.A(n_1983),
.B(n_1939),
.C(n_1819),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1954),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1977),
.A2(n_1942),
.B1(n_1943),
.B2(n_1947),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1977),
.A2(n_1942),
.B1(n_1891),
.B2(n_1877),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1949),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1961),
.A2(n_1877),
.B1(n_1913),
.B2(n_1943),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1973),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1949),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1952),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1973),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1967),
.B(n_1947),
.Y(n_1997)
);

OAI322xp33_ASAP7_75t_L g1998 ( 
.A1(n_1979),
.A2(n_1908),
.A3(n_1906),
.B1(n_1902),
.B2(n_1910),
.C1(n_1932),
.C2(n_1936),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1950),
.B(n_1941),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1982),
.B(n_1930),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1951),
.A2(n_1877),
.B1(n_1935),
.B2(n_1930),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1948),
.B(n_1970),
.Y(n_2002)
);

INVxp67_ASAP7_75t_L g2003 ( 
.A(n_1959),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1957),
.A2(n_1906),
.B(n_1902),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1957),
.B(n_1935),
.Y(n_2005)
);

AOI222xp33_ASAP7_75t_L g2006 ( 
.A1(n_1972),
.A2(n_1924),
.B1(n_1928),
.B2(n_1792),
.C1(n_1779),
.C2(n_1776),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

NOR4xp25_ASAP7_75t_SL g2008 ( 
.A(n_1952),
.B(n_1940),
.C(n_1938),
.D(n_1937),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1972),
.B(n_1906),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1974),
.B(n_1924),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1959),
.Y(n_2011)
);

A2O1A1Ixp33_ASAP7_75t_L g2012 ( 
.A1(n_1974),
.A2(n_1702),
.B(n_1822),
.C(n_1792),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1997),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1988),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1988),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1985),
.A2(n_1959),
.B1(n_1956),
.B2(n_1963),
.C(n_1954),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1991),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1994),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_2011),
.Y(n_2019)
);

OAI33xp33_ASAP7_75t_L g2020 ( 
.A1(n_2003),
.A2(n_1953),
.A3(n_1955),
.B1(n_1964),
.B2(n_1976),
.B3(n_1971),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1987),
.A2(n_1963),
.B(n_1956),
.Y(n_2021)
);

NOR2x1_ASAP7_75t_L g2022 ( 
.A(n_2011),
.B(n_1960),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2007),
.B(n_1986),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_2005),
.B(n_1981),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1999),
.B(n_1978),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2010),
.B(n_1978),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1995),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2007),
.B(n_1981),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1993),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2009),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2009),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_2004),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1986),
.A2(n_1969),
.B1(n_1908),
.B2(n_1910),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2014),
.Y(n_2034)
);

NOR3xp33_ASAP7_75t_L g2035 ( 
.A(n_2016),
.B(n_1998),
.C(n_2000),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_SL g2036 ( 
.A(n_2025),
.B(n_1996),
.Y(n_2036)
);

AOI21xp33_ASAP7_75t_SL g2037 ( 
.A1(n_2032),
.A2(n_2002),
.B(n_1989),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2015),
.Y(n_2038)
);

AOI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_2032),
.A2(n_1989),
.B1(n_1990),
.B2(n_2012),
.C(n_1992),
.Y(n_2039)
);

OAI222xp33_ASAP7_75t_L g2040 ( 
.A1(n_2022),
.A2(n_2001),
.B1(n_2008),
.B2(n_1968),
.C1(n_1965),
.C2(n_1984),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_2023),
.B(n_2012),
.Y(n_2041)
);

OAI21xp33_ASAP7_75t_L g2042 ( 
.A1(n_2028),
.A2(n_2006),
.B(n_1968),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2024),
.B(n_1928),
.Y(n_2043)
);

OAI21xp33_ASAP7_75t_SL g2044 ( 
.A1(n_2021),
.A2(n_1965),
.B(n_1962),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2029),
.Y(n_2045)
);

AOI211xp5_ASAP7_75t_L g2046 ( 
.A1(n_2019),
.A2(n_1960),
.B(n_1966),
.C(n_1962),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2036),
.B(n_2030),
.Y(n_2047)
);

NOR3xp33_ASAP7_75t_L g2048 ( 
.A(n_2037),
.B(n_2013),
.C(n_2031),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_2045),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_2040),
.A2(n_2020),
.B(n_2033),
.Y(n_2050)
);

OAI211xp5_ASAP7_75t_L g2051 ( 
.A1(n_2041),
.A2(n_2035),
.B(n_2039),
.C(n_2044),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_L g2052 ( 
.A1(n_2039),
.A2(n_2029),
.B(n_2027),
.C(n_2017),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2043),
.B(n_2024),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_L g2054 ( 
.A(n_2034),
.B(n_2018),
.C(n_2025),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_2042),
.A2(n_2026),
.B1(n_1966),
.B2(n_1984),
.C(n_1910),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2046),
.A2(n_2026),
.B(n_1908),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_2038),
.B(n_1980),
.C(n_1936),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2043),
.B(n_1980),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2041),
.A2(n_1932),
.B1(n_1865),
.B2(n_1873),
.Y(n_2059)
);

NAND4xp25_ASAP7_75t_L g2060 ( 
.A(n_2051),
.B(n_2050),
.C(n_2048),
.D(n_2053),
.Y(n_2060)
);

NAND3xp33_ASAP7_75t_L g2061 ( 
.A(n_2052),
.B(n_1937),
.C(n_1929),
.Y(n_2061)
);

OAI21xp5_ASAP7_75t_SL g2062 ( 
.A1(n_2047),
.A2(n_1873),
.B(n_1865),
.Y(n_2062)
);

AND4x1_ASAP7_75t_L g2063 ( 
.A(n_2054),
.B(n_1688),
.C(n_1647),
.D(n_1938),
.Y(n_2063)
);

AOI221x1_ASAP7_75t_L g2064 ( 
.A1(n_2056),
.A2(n_1940),
.B1(n_1946),
.B2(n_1879),
.C(n_1897),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_SL g2065 ( 
.A1(n_2049),
.A2(n_1647),
.B1(n_1688),
.B2(n_1697),
.Y(n_2065)
);

OAI211xp5_ASAP7_75t_SL g2066 ( 
.A1(n_2055),
.A2(n_1696),
.B(n_1946),
.C(n_1933),
.Y(n_2066)
);

AOI211xp5_ASAP7_75t_L g2067 ( 
.A1(n_2059),
.A2(n_1696),
.B(n_1811),
.C(n_1779),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2061),
.Y(n_2068)
);

AOI211xp5_ASAP7_75t_SL g2069 ( 
.A1(n_2065),
.A2(n_2058),
.B(n_2057),
.C(n_1740),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2060),
.A2(n_2066),
.B1(n_1850),
.B2(n_1846),
.Y(n_2070)
);

AOI211xp5_ASAP7_75t_L g2071 ( 
.A1(n_2062),
.A2(n_1710),
.B(n_1715),
.C(n_1786),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2067),
.A2(n_1786),
.B(n_1776),
.C(n_1774),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2064),
.Y(n_2073)
);

NAND4xp25_ASAP7_75t_L g2074 ( 
.A(n_2063),
.B(n_1850),
.C(n_1846),
.D(n_1706),
.Y(n_2074)
);

OAI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_2068),
.A2(n_1846),
.B(n_1850),
.C(n_1799),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2074),
.B(n_1697),
.Y(n_2076)
);

NAND4xp75_ASAP7_75t_L g2077 ( 
.A(n_2073),
.B(n_1648),
.C(n_1646),
.D(n_1624),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_2069),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2070),
.B(n_1879),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2071),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2078),
.B(n_2072),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_L g2082 ( 
.A(n_2075),
.B(n_1843),
.C(n_1851),
.Y(n_2082)
);

NAND3x1_ASAP7_75t_L g2083 ( 
.A(n_2076),
.B(n_1897),
.C(n_1894),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2081),
.A2(n_2077),
.B(n_2080),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_2082),
.B1(n_2079),
.B2(n_2083),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2085),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2085),
.Y(n_2087)
);

OA22x2_ASAP7_75t_L g2088 ( 
.A1(n_2086),
.A2(n_1894),
.B1(n_1880),
.B2(n_1851),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2087),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_2089),
.A2(n_1880),
.B(n_1895),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2088),
.A2(n_1656),
.B(n_1616),
.C(n_1834),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_1895),
.B(n_1874),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2092),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2093),
.Y(n_2094)
);

OAI221xp5_ASAP7_75t_R g2095 ( 
.A1(n_2094),
.A2(n_2090),
.B1(n_1712),
.B2(n_1817),
.C(n_1874),
.Y(n_2095)
);

AOI211xp5_ASAP7_75t_L g2096 ( 
.A1(n_2095),
.A2(n_1656),
.B(n_1694),
.C(n_1698),
.Y(n_2096)
);


endmodule