module fake_jpeg_777_n_69 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_19),
.Y(n_31)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_21),
.C(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_24),
.C(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_20),
.B1(n_29),
.B2(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_22),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_28),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_39),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_28),
.C(n_21),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.C(n_38),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_2),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_21),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_22),
.C(n_13),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_49),
.B(n_26),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_59),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_11),
.C(n_10),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_61),
.CI(n_60),
.CON(n_65),
.SN(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_1),
.B(n_4),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_65),
.B(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_6),
.C(n_7),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_7),
.Y(n_69)
);


endmodule