module real_jpeg_451_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_49),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_63),
.B1(n_70),
.B2(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_63),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_63),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_69),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_69),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_70),
.B1(n_73),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_84),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_84),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_84),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_70),
.B1(n_73),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_8),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_131),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_131),
.Y(n_244)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_10),
.A2(n_39),
.B1(n_55),
.B2(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_39),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_13),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_73),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_15),
.B(n_132),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_15),
.A2(n_54),
.B(n_55),
.C(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_15),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_15),
.B(n_60),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_15),
.B(n_27),
.C(n_45),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_15),
.A2(n_40),
.B1(n_42),
.B2(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_15),
.B(n_33),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_15),
.B(n_50),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_20),
.B(n_112),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.C(n_66),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_22),
.A2(n_23),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_24),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_26),
.A2(n_33),
.B1(n_100),
.B2(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_32),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_31),
.A2(n_32),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_31),
.A2(n_32),
.B1(n_159),
.B2(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_31),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_31),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_31),
.A2(n_32),
.B1(n_215),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_32),
.A2(n_174),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_32),
.B(n_188),
.Y(n_217)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_33),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_33),
.A2(n_187),
.B(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_42),
.B1(n_54),
.B2(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_40),
.B(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_42),
.A2(n_61),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_43),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_43),
.B(n_180),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_47),
.A2(n_89),
.B1(n_90),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_47),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_47),
.A2(n_200),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_47),
.A2(n_89),
.B1(n_177),
.B2(n_211),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_50),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_51),
.B(n_66),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_64),
.B1(n_65),
.B2(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_52),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_52),
.A2(n_152),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_60),
.B1(n_151),
.B2(n_168),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_59),
.C(n_60),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_56),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_55),
.A2(n_70),
.A3(n_77),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_56),
.B(n_79),
.Y(n_156)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_60),
.B(n_128),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_62),
.A2(n_64),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_64),
.A2(n_127),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_81),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_75),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_70),
.A2(n_74),
.B(n_184),
.C(n_193),
.Y(n_192)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_76),
.A2(n_105),
.B(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_77),
.Y(n_79)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_82),
.B(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_94),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_89),
.A2(n_179),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_108),
.B2(n_111),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_107),
.B1(n_109),
.B2(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_100),
.A2(n_184),
.B(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_129),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_120),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_121),
.B(n_123),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_161),
.B(n_279),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_137),
.B(n_139),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_140),
.B(n_144),
.Y(n_264)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_146),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_153),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_147),
.B(n_149),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_153),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_157),
.B1(n_158),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI31xp33_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_261),
.A3(n_271),
.B(n_276),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_205),
.B(n_260),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_189),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_164),
.B(n_189),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_175),
.C(n_181),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_165),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_170),
.C(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_175),
.B(n_181),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_185),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_190),
.B(n_202),
.C(n_204),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_255),
.B(n_259),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_224),
.B(n_254),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_214),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_236),
.B(n_253),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_247),
.B(n_252),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_246),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_245),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);


endmodule