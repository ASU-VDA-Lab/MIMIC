module real_jpeg_25856_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_32),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_1),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_1),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_111),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_111),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_111),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_62),
.B1(n_158),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_163),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_163),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_163),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_72),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_8),
.B(n_26),
.C(n_39),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_92),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_44),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_47),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_107)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_13),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_154),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_154),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_154),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_89),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_63),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_14),
.A2(n_26),
.B1(n_33),
.B2(n_89),
.Y(n_177)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_94),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_21),
.A2(n_74),
.B1(n_75),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_21),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_49),
.B2(n_73),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_22),
.A2(n_50),
.B(n_52),
.Y(n_133)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_24),
.A2(n_34),
.B1(n_50),
.B2(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_25),
.A2(n_28),
.B1(n_144),
.B2(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_25),
.A2(n_100),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_25),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_25),
.A2(n_223),
.B1(n_230),
.B2(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_33),
.B1(n_39),
.B2(n_41),
.Y(n_42)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_27),
.Y(n_195)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_102),
.Y(n_146)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_29),
.B(n_31),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_31),
.A2(n_146),
.B(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_33),
.B(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_34),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_45),
.Y(n_34)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_35),
.A2(n_42),
.B1(n_43),
.B2(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_35),
.A2(n_42),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_35),
.A2(n_45),
.B(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_35),
.A2(n_42),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_35),
.A2(n_42),
.B1(n_208),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_35),
.A2(n_77),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_38),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_37),
.B(n_59),
.C(n_85),
.Y(n_249)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_38),
.B(n_204),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_38),
.A2(n_84),
.B(n_248),
.C(n_249),
.Y(n_247)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_42),
.A2(n_79),
.B(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_42),
.B(n_159),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_48),
.A2(n_80),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_66),
.B(n_68),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_109),
.B(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_53),
.A2(n_55),
.B1(n_162),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_69),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_72),
.B1(n_157),
.B2(n_161),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_54),
.A2(n_72),
.B1(n_110),
.B2(n_169),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_55),
.A2(n_118),
.B(n_121),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_65),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_56),
.A2(n_59),
.B(n_160),
.C(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_57),
.B(n_58),
.C(n_70),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_59),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_59),
.B(n_159),
.CON(n_248),
.SN(n_248)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_70),
.B(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_81),
.B(n_93),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_81),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_92),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_92),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_82),
.A2(n_92),
.B1(n_189),
.B2(n_248),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_88),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_83),
.A2(n_125),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_92),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_115),
.B1(n_131),
.B2(n_132),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_94),
.B(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.C(n_108),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_95),
.A2(n_96),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_101),
.A2(n_177),
.B(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_103),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_105),
.B(n_108),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_133),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_130),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_125),
.A2(n_126),
.B(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_309),
.B(n_314),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_298),
.B(n_308),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_196),
.B(n_280),
.C(n_297),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_181),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_139),
.B(n_181),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_164),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_148),
.B2(n_149),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_141),
.B(n_149),
.C(n_164),
.Y(n_281)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_143),
.B(n_147),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_183),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_174),
.B2(n_180),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_167),
.B(n_170),
.C(n_180),
.Y(n_296)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_173),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_182),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_185),
.B(n_186),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_193),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_279),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_274),
.B(n_278),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_260),
.B(n_273),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_244),
.B(n_259),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_218),
.B(n_243),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_217),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_242),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_225),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_236),
.B(n_241),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_258),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_258),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_254),
.C(n_257),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_296),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);


endmodule