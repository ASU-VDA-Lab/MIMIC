module fake_jpeg_23622_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_21),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_23),
.B1(n_29),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_27),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_15),
.B1(n_28),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_15),
.B1(n_20),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_29),
.B1(n_20),
.B2(n_19),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_22),
.B1(n_16),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_67),
.B1(n_55),
.B2(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_61),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_22),
.B1(n_37),
.B2(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_74),
.C(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_79),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_53),
.B1(n_51),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_92),
.B1(n_60),
.B2(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_42),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_63),
.Y(n_99)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_70),
.B1(n_66),
.B2(n_69),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_54),
.B(n_27),
.C(n_35),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_69),
.B(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_106),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_52),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_99),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_109),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_83),
.B(n_94),
.C(n_78),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_107),
.B1(n_78),
.B2(n_85),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_72),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_72),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_53),
.C(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_45),
.C(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_120),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_117),
.B1(n_100),
.B2(n_97),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_98),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_82),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_78),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_98),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_27),
.B(n_18),
.C(n_24),
.D(n_45),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_24),
.C(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_113),
.B1(n_121),
.B2(n_112),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_129),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_117),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_97),
.B1(n_109),
.B2(n_18),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_27),
.B1(n_24),
.B2(n_9),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_24),
.C(n_13),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_143),
.B1(n_147),
.B2(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_144),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_116),
.B1(n_124),
.B2(n_9),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_24),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_145),
.B(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_1),
.B(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_131),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_136),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_153),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_155),
.Y(n_157)
);

AOI31xp67_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_128),
.A3(n_133),
.B(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

FAx1_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_139),
.CI(n_147),
.CON(n_161),
.SN(n_161)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_150),
.B1(n_153),
.B2(n_12),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_164),
.Y(n_169)
);

AOI31xp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_7),
.A3(n_8),
.B(n_157),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_8),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_162),
.B(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);


endmodule