module fake_ariane_869_n_1837 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1837);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1837;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_95),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_116),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_24),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_20),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_94),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_174),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_31),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_80),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_6),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_108),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_61),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_82),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_65),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_58),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_151),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_14),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_70),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_59),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_92),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_90),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_170),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_68),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_19),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_141),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_45),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_119),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_74),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_153),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_17),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_180),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_40),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_87),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_38),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_73),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_76),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_42),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_30),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_166),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_19),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_71),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_88),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_67),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_117),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_35),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_110),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_69),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_85),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_142),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_52),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_33),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_157),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_24),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_79),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_50),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_34),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_15),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_115),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_18),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_30),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_137),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_107),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_36),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_15),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_51),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_34),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_165),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_46),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_9),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_81),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_64),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_132),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_118),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_25),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_12),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_121),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_123),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_101),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_160),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_48),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_124),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_172),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_158),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_148),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_37),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_140),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_2),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_48),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_21),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_138),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_83),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_182),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_113),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_12),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_86),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_155),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_36),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_100),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_126),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_46),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_125),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_14),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_13),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_28),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_11),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_41),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_18),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_33),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_175),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_10),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_185),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_35),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_60),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_104),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_66),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_199),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_199),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_199),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_240),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_199),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_239),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_239),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_235),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_239),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_241),
.B(n_4),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_239),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_225),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_293),
.B(n_6),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_239),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_233),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_247),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_250),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_252),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_219),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_230),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_226),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_306),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_249),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_255),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_259),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_226),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_276),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_233),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_276),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_261),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_304),
.B(n_7),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_262),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_286),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_193),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_190),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_187),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_266),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_191),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_190),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_205),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_205),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_216),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_193),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_272),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_195),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_216),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_280),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_283),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_280),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_269),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_287),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_341),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_201),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_287),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_222),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_284),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_294),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_204),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_297),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_188),
.B(n_8),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_197),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_296),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_233),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_292),
.B(n_8),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_243),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_213),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_298),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_299),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_243),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_254),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_291),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_197),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_282),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_300),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_302),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_301),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_308),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_307),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_319),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_204),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_436),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_189),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_433),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_383),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_372),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_408),
.B(n_316),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_387),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_416),
.B(n_192),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_420),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_373),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_426),
.A2(n_315),
.B1(n_344),
.B2(n_268),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_376),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_391),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_397),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_420),
.B(n_200),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_378),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_439),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_439),
.B(n_206),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_394),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_210),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_212),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_377),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_384),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_431),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_403),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_405),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_444),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_411),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_448),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_413),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_400),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_400),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_396),
.B(n_253),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_408),
.B(n_215),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_221),
.B(n_218),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_408),
.B(n_316),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_421),
.B(n_253),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_418),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_442),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_402),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_422),
.B(n_224),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_453),
.B(n_282),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_422),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_483),
.Y(n_542)
);

INVxp33_ASAP7_75t_SL g543 ( 
.A(n_465),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_478),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_466),
.B(n_198),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_466),
.B(n_390),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_388),
.Y(n_548)
);

INVx4_ASAP7_75t_SL g549 ( 
.A(n_495),
.Y(n_549)
);

AND2x2_ASAP7_75t_SL g550 ( 
.A(n_540),
.B(n_446),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_480),
.B(n_425),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_472),
.B(n_198),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_480),
.B(n_429),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_471),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_471),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_480),
.A2(n_451),
.B1(n_440),
.B2(n_461),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_471),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_536),
.Y(n_561)
);

NOR2x1p5_ASAP7_75t_L g562 ( 
.A(n_489),
.B(n_437),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_478),
.B(n_409),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_476),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_484),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_478),
.B(n_438),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_502),
.B(n_456),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_472),
.B(n_530),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_480),
.B(n_512),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_517),
.B(n_459),
.C(n_452),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_502),
.B(n_398),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_520),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_472),
.B(n_423),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_538),
.A2(n_434),
.B1(n_454),
.B2(n_458),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

BUFx8_ASAP7_75t_SL g586 ( 
.A(n_513),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_472),
.B(n_198),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_528),
.B(n_468),
.Y(n_589)
);

AND3x2_ASAP7_75t_L g590 ( 
.A(n_540),
.B(n_359),
.C(n_265),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_530),
.B(n_410),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_480),
.B(n_229),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_516),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_528),
.B(n_423),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_504),
.Y(n_596)
);

OR2x2_ASAP7_75t_SL g597 ( 
.A(n_469),
.B(n_463),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_509),
.B(n_417),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

NOR2x1p5_ASAP7_75t_L g600 ( 
.A(n_470),
.B(n_203),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_487),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_509),
.B(n_419),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_504),
.B(n_457),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_481),
.A2(n_273),
.B1(n_360),
.B2(n_349),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_512),
.A2(n_310),
.B1(n_353),
.B2(n_356),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_530),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_510),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_487),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_530),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_510),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_512),
.B(n_234),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_512),
.B(n_236),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_468),
.B(n_427),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_511),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_496),
.B(n_450),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_512),
.B(n_237),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_511),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_477),
.B(n_427),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_541),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_495),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_481),
.A2(n_327),
.B1(n_366),
.B2(n_333),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_492),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_500),
.B(n_525),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_521),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_SL g635 ( 
.A(n_500),
.B(n_203),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_L g636 ( 
.A1(n_525),
.A2(n_220),
.B1(n_279),
.B2(n_311),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_492),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_524),
.B(n_198),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

AND3x2_ASAP7_75t_L g641 ( 
.A(n_533),
.B(n_455),
.C(n_450),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_477),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

OAI22xp33_ASAP7_75t_L g645 ( 
.A1(n_533),
.A2(n_327),
.B1(n_333),
.B2(n_366),
.Y(n_645)
);

NOR2x1p5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_220),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_529),
.B(n_245),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_485),
.B(n_455),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_534),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_508),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_474),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_529),
.A2(n_430),
.B1(n_428),
.B2(n_432),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_539),
.B(n_320),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_537),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_531),
.B(n_428),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_474),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_495),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_531),
.B(n_430),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_482),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_539),
.B(n_251),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_508),
.B(n_256),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_474),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_485),
.B(n_493),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_493),
.B(n_432),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_508),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_515),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_498),
.B(n_460),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_498),
.B(n_435),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_499),
.B(n_435),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_495),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_491),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_499),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_491),
.A2(n_363),
.B1(n_364),
.B2(n_361),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_495),
.B(n_326),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_491),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_535),
.A2(n_443),
.B1(n_445),
.B2(n_447),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_491),
.B(n_443),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_467),
.A2(n_445),
.B1(n_447),
.B2(n_449),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_508),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_518),
.B(n_449),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_467),
.A2(n_362),
.B1(n_338),
.B2(n_352),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_518),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_467),
.B(n_198),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_586),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_604),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_547),
.B(n_519),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_632),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_589),
.B(n_523),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_632),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_604),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_607),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_593),
.Y(n_696)
);

BUFx8_ASAP7_75t_L g697 ( 
.A(n_668),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_589),
.B(n_523),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_550),
.B(n_196),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_548),
.B(n_523),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_548),
.B(n_674),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_655),
.A2(n_535),
.B1(n_475),
.B2(n_522),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_559),
.B(n_202),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_621),
.B(n_523),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_607),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_570),
.B(n_460),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_551),
.B(n_358),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_577),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_551),
.B(n_279),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_642),
.B(n_508),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_636),
.B(n_314),
.C(n_311),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_621),
.B(n_202),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_SL g713 ( 
.A(n_573),
.B(n_581),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_610),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_545),
.B(n_347),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_624),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_554),
.B(n_314),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_545),
.B(n_207),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_624),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_665),
.B(n_207),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_574),
.B(n_209),
.Y(n_721)
);

BUFx5_ASAP7_75t_L g722 ( 
.A(n_634),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_648),
.B(n_209),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_655),
.A2(n_630),
.B1(n_676),
.B2(n_685),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_554),
.B(n_211),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_594),
.B(n_211),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_626),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_609),
.B(n_214),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_630),
.A2(n_535),
.B1(n_522),
.B2(n_507),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_594),
.B(n_618),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_609),
.B(n_214),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_618),
.B(n_217),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_625),
.B(n_217),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_592),
.A2(n_616),
.B1(n_622),
.B2(n_617),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_625),
.B(n_223),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_582),
.B(n_223),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_564),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_684),
.A2(n_522),
.B(n_507),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_670),
.B(n_267),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_598),
.B(n_462),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_596),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_555),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_582),
.B(n_267),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_576),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_598),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_566),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_670),
.B(n_278),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_312),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_684),
.Y(n_749)
);

INVx8_ASAP7_75t_L g750 ( 
.A(n_602),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_555),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_557),
.Y(n_752)
);

BUFx8_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_679),
.A2(n_368),
.B(n_370),
.C(n_271),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_592),
.B(n_317),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_616),
.B(n_322),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_313),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_617),
.B(n_322),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_313),
.Y(n_759)
);

BUFx5_ASAP7_75t_L g760 ( 
.A(n_634),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_569),
.B(n_321),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_608),
.B(n_321),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_565),
.B(n_462),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_557),
.B(n_227),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_573),
.B(n_323),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_569),
.B(n_323),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_L g767 ( 
.A1(n_647),
.A2(n_507),
.B(n_506),
.C(n_503),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_622),
.B(n_324),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_676),
.A2(n_571),
.B1(n_591),
.B2(n_568),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_558),
.B(n_342),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_578),
.B(n_341),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_543),
.B(n_542),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_542),
.B(n_324),
.Y(n_773)
);

AO22x1_ASAP7_75t_L g774 ( 
.A1(n_661),
.A2(n_342),
.B1(n_349),
.B2(n_343),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_341),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_602),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_585),
.A2(n_343),
.B1(n_334),
.B2(n_340),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_562),
.B(n_404),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_SL g780 ( 
.A(n_600),
.B(n_331),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_595),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_591),
.B(n_331),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_561),
.B(n_334),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_658),
.A2(n_506),
.B(n_503),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_599),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_560),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_563),
.B(n_340),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_666),
.B(n_345),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_560),
.B(n_345),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_671),
.B(n_346),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_675),
.B(n_346),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_603),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_685),
.A2(n_506),
.B1(n_475),
.B2(n_503),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_662),
.B(n_350),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_635),
.B(n_350),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_662),
.A2(n_475),
.B1(n_486),
.B2(n_282),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_584),
.B(n_367),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_579),
.A2(n_414),
.B1(n_337),
.B2(n_369),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_585),
.A2(n_486),
.B(n_257),
.C(n_330),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_553),
.A2(n_588),
.B1(n_663),
.B2(n_651),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_679),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_584),
.B(n_367),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_651),
.B(n_369),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_605),
.B(n_414),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_611),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_636),
.A2(n_337),
.B1(n_295),
.B2(n_339),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_645),
.B(n_228),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_SL g808 ( 
.A1(n_606),
.A2(n_289),
.B1(n_270),
.B2(n_275),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_664),
.A2(n_673),
.B(n_686),
.C(n_677),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_572),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_615),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_641),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_680),
.B(n_486),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_572),
.A2(n_318),
.B(n_336),
.C(n_348),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_680),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_546),
.B(n_231),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_575),
.A2(n_281),
.B(n_332),
.C(n_328),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_552),
.B(n_556),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_619),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_647),
.A2(n_277),
.B(n_335),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_623),
.A2(n_285),
.B1(n_232),
.B2(n_238),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_633),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_575),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_597),
.B(n_242),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_639),
.A2(n_505),
.B1(n_497),
.B2(n_495),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_SL g826 ( 
.A1(n_590),
.A2(n_288),
.B1(n_244),
.B2(n_246),
.Y(n_826)
);

BUFx6f_ASAP7_75t_SL g827 ( 
.A(n_553),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_546),
.B(n_248),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_590),
.B(n_258),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_583),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_645),
.B(n_309),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_629),
.B(n_305),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_583),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_546),
.B(n_351),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_643),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_641),
.B(n_497),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_629),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_646),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_553),
.A2(n_303),
.B1(n_260),
.B2(n_263),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_587),
.A2(n_505),
.B(n_497),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_657),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_544),
.B(n_10),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_784),
.A2(n_663),
.B(n_644),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_801),
.A2(n_628),
.B(n_587),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_730),
.B(n_601),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_694),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_750),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_692),
.A2(n_631),
.B(n_640),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_750),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_744),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_698),
.A2(n_631),
.B(n_640),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_688),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_724),
.A2(n_553),
.B1(n_588),
.B2(n_653),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_708),
.B(n_678),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_701),
.B(n_612),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_767),
.A2(n_613),
.B(n_627),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_767),
.A2(n_627),
.B(n_612),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_700),
.B(n_613),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_649),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_809),
.A2(n_650),
.B(n_637),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_820),
.A2(n_656),
.B(n_654),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_710),
.A2(n_637),
.B(n_682),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_715),
.A2(n_682),
.B1(n_667),
.B2(n_650),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_813),
.A2(n_667),
.B(n_683),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_738),
.A2(n_629),
.B(n_659),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_742),
.A2(n_672),
.B(n_659),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_740),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_818),
.A2(n_652),
.B(n_553),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_709),
.B(n_652),
.C(n_660),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_751),
.A2(n_659),
.B(n_672),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_752),
.A2(n_659),
.B(n_672),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_718),
.A2(n_672),
.B1(n_678),
.B2(n_681),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_786),
.A2(n_290),
.B(n_357),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_741),
.B(n_549),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_749),
.B(n_546),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_724),
.B(n_546),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_810),
.A2(n_830),
.B(n_823),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_734),
.A2(n_681),
.B1(n_505),
.B2(n_497),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_769),
.B(n_588),
.Y(n_879)
);

AO21x1_ASAP7_75t_L g880 ( 
.A1(n_709),
.A2(n_549),
.B(n_588),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_833),
.A2(n_264),
.B(n_274),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_818),
.A2(n_588),
.B(n_638),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_781),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_691),
.B(n_549),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_749),
.A2(n_354),
.B(n_355),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_761),
.A2(n_365),
.B(n_227),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_726),
.A2(n_495),
.B1(n_497),
.B2(n_505),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_785),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_766),
.A2(n_227),
.B(n_505),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_740),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_792),
.B(n_505),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_750),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_765),
.A2(n_227),
.B(n_505),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_840),
.A2(n_638),
.B(n_687),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_SL g895 ( 
.A1(n_725),
.A2(n_11),
.B(n_13),
.C(n_17),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_695),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_705),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_717),
.A2(n_638),
.B1(n_687),
.B2(n_497),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_806),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_716),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_805),
.B(n_638),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_806),
.A2(n_22),
.B(n_23),
.C(n_27),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_803),
.A2(n_227),
.B(n_638),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_811),
.B(n_819),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_720),
.A2(n_687),
.B(n_98),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_800),
.A2(n_687),
.B(n_106),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_717),
.A2(n_687),
.B1(n_28),
.B2(n_32),
.Y(n_907)
);

AND2x2_ASAP7_75t_SL g908 ( 
.A(n_711),
.B(n_776),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_822),
.B(n_835),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_712),
.A2(n_96),
.B(n_178),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_815),
.B(n_27),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_756),
.A2(n_32),
.B(n_38),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_696),
.B(n_44),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_689),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_757),
.A2(n_127),
.B(n_173),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_815),
.B(n_45),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_707),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_693),
.B(n_49),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_753),
.B(n_51),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_732),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_733),
.B(n_53),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_756),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_714),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_711),
.A2(n_56),
.B(n_63),
.C(n_75),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_740),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_758),
.A2(n_112),
.B(n_120),
.C(n_128),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_737),
.B(n_183),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_735),
.B(n_129),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_759),
.A2(n_131),
.B(n_136),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_746),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_739),
.B(n_747),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_758),
.A2(n_145),
.B1(n_150),
.B2(n_154),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_719),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_779),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_842),
.A2(n_159),
.B(n_161),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_736),
.A2(n_743),
.B(n_790),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_707),
.B(n_167),
.C(n_169),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_737),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_788),
.A2(n_789),
.B(n_728),
.Y(n_939)
);

NOR2x1p5_ASAP7_75t_SL g940 ( 
.A(n_722),
.B(n_760),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_731),
.A2(n_723),
.B(n_832),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_704),
.A2(n_702),
.B(n_825),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_775),
.B(n_727),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_827),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_779),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_706),
.B(n_804),
.Y(n_946)
);

AO22x1_ASAP7_75t_L g947 ( 
.A1(n_753),
.A2(n_697),
.B1(n_776),
.B2(n_745),
.Y(n_947)
);

INVx8_ASAP7_75t_L g948 ( 
.A(n_827),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_779),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_771),
.B(n_763),
.Y(n_950)
);

BUFx8_ASAP7_75t_L g951 ( 
.A(n_690),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_755),
.A2(n_704),
.B1(n_787),
.B2(n_699),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_787),
.B(n_841),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_713),
.A2(n_828),
.B(n_834),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_779),
.A2(n_837),
.B(n_768),
.Y(n_955)
);

AOI22x1_ASAP7_75t_L g956 ( 
.A1(n_837),
.A2(n_778),
.B1(n_799),
.B2(n_838),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_697),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_722),
.B(n_760),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_842),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_837),
.A2(n_783),
.B(n_782),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_722),
.B(n_760),
.Y(n_961)
);

AO22x1_ASAP7_75t_L g962 ( 
.A1(n_812),
.A2(n_829),
.B1(n_824),
.B2(n_797),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_837),
.A2(n_783),
.B(n_794),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_722),
.B(n_760),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_807),
.A2(n_831),
.B(n_754),
.C(n_703),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_762),
.A2(n_798),
.B(n_791),
.C(n_770),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_721),
.A2(n_773),
.B(n_795),
.C(n_814),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_836),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_772),
.B(n_802),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_722),
.B(n_760),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_816),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_770),
.A2(n_748),
.B(n_821),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_780),
.A2(n_796),
.B(n_817),
.C(n_702),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_825),
.A2(n_722),
.B(n_760),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_777),
.B(n_826),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_796),
.A2(n_808),
.B(n_839),
.C(n_729),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_808),
.A2(n_729),
.B(n_793),
.C(n_798),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_793),
.B(n_774),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_764),
.A2(n_801),
.B(n_730),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_764),
.A2(n_730),
.B1(n_801),
.B2(n_715),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_764),
.A2(n_801),
.B(n_730),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_764),
.A2(n_801),
.B(n_730),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_764),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_779),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_696),
.B(n_593),
.C(n_580),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_730),
.B(n_801),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_734),
.A2(n_548),
.B(n_758),
.C(n_756),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_763),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_701),
.A2(n_806),
.B(n_715),
.C(n_548),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_694),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_779),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_708),
.B(n_466),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_694),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_784),
.A2(n_647),
.B(n_820),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_801),
.A2(n_730),
.B(n_698),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_694),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_730),
.B(n_801),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_730),
.B(n_801),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_724),
.A2(n_550),
.B1(n_717),
.B2(n_709),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_688),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_708),
.B(n_466),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_767),
.A2(n_809),
.B(n_730),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_724),
.A2(n_550),
.B1(n_717),
.B2(n_709),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_730),
.B(n_801),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_730),
.B(n_801),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_744),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_744),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_779),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_801),
.A2(n_730),
.B(n_698),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_801),
.A2(n_730),
.B(n_698),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_779),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_767),
.A2(n_809),
.B(n_730),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_701),
.A2(n_806),
.B(n_715),
.C(n_548),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_1011),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_856),
.A2(n_974),
.B(n_961),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_946),
.B(n_986),
.Y(n_1017)
);

INVx6_ASAP7_75t_L g1018 ( 
.A(n_847),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_997),
.B(n_998),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_999),
.A2(n_1003),
.B1(n_978),
.B2(n_854),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_975),
.A2(n_987),
.B1(n_1013),
.B2(n_989),
.C(n_977),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_951),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_948),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_992),
.B(n_1001),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_954),
.A2(n_980),
.B(n_963),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_938),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_958),
.A2(n_964),
.B(n_961),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_SL g1030 ( 
.A1(n_931),
.A2(n_921),
.B(n_916),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_950),
.B(n_988),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_952),
.B(n_995),
.Y(n_1032)
);

BUFx8_ASAP7_75t_SL g1033 ( 
.A(n_1000),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_931),
.B(n_859),
.Y(n_1034)
);

NAND3x1_ASAP7_75t_L g1035 ( 
.A(n_917),
.B(n_913),
.C(n_907),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_979),
.A2(n_982),
.B(n_981),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_970),
.A2(n_994),
.B(n_1002),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_970),
.A2(n_1012),
.B(n_857),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_930),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_953),
.B(n_904),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_928),
.A2(n_866),
.B(n_955),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_884),
.Y(n_1043)
);

AND2x2_ASAP7_75t_SL g1044 ( 
.A(n_876),
.B(n_908),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_866),
.A2(n_865),
.B(n_851),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_928),
.A2(n_865),
.B(n_843),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_953),
.B(n_904),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_914),
.Y(n_1048)
);

OA21x2_ASAP7_75t_L g1049 ( 
.A1(n_860),
.A2(n_935),
.B(n_905),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_844),
.A2(n_921),
.B(n_845),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_959),
.A2(n_889),
.B(n_960),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_845),
.A2(n_858),
.B(n_848),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_869),
.A2(n_855),
.B(n_972),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_909),
.B(n_943),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_925),
.B(n_985),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_880),
.A2(n_886),
.B(n_939),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_936),
.A2(n_893),
.B(n_962),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_862),
.A2(n_942),
.B(n_870),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_966),
.A2(n_906),
.B(n_932),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_867),
.B(n_890),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_943),
.B(n_909),
.Y(n_1061)
);

BUFx10_ASAP7_75t_L g1062 ( 
.A(n_927),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_L g1063 ( 
.A(n_875),
.B(n_991),
.Y(n_1063)
);

AO21x2_ASAP7_75t_L g1064 ( 
.A1(n_876),
.A2(n_868),
.B(n_858),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_847),
.B(n_849),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_887),
.A2(n_916),
.B(n_911),
.Y(n_1066)
);

BUFx12f_ASAP7_75t_L g1067 ( 
.A(n_957),
.Y(n_1067)
);

BUFx4_ASAP7_75t_R g1068 ( 
.A(n_852),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_911),
.A2(n_941),
.B(n_903),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_855),
.A2(n_864),
.B(n_863),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_849),
.B(n_892),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_847),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_883),
.B(n_888),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_871),
.A2(n_877),
.B(n_894),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_872),
.A2(n_891),
.B(n_901),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_891),
.A2(n_967),
.B(n_882),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_915),
.A2(n_929),
.B(n_910),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1080)
);

AND2x2_ASAP7_75t_SL g1081 ( 
.A(n_937),
.B(n_853),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_879),
.A2(n_901),
.B(n_874),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_965),
.A2(n_945),
.B(n_949),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_976),
.A2(n_973),
.B(n_879),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_968),
.B(n_969),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_926),
.A2(n_878),
.B(n_983),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1011),
.B(n_944),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_934),
.A2(n_984),
.B(n_1008),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_912),
.A2(n_899),
.B(n_902),
.C(n_924),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_969),
.B(n_846),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_944),
.B(n_884),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_948),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_896),
.B(n_993),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_922),
.A2(n_920),
.B(n_940),
.C(n_918),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_934),
.A2(n_1008),
.B(n_984),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_897),
.B(n_933),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_983),
.A2(n_956),
.B(n_971),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_SL g1098 ( 
.A1(n_900),
.A2(n_996),
.B(n_990),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_SL g1099 ( 
.A1(n_895),
.A2(n_885),
.B(n_1011),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1011),
.B(n_991),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_873),
.A2(n_881),
.B(n_875),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_SL g1102 ( 
.A1(n_991),
.A2(n_987),
.B1(n_989),
.B2(n_1013),
.C(n_806),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_875),
.A2(n_898),
.B(n_919),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_875),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_875),
.A2(n_987),
.B(n_981),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_987),
.A2(n_999),
.B(n_1003),
.C(n_989),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_946),
.B(n_701),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_957),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_861),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_905),
.A2(n_876),
.B(n_954),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_999),
.B(n_1003),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_987),
.A2(n_981),
.B(n_979),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_876),
.A2(n_977),
.A3(n_980),
.B(n_976),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_876),
.A2(n_977),
.A3(n_980),
.B(n_976),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_856),
.A2(n_974),
.B(n_961),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_849),
.B(n_892),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_946),
.B(n_701),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_SL g1126 ( 
.A1(n_931),
.A2(n_921),
.B(n_986),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_981),
.B(n_979),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_861),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_861),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_987),
.A2(n_1003),
.B1(n_999),
.B2(n_997),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_987),
.A2(n_1003),
.B1(n_999),
.B2(n_997),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_987),
.A2(n_999),
.B(n_1003),
.C(n_989),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_884),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_954),
.A2(n_974),
.B(n_980),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_946),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_987),
.A2(n_981),
.B(n_979),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_946),
.B(n_701),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_946),
.B(n_701),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1141)
);

INVx3_ASAP7_75t_SL g1142 ( 
.A(n_847),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_987),
.A2(n_981),
.B(n_979),
.Y(n_1143)
);

NAND2x1p5_ASAP7_75t_L g1144 ( 
.A(n_1011),
.B(n_849),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_884),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_987),
.A2(n_999),
.B(n_1003),
.C(n_989),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_992),
.B(n_1001),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_987),
.A2(n_1003),
.B1(n_999),
.B2(n_997),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_856),
.A2(n_974),
.B(n_961),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_852),
.B(n_688),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_954),
.A2(n_974),
.B(n_980),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_974),
.A2(n_856),
.B(n_958),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_850),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1011),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_986),
.A2(n_998),
.B(n_997),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_SL g1159 ( 
.A1(n_977),
.A2(n_961),
.B(n_958),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_987),
.A2(n_981),
.B(n_979),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_948),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1032),
.A2(n_1112),
.B(n_1014),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_1015),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1062),
.B(n_1034),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1033),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1061),
.B(n_1017),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1032),
.A2(n_1117),
.B(n_1113),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1061),
.B(n_1107),
.Y(n_1168)
);

INVx3_ASAP7_75t_SL g1169 ( 
.A(n_1073),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_1018),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1033),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1074),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1062),
.B(n_1019),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1022),
.B(n_1133),
.C(n_1106),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1106),
.A2(n_1146),
.B(n_1133),
.C(n_1155),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1021),
.A2(n_1023),
.B(n_1124),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_SL g1177 ( 
.A1(n_1041),
.A2(n_1116),
.B(n_1138),
.C(n_1160),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1026),
.B(n_1147),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1028),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1150),
.A2(n_1158),
.B(n_1152),
.Y(n_1181)
);

CKINVDCx6p67_ASAP7_75t_R g1182 ( 
.A(n_1142),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1031),
.B(n_1136),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1142),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1125),
.B(n_1139),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1146),
.A2(n_1131),
.B1(n_1132),
.B2(n_1148),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1136),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1089),
.A2(n_1094),
.B(n_1140),
.C(n_1054),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1091),
.B(n_1079),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1020),
.B(n_1116),
.Y(n_1190)
);

AND2x2_ASAP7_75t_SL g1191 ( 
.A(n_1020),
.B(n_1044),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1035),
.A2(n_1089),
.B1(n_1081),
.B2(n_1080),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1025),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1055),
.B(n_1060),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1015),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1052),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1161),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1015),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1015),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1159),
.A2(n_1070),
.B(n_1050),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1067),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1156),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1048),
.B(n_1072),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1161),
.B(n_1100),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1102),
.B(n_1119),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1048),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1035),
.A2(n_1084),
.B1(n_1094),
.B2(n_1103),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1068),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1053),
.A2(n_1105),
.B1(n_1077),
.B2(n_1085),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1091),
.B(n_1024),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1073),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1096),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1076),
.A2(n_1127),
.B1(n_1118),
.B2(n_1143),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

CKINVDCx6p67_ASAP7_75t_R g1215 ( 
.A(n_1108),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1068),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1043),
.B(n_1134),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1043),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1134),
.B(n_1145),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1038),
.A2(n_1037),
.B(n_1086),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1093),
.A2(n_1062),
.B1(n_1090),
.B2(n_1064),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1157),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1091),
.B(n_1092),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1065),
.A2(n_1087),
.B(n_1144),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1145),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1119),
.B(n_1120),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1071),
.B(n_1122),
.Y(n_1227)
);

NOR2x1_ASAP7_75t_L g1228 ( 
.A(n_1151),
.B(n_1122),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_1029),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1064),
.A2(n_1122),
.B1(n_1100),
.B2(n_1104),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1051),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1157),
.Y(n_1232)
);

AO32x1_ASAP7_75t_L g1233 ( 
.A1(n_1114),
.A2(n_1129),
.A3(n_1128),
.B1(n_1126),
.B2(n_1030),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_L g1234 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1087),
.B(n_1120),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1104),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1119),
.B(n_1120),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1083),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1119),
.B(n_1120),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1045),
.A2(n_1086),
.B(n_1154),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1101),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1082),
.B(n_1057),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1115),
.A2(n_1129),
.B1(n_1128),
.B2(n_1097),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1110),
.B(n_1141),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1058),
.B(n_1075),
.Y(n_1245)
);

NOR2x1_ASAP7_75t_L g1246 ( 
.A(n_1099),
.B(n_1056),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1069),
.B(n_1042),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1027),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1066),
.B(n_1046),
.Y(n_1249)
);

INVx3_ASAP7_75t_SL g1250 ( 
.A(n_1135),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_1153),
.Y(n_1251)
);

BUFx5_ASAP7_75t_L g1252 ( 
.A(n_1109),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1110),
.A2(n_1130),
.B1(n_1111),
.B2(n_1141),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1016),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1111),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1121),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1123),
.B(n_1130),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_1123),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1137),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1137),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1154),
.B(n_543),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1034),
.B(n_946),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1034),
.B(n_946),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1015),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1074),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1142),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1015),
.Y(n_1267)
);

O2A1O1Ixp5_ASAP7_75t_L g1268 ( 
.A1(n_1059),
.A2(n_1032),
.B(n_1133),
.C(n_1106),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1074),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1089),
.A2(n_912),
.B1(n_1084),
.B2(n_1133),
.C(n_1106),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1022),
.A2(n_1003),
.B(n_999),
.C(n_987),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1034),
.B(n_946),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1032),
.A2(n_997),
.B(n_986),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1074),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_SL g1275 ( 
.A(n_1073),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1022),
.A2(n_1003),
.B(n_999),
.C(n_987),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1074),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1074),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1074),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1039),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1025),
.B(n_849),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1034),
.B(n_946),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1028),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1032),
.A2(n_997),
.B(n_986),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1074),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1028),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1032),
.A2(n_997),
.B(n_986),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1028),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1032),
.A2(n_997),
.B(n_986),
.Y(n_1289)
);

O2A1O1Ixp5_ASAP7_75t_SL g1290 ( 
.A1(n_1041),
.A2(n_1032),
.B(n_647),
.C(n_1116),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1222),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1174),
.A2(n_1186),
.B1(n_1192),
.B2(n_1271),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1165),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1191),
.A2(n_1207),
.B1(n_1192),
.B2(n_1190),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1216),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1230),
.B(n_1235),
.Y(n_1296)
);

AOI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1196),
.A2(n_1167),
.B(n_1162),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1184),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1260),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1207),
.A2(n_1190),
.B1(n_1186),
.B2(n_1174),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_SL g1301 ( 
.A1(n_1188),
.A2(n_1213),
.B(n_1273),
.Y(n_1301)
);

CKINVDCx6p67_ASAP7_75t_R g1302 ( 
.A(n_1215),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1241),
.Y(n_1303)
);

AO21x1_ASAP7_75t_L g1304 ( 
.A1(n_1213),
.A2(n_1200),
.B(n_1205),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1237),
.B(n_1239),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1284),
.A2(n_1289),
.B(n_1287),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1205),
.B(n_1172),
.Y(n_1307)
);

AO21x1_ASAP7_75t_SL g1308 ( 
.A1(n_1220),
.A2(n_1226),
.B(n_1231),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1276),
.A2(n_1175),
.B1(n_1166),
.B2(n_1168),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1265),
.B(n_1269),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1226),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1274),
.B(n_1277),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1216),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1181),
.A2(n_1244),
.B(n_1229),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1243),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1249),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1206),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1250),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1259),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1185),
.B(n_1262),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1233),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1180),
.A2(n_1272),
.B1(n_1263),
.B2(n_1282),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1285),
.B(n_1183),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1180),
.B(n_1178),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1203),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1179),
.B(n_1283),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_1173),
.B1(n_1238),
.B2(n_1182),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1220),
.A2(n_1268),
.B(n_1247),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1194),
.A2(n_1212),
.B1(n_1286),
.B2(n_1221),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1171),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1179),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1233),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1233),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1177),
.A2(n_1290),
.B(n_1253),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1266),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1253),
.A2(n_1246),
.B(n_1255),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1275),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1202),
.B(n_1261),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1247),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1230),
.B(n_1227),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1209),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1189),
.B(n_1288),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1255),
.A2(n_1234),
.B(n_1242),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1283),
.B(n_1288),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1176),
.B(n_1225),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1208),
.A2(n_1169),
.B1(n_1280),
.B2(n_1266),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1248),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1163),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1236),
.B(n_1218),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1251),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1257),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1214),
.A2(n_1270),
.B(n_1199),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1251),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1210),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_SL g1358 ( 
.A1(n_1224),
.A2(n_1197),
.B(n_1193),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1218),
.B(n_1267),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1266),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1257),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1245),
.A2(n_1258),
.B(n_1219),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1210),
.A2(n_1228),
.B1(n_1223),
.B2(n_1201),
.Y(n_1363)
);

BUFx2_ASAP7_75t_R g1364 ( 
.A(n_1211),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1245),
.A2(n_1217),
.B(n_1204),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1254),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1256),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1232),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1252),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1252),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1252),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1195),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1195),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1199),
.A2(n_1264),
.B(n_1267),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1264),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1198),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1281),
.A2(n_1200),
.B(n_1240),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1170),
.B(n_1237),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1170),
.B(n_543),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1187),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1168),
.B(n_543),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1165),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1192),
.A2(n_975),
.B1(n_1003),
.B2(n_999),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1200),
.A2(n_1240),
.B(n_1027),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1216),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1186),
.A2(n_1174),
.B(n_1022),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1260),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1191),
.A2(n_1003),
.B1(n_999),
.B2(n_1116),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1237),
.B(n_1239),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1181),
.A2(n_1243),
.B(n_1036),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1165),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1196),
.A2(n_1041),
.B(n_1162),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1200),
.A2(n_1240),
.B(n_1027),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1187),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1189),
.Y(n_1396)
);

BUFx2_ASAP7_75t_R g1397 ( 
.A(n_1208),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1222),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1186),
.A2(n_987),
.B(n_999),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1303),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1321),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1305),
.B(n_1390),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1354),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1354),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1303),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1324),
.B(n_1322),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1387),
.A2(n_1292),
.B(n_1399),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1315),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1336),
.A2(n_1306),
.B(n_1384),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1381),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1302),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1309),
.A2(n_1329),
.B(n_1295),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1395),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1333),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1305),
.B(n_1390),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1300),
.A2(n_1294),
.B(n_1389),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1396),
.B(n_1348),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1341),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1318),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1328),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1301),
.A2(n_1334),
.B(n_1323),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1320),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1293),
.Y(n_1423)
);

AO21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1340),
.A2(n_1344),
.B(n_1361),
.Y(n_1424)
);

BUFx4f_ASAP7_75t_SL g1425 ( 
.A(n_1302),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1319),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1299),
.B(n_1388),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1296),
.B(n_1343),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1293),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1311),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1307),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1311),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1345),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1358),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1362),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1307),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1393),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1299),
.A2(n_1331),
.B1(n_1343),
.B2(n_1327),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1345),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1361),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1304),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1382),
.A2(n_1355),
.B(n_1340),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1326),
.B(n_1325),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1394),
.A2(n_1393),
.B(n_1297),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1339),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1347),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1325),
.B(n_1344),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1359),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1342),
.B(n_1379),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1362),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1348),
.Y(n_1451)
);

INVx5_ASAP7_75t_L g1452 ( 
.A(n_1396),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1355),
.A2(n_1380),
.B(n_1353),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1338),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1297),
.A2(n_1316),
.B(n_1378),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1353),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1457)
);

AOI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1356),
.A2(n_1334),
.B(n_1323),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1332),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1314),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1352),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_1308),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1356),
.B(n_1373),
.C(n_1377),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1313),
.B(n_1327),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1391),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1350),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1308),
.B(n_1313),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1373),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1330),
.B(n_1296),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1366),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1366),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1335),
.A2(n_1338),
.B(n_1346),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1367),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1335),
.A2(n_1367),
.B(n_1346),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1378),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1407),
.A2(n_1314),
.B1(n_1386),
.B2(n_1295),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1402),
.B(n_1330),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1424),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1431),
.B(n_1330),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1401),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1402),
.B(n_1369),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1401),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1415),
.B(n_1372),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1415),
.B(n_1372),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1434),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1462),
.B(n_1371),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1422),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1406),
.B(n_1350),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1365),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1436),
.B(n_1370),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1436),
.B(n_1374),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1458),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1422),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1470),
.B(n_1376),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1470),
.B(n_1376),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1434),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1375),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1463),
.B(n_1291),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1472),
.B(n_1424),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1375),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1421),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1434),
.B(n_1291),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1419),
.B(n_1398),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1464),
.B(n_1357),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1430),
.B(n_1291),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1416),
.A2(n_1314),
.B1(n_1386),
.B2(n_1351),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1412),
.A2(n_1386),
.B1(n_1364),
.B2(n_1363),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1421),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1448),
.B(n_1349),
.Y(n_1513)
);

INVx8_ASAP7_75t_L g1514 ( 
.A(n_1452),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1421),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1441),
.B(n_1368),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1477),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1477),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1414),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1481),
.A2(n_1442),
.B(n_1453),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1505),
.A2(n_1416),
.B1(n_1512),
.B2(n_1515),
.C(n_1517),
.Y(n_1521)
);

AOI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1505),
.A2(n_1420),
.B1(n_1476),
.B2(n_1474),
.C(n_1473),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1511),
.A2(n_1412),
.B1(n_1427),
.B2(n_1386),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1491),
.B(n_1408),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1495),
.A2(n_1455),
.B(n_1444),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1480),
.B(n_1403),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1511),
.B(n_1465),
.C(n_1456),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1481),
.B(n_1456),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1410),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1413),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1487),
.B(n_1418),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1510),
.B(n_1404),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1486),
.B(n_1446),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1486),
.B(n_1400),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1405),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1503),
.B(n_1404),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1510),
.A2(n_1427),
.B1(n_1438),
.B2(n_1428),
.C(n_1457),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1474),
.C(n_1473),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1484),
.B(n_1459),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1494),
.B(n_1443),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1513),
.B(n_1469),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1503),
.B(n_1428),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1476),
.C(n_1469),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1494),
.B(n_1432),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1479),
.A2(n_1513),
.B(n_1499),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1494),
.B(n_1432),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1479),
.A2(n_1428),
.B(n_1461),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.B(n_1433),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1492),
.B(n_1426),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1426),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1471),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1500),
.B(n_1433),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1517),
.B(n_1518),
.C(n_1516),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1495),
.A2(n_1455),
.B(n_1444),
.Y(n_1554)
);

NOR3xp33_ASAP7_75t_SL g1555 ( 
.A(n_1509),
.B(n_1332),
.C(n_1392),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1502),
.A2(n_1437),
.B(n_1468),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1493),
.B(n_1439),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1516),
.B(n_1440),
.C(n_1435),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1504),
.B(n_1449),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1490),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1504),
.B(n_1475),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1435),
.C(n_1450),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1497),
.B(n_1498),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1493),
.B(n_1507),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_1467),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1488),
.A2(n_1417),
.B(n_1454),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1507),
.B(n_1409),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1569),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1561),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1478),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1551),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1550),
.B(n_1508),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1560),
.B(n_1483),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1548),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1546),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1562),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1497),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1524),
.B(n_1429),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1542),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1564),
.B(n_1478),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1560),
.B(n_1483),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1498),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1558),
.B(n_1478),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1526),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.B(n_1482),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1566),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1562),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1556),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1563),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1525),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1525),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1522),
.B(n_1485),
.Y(n_1602)
);

AND2x4_ASAP7_75t_SL g1603 ( 
.A(n_1527),
.B(n_1506),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1525),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1556),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1541),
.B(n_1485),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1553),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1557),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1536),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1554),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1589),
.B(n_1533),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1602),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1602),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1606),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1580),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1589),
.B(n_1545),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1572),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1529),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1595),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1595),
.B(n_1530),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1571),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1579),
.B(n_1539),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1571),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1607),
.B(n_1520),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1574),
.B(n_1552),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1603),
.A2(n_1523),
.B1(n_1537),
.B2(n_1532),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1606),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1576),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1575),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1577),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1577),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1607),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1603),
.A2(n_1521),
.B(n_1534),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1608),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1540),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1580),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1576),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1574),
.B(n_1568),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1574),
.B(n_1496),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1574),
.B(n_1496),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1609),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1610),
.B(n_1496),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1581),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1581),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1639),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1637),
.B(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1634),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1622),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1640),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1620),
.C(n_1625),
.D(n_1614),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1643),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1645),
.B(n_1583),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1615),
.B(n_1594),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1648),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1668)
);

NAND2x2_ASAP7_75t_L g1669 ( 
.A(n_1622),
.B(n_1572),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_L g1670 ( 
.A(n_1616),
.B(n_1645),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1613),
.B(n_1578),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1626),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1649),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1578),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1650),
.B(n_1528),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1619),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1626),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1617),
.B(n_1587),
.Y(n_1680)
);

NAND2x2_ASAP7_75t_L g1681 ( 
.A(n_1623),
.B(n_1596),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1641),
.B(n_1587),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1628),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1632),
.B(n_1570),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1628),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1630),
.B(n_1611),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1630),
.B(n_1611),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1618),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1618),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1621),
.Y(n_1690)
);

NAND2x2_ASAP7_75t_L g1691 ( 
.A(n_1616),
.B(n_1596),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1621),
.B(n_1570),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1633),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1633),
.B(n_1590),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1646),
.B(n_1647),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.B(n_1592),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1644),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1688),
.A2(n_1598),
.B(n_1597),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1683),
.B(n_1651),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1664),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1661),
.A2(n_1631),
.B(n_1638),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1678),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1665),
.B(n_1646),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1688),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1664),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1647),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1695),
.B(n_1582),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1679),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1691),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1683),
.B(n_1654),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1668),
.B(n_1651),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1689),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1653),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1662),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1654),
.B(n_1652),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1653),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1690),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1652),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1686),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1675),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1693),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1687),
.B(n_1582),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1670),
.B(n_1582),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1664),
.B(n_1582),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1657),
.B(n_1656),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1659),
.B(n_1596),
.Y(n_1730)
);

AND3x1_ASAP7_75t_L g1731 ( 
.A(n_1657),
.B(n_1584),
.C(n_1649),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1659),
.B(n_1601),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1701),
.A2(n_1677),
.B1(n_1681),
.B2(n_1663),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

OAI322xp33_ASAP7_75t_L g1735 ( 
.A1(n_1716),
.A2(n_1655),
.A3(n_1658),
.B1(n_1672),
.B2(n_1667),
.C1(n_1671),
.C2(n_1684),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1701),
.A2(n_1677),
.B1(n_1681),
.B2(n_1691),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1723),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_SL g1738 ( 
.A1(n_1716),
.A2(n_1696),
.B(n_1610),
.C(n_1694),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_1692),
.B(n_1680),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1702),
.B(n_1673),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1707),
.B(n_1682),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1731),
.A2(n_1669),
.B1(n_1676),
.B2(n_1585),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1723),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1698),
.A2(n_1601),
.B1(n_1669),
.B2(n_1597),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1720),
.A2(n_1601),
.B1(n_1600),
.B2(n_1604),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1707),
.A2(n_1718),
.B1(n_1732),
.B2(n_1713),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1709),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1731),
.B(n_1591),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1710),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_R g1751 ( 
.A(n_1700),
.B(n_1383),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1590),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1717),
.B(n_1583),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1713),
.A2(n_1612),
.B(n_1600),
.C(n_1604),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1698),
.A2(n_1601),
.B1(n_1597),
.B2(n_1605),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1729),
.A2(n_1591),
.B(n_1586),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1723),
.A2(n_1585),
.B1(n_1586),
.B2(n_1591),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1732),
.A2(n_1604),
.B1(n_1600),
.B2(n_1612),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1737),
.B(n_1717),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1743),
.B(n_1703),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1747),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1749),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1750),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1740),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1746),
.B(n_1717),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1746),
.B(n_1724),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1752),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1741),
.B(n_1697),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1770)
);

NAND2x1_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1753),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1739),
.B(n_1724),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1703),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1751),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1738),
.B(n_1724),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1756),
.B(n_1729),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1735),
.B(n_1729),
.Y(n_1778)
);

AOI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1745),
.B(n_1742),
.C(n_1712),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1760),
.B(n_1706),
.Y(n_1780)
);

NOR2x1p5_ASAP7_75t_SL g1781 ( 
.A(n_1769),
.B(n_1704),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1766),
.A2(n_1767),
.B(n_1778),
.C(n_1773),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1776),
.B(n_1777),
.C(n_1765),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1771),
.A2(n_1758),
.B1(n_1744),
.B2(n_1754),
.C(n_1755),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1775),
.A2(n_1698),
.B1(n_1712),
.B2(n_1758),
.Y(n_1785)
);

OAI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1761),
.A2(n_1770),
.B(n_1762),
.C(n_1774),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1760),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1762),
.A2(n_1699),
.B(n_1711),
.C(n_1710),
.Y(n_1788)
);

OA22x2_ASAP7_75t_L g1789 ( 
.A1(n_1774),
.A2(n_1712),
.B1(n_1727),
.B2(n_1757),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1770),
.A2(n_1768),
.B1(n_1772),
.B2(n_1759),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1787),
.Y(n_1791)
);

NAND4xp25_ASAP7_75t_L g1792 ( 
.A(n_1782),
.B(n_1759),
.C(n_1769),
.D(n_1768),
.Y(n_1792)
);

NOR3xp33_ASAP7_75t_L g1793 ( 
.A(n_1786),
.B(n_1762),
.C(n_1763),
.Y(n_1793)
);

NOR3x1_ASAP7_75t_L g1794 ( 
.A(n_1780),
.B(n_1764),
.C(n_1699),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1788),
.B(n_1759),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1779),
.B(n_1704),
.C(n_1700),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1781),
.Y(n_1797)
);

NOR3x1_ASAP7_75t_L g1798 ( 
.A(n_1784),
.B(n_1715),
.C(n_1711),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1790),
.C(n_1785),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1789),
.B(n_1700),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1782),
.B(n_1705),
.C(n_1715),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1792),
.B(n_1705),
.Y(n_1802)
);

NAND4xp75_ASAP7_75t_L g1803 ( 
.A(n_1798),
.B(n_1727),
.C(n_1728),
.D(n_1706),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1791),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1799),
.B(n_1705),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1797),
.A2(n_1705),
.B(n_1411),
.C(n_1445),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1801),
.B(n_1697),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_L g1808 ( 
.A(n_1796),
.B(n_1727),
.C(n_1728),
.D(n_1706),
.Y(n_1808)
);

NOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1795),
.B(n_1800),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1809),
.Y(n_1810)
);

NOR2x1_ASAP7_75t_L g1811 ( 
.A(n_1802),
.B(n_1721),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1807),
.A2(n_1793),
.B1(n_1803),
.B2(n_1806),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1805),
.B(n_1804),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1808),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1802),
.B(n_1794),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1809),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1815),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1810),
.Y(n_1818)
);

AOI21xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1816),
.A2(n_1392),
.B(n_1383),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1811),
.Y(n_1820)
);

AND3x4_ASAP7_75t_L g1821 ( 
.A(n_1813),
.B(n_1732),
.C(n_1425),
.Y(n_1821)
);

AND3x4_ASAP7_75t_L g1822 ( 
.A(n_1812),
.B(n_1732),
.C(n_1429),
.Y(n_1822)
);

INVx5_ASAP7_75t_L g1823 ( 
.A(n_1818),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1820),
.Y(n_1824)
);

NAND2xp33_ASAP7_75t_L g1825 ( 
.A(n_1817),
.B(n_1814),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1825),
.A2(n_1823),
.B1(n_1821),
.B2(n_1822),
.Y(n_1826)
);

NAND5xp2_ASAP7_75t_L g1827 ( 
.A(n_1826),
.B(n_1824),
.C(n_1823),
.D(n_1819),
.E(n_1728),
.Y(n_1827)
);

OA21x2_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1725),
.B(n_1721),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1827),
.A2(n_1719),
.B(n_1725),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1828),
.A2(n_1698),
.B1(n_1732),
.B2(n_1719),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1829),
.A2(n_1722),
.B(n_1697),
.C(n_1714),
.Y(n_1831)
);

OR3x1_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1460),
.C(n_1423),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1831),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1832),
.B(n_1722),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1834),
.A2(n_1722),
.B1(n_1714),
.B2(n_1730),
.Y(n_1835)
);

OAI221xp5_ASAP7_75t_R g1836 ( 
.A1(n_1835),
.A2(n_1730),
.B1(n_1708),
.B2(n_1726),
.C(n_1397),
.Y(n_1836)
);

AOI211xp5_ASAP7_75t_L g1837 ( 
.A1(n_1836),
.A2(n_1298),
.B(n_1360),
.C(n_1337),
.Y(n_1837)
);


endmodule