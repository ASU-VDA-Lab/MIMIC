module real_aes_8110_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g424 ( .A(n_0), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_1), .A2(n_124), .B(n_128), .C(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_2), .A2(n_153), .B(n_154), .Y(n_152) );
INVx1_ASAP7_75t_L g528 ( .A(n_3), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_4), .B(n_165), .Y(n_164) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_5), .A2(n_153), .B(n_495), .Y(n_494) );
AND2x6_ASAP7_75t_L g124 ( .A(n_6), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g270 ( .A(n_7), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_8), .B(n_40), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_9), .A2(n_174), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_10), .B(n_136), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_11), .B(n_158), .Y(n_483) );
INVx1_ASAP7_75t_L g499 ( .A(n_12), .Y(n_499) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g453 ( .A(n_14), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_15), .A2(n_134), .B(n_226), .C(n_228), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_16), .B(n_165), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_17), .B(n_463), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_18), .B(n_153), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_19), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_20), .A2(n_158), .B(n_235), .C(n_237), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_21), .B(n_165), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_22), .B(n_136), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_23), .A2(n_181), .B(n_228), .C(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_24), .B(n_136), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_25), .Y(n_189) );
INVx1_ASAP7_75t_L g132 ( .A(n_26), .Y(n_132) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_27), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_29), .B(n_136), .Y(n_529) );
INVx1_ASAP7_75t_L g179 ( .A(n_30), .Y(n_179) );
INVx1_ASAP7_75t_L g507 ( .A(n_31), .Y(n_507) );
INVx2_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_33), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_34), .A2(n_158), .B(n_159), .C(n_161), .Y(n_157) );
INVxp67_ASAP7_75t_L g180 ( .A(n_35), .Y(n_180) );
CKINVDCx14_ASAP7_75t_R g155 ( .A(n_36), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_37), .A2(n_128), .B(n_131), .C(n_139), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_38), .A2(n_124), .B(n_128), .C(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_39), .A2(n_68), .B1(n_710), .B2(n_711), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_39), .Y(n_710) );
INVx1_ASAP7_75t_L g506 ( .A(n_41), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_42), .A2(n_197), .B(n_268), .C(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_43), .B(n_136), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_44), .A2(n_84), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_44), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_45), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_46), .Y(n_176) );
INVx1_ASAP7_75t_L g233 ( .A(n_47), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_48), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_49), .B(n_153), .Y(n_485) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_50), .A2(n_709), .B1(n_712), .B2(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_50), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_51), .A2(n_128), .B1(n_237), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_52), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_53), .Y(n_525) );
CKINVDCx14_ASAP7_75t_R g266 ( .A(n_54), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_55), .A2(n_161), .B(n_268), .C(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_56), .Y(n_474) );
INVx1_ASAP7_75t_L g496 ( .A(n_57), .Y(n_496) );
INVx1_ASAP7_75t_L g125 ( .A(n_58), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
INVx1_ASAP7_75t_SL g160 ( .A(n_60), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_61), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_62), .B(n_165), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_63), .Y(n_427) );
INVx1_ASAP7_75t_L g192 ( .A(n_64), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_SL g515 ( .A1(n_65), .A2(n_161), .B(n_463), .C(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g517 ( .A(n_66), .Y(n_517) );
INVx1_ASAP7_75t_L g437 ( .A(n_67), .Y(n_437) );
INVx1_ASAP7_75t_L g711 ( .A(n_68), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_69), .A2(n_153), .B(n_265), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_70), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_71), .A2(n_153), .B(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_72), .Y(n_510) );
INVx1_ASAP7_75t_L g468 ( .A(n_73), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_74), .A2(n_174), .B(n_175), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_75), .Y(n_126) );
INVx1_ASAP7_75t_L g224 ( .A(n_76), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_77), .A2(n_124), .B(n_128), .C(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_78), .A2(n_153), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g227 ( .A(n_79), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_80), .B(n_133), .Y(n_461) );
INVx2_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx1_ASAP7_75t_L g216 ( .A(n_82), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_83), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_84), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_85), .A2(n_124), .B(n_128), .C(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g421 ( .A(n_86), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g706 ( .A(n_86), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_86), .B(n_423), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_87), .A2(n_128), .B(n_191), .C(n_199), .Y(n_190) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_88), .A2(n_440), .B1(n_708), .B2(n_714), .C1(n_721), .C2(n_722), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_89), .B(n_140), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_90), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_91), .A2(n_124), .B(n_128), .C(n_481), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_92), .A2(n_103), .B1(n_429), .B2(n_438), .C1(n_725), .C2(n_730), .Y(n_102) );
OAI22xp33_ASAP7_75t_SL g105 ( .A1(n_92), .A2(n_106), .B1(n_417), .B2(n_418), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_92), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_93), .Y(n_487) );
INVx1_ASAP7_75t_L g514 ( .A(n_94), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_95), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_96), .B(n_133), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_97), .B(n_148), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_98), .B(n_148), .Y(n_454) );
INVx2_ASAP7_75t_L g236 ( .A(n_99), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_100), .B(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_101), .A2(n_153), .B(n_513), .Y(n_512) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_419), .B(n_426), .Y(n_104) );
INVx1_ASAP7_75t_L g418 ( .A(n_106), .Y(n_418) );
XOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_110), .A2(n_441), .B1(n_705), .B2(n_707), .Y(n_440) );
INVx1_ASAP7_75t_L g718 ( .A(n_110), .Y(n_718) );
OR3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_328), .C(n_375), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_274), .C(n_299), .Y(n_111) );
AOI221xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_209), .B1(n_240), .B2(n_243), .C(n_251), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_166), .B(n_202), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_115), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_115), .B(n_256), .Y(n_372) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_150), .Y(n_115) );
AND2x2_ASAP7_75t_L g242 ( .A(n_116), .B(n_208), .Y(n_242) );
AND2x2_ASAP7_75t_L g292 ( .A(n_116), .B(n_207), .Y(n_292) );
AND2x2_ASAP7_75t_L g313 ( .A(n_116), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g318 ( .A(n_116), .B(n_285), .Y(n_318) );
OR2x2_ASAP7_75t_L g326 ( .A(n_116), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g398 ( .A(n_116), .B(n_186), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_116), .B(n_347), .Y(n_412) );
INVx3_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g257 ( .A(n_117), .B(n_150), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_117), .B(n_186), .Y(n_258) );
AND2x4_ASAP7_75t_L g280 ( .A(n_117), .B(n_208), .Y(n_280) );
AND2x2_ASAP7_75t_L g310 ( .A(n_117), .B(n_168), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_117), .B(n_309), .Y(n_319) );
AND2x2_ASAP7_75t_L g335 ( .A(n_117), .B(n_187), .Y(n_335) );
OR2x2_ASAP7_75t_L g344 ( .A(n_117), .B(n_327), .Y(n_344) );
AND2x2_ASAP7_75t_L g350 ( .A(n_117), .B(n_285), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_117), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g364 ( .A(n_117), .B(n_204), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_117), .B(n_253), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_117), .B(n_314), .Y(n_403) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_145), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_127), .C(n_140), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_119), .A2(n_189), .B(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_119), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_119), .A2(n_468), .B(n_469), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_119), .A2(n_163), .B1(n_504), .B2(n_508), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_119), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
AND2x4_ASAP7_75t_L g153 ( .A(n_120), .B(n_124), .Y(n_153) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
INVx1_ASAP7_75t_L g238 ( .A(n_122), .Y(n_238) );
INVx1_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
INVx3_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_123), .Y(n_182) );
INVx1_ASAP7_75t_L g463 ( .A(n_123), .Y(n_463) );
BUFx3_ASAP7_75t_L g139 ( .A(n_124), .Y(n_139) );
INVx4_ASAP7_75t_SL g163 ( .A(n_124), .Y(n_163) );
INVx5_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
BUFx3_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_135), .C(n_137), .Y(n_131) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_133), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_133), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_134), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_134), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_134), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
INVx2_ASAP7_75t_L g268 ( .A(n_136), .Y(n_268) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_138), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_140), .A2(n_264), .B(n_271), .Y(n_263) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_140), .A2(n_448), .B(n_454), .Y(n_447) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g149 ( .A(n_141), .B(n_142), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx3_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_147), .A2(n_188), .B(n_200), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_147), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_SL g464 ( .A(n_147), .B(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_148), .A2(n_512), .B(n_518), .Y(n_511) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx2_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
AND2x2_ASAP7_75t_L g309 ( .A(n_150), .B(n_186), .Y(n_309) );
AND2x2_ASAP7_75t_L g314 ( .A(n_150), .B(n_187), .Y(n_314) );
INVx1_ASAP7_75t_L g370 ( .A(n_150), .Y(n_370) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_164), .Y(n_150) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_222), .B(n_229), .Y(n_221) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_151), .A2(n_231), .B(n_239), .Y(n_230) );
BUFx2_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_157), .C(n_163), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_156), .A2(n_163), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_156), .A2(n_163), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_156), .A2(n_163), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_156), .A2(n_163), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_156), .A2(n_163), .B(n_450), .C(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_156), .A2(n_163), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_156), .A2(n_163), .B(n_514), .C(n_515), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_158), .B(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_162), .Y(n_484) );
INVx1_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_165), .A2(n_494), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g279 ( .A(n_167), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_186), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_168), .B(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g256 ( .A(n_168), .Y(n_256) );
OR2x2_ASAP7_75t_L g327 ( .A(n_168), .B(n_186), .Y(n_327) );
OR2x2_ASAP7_75t_L g388 ( .A(n_168), .B(n_295), .Y(n_388) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_183), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_205), .B(n_206), .Y(n_204) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_170), .A2(n_467), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_SL g457 ( .A1(n_171), .A2(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_172), .A2(n_503), .B(n_509), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_172), .B(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_172), .A2(n_524), .B(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g205 ( .A(n_173), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_181), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_181), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_181), .B(n_453), .Y(n_452) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g194 ( .A(n_182), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_182), .A2(n_194), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_185), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_185), .A2(n_479), .B(n_486), .Y(n_478) );
AND2x2_ASAP7_75t_L g207 ( .A(n_186), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g347 ( .A(n_186), .B(n_204), .Y(n_347) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g286 ( .A(n_187), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_193), .A2(n_196), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_196), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_196), .A2(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g228 ( .A(n_198), .Y(n_228) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_203), .A2(n_392), .B1(n_396), .B2(n_399), .C(n_400), .Y(n_391) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_207), .Y(n_203) );
INVx1_ASAP7_75t_SL g254 ( .A(n_204), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_204), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g386 ( .A(n_204), .B(n_242), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_207), .B(n_256), .Y(n_378) );
AND2x2_ASAP7_75t_L g285 ( .A(n_208), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g289 ( .A(n_209), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_209), .B(n_295), .Y(n_325) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AND2x2_ASAP7_75t_L g250 ( .A(n_210), .B(n_221), .Y(n_250) );
INVx4_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
BUFx3_ASAP7_75t_L g305 ( .A(n_210), .Y(n_305) );
AND3x2_ASAP7_75t_L g320 ( .A(n_210), .B(n_321), .C(n_322), .Y(n_320) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_211), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_211), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_211), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g402 ( .A(n_220), .B(n_316), .Y(n_402) );
AND2x2_ASAP7_75t_L g410 ( .A(n_220), .B(n_295), .Y(n_410) );
INVx1_ASAP7_75t_SL g415 ( .A(n_220), .Y(n_415) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
INVx1_ASAP7_75t_SL g273 ( .A(n_221), .Y(n_273) );
AND2x2_ASAP7_75t_L g296 ( .A(n_221), .B(n_262), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_221), .B(n_246), .Y(n_298) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_221), .Y(n_338) );
OR2x2_ASAP7_75t_L g343 ( .A(n_221), .B(n_262), .Y(n_343) );
INVx2_ASAP7_75t_L g248 ( .A(n_230), .Y(n_248) );
AND2x2_ASAP7_75t_L g283 ( .A(n_230), .B(n_263), .Y(n_283) );
OR2x2_ASAP7_75t_L g303 ( .A(n_230), .B(n_263), .Y(n_303) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_230), .Y(n_323) );
INVx2_ASAP7_75t_L g530 ( .A(n_237), .Y(n_530) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_241), .A2(n_282), .B(n_374), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g409 ( .A1(n_243), .A2(n_253), .A3(n_280), .B1(n_410), .B2(n_411), .C1(n_413), .C2(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_245), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_246), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g340 ( .A(n_248), .B(n_262), .Y(n_340) );
AND2x2_ASAP7_75t_L g407 ( .A(n_248), .B(n_263), .Y(n_407) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g348 ( .A(n_250), .B(n_302), .Y(n_348) );
AOI31xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_255), .A3(n_258), .B(n_259), .Y(n_251) );
AND2x2_ASAP7_75t_L g307 ( .A(n_253), .B(n_285), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_253), .B(n_277), .Y(n_389) );
AND2x2_ASAP7_75t_L g408 ( .A(n_253), .B(n_313), .Y(n_408) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_256), .B(n_285), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_256), .B(n_314), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_256), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_256), .B(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_257), .B(n_314), .Y(n_346) );
INVx1_ASAP7_75t_L g390 ( .A(n_257), .Y(n_390) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_272), .Y(n_260) );
INVxp67_ASAP7_75t_L g342 ( .A(n_261), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_262), .B(n_273), .Y(n_278) );
INVx1_ASAP7_75t_L g384 ( .A(n_262), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_262), .B(n_361), .Y(n_395) );
BUFx3_ASAP7_75t_L g295 ( .A(n_263), .Y(n_295) );
AND2x2_ASAP7_75t_L g321 ( .A(n_263), .B(n_273), .Y(n_321) );
INVx2_ASAP7_75t_L g361 ( .A(n_263), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_272), .B(n_394), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_281), .C(n_290), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_276), .A2(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_277), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_277), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g357 ( .A(n_278), .B(n_303), .Y(n_357) );
INVx3_ASAP7_75t_L g288 ( .A(n_280), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_284), .B1(n_287), .B2(n_289), .Y(n_281) );
OAI21xp5_ASAP7_75t_SL g306 ( .A1(n_283), .A2(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g332 ( .A(n_283), .B(n_296), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_283), .B(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g287 ( .A(n_286), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g356 ( .A(n_286), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g300 ( .A1(n_287), .A2(n_301), .B(n_306), .Y(n_300) );
OAI22xp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B1(n_297), .B2(n_298), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_292), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_338), .Y(n_337) );
NOR3xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_311), .C(n_324), .Y(n_299) );
OAI22xp5_ASAP7_75t_SL g366 ( .A1(n_301), .A2(n_367), .B1(n_371), .B2(n_372), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g371 ( .A(n_303), .B(n_304), .Y(n_371) );
AND2x2_ASAP7_75t_L g379 ( .A(n_304), .B(n_360), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_305), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_SL g387 ( .A1(n_305), .A2(n_388), .B(n_389), .C(n_390), .Y(n_387) );
OR2x2_ASAP7_75t_L g414 ( .A(n_305), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B(n_317), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_313), .A2(n_350), .B(n_351), .C(n_354), .Y(n_349) );
OAI21xp33_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g382 ( .A(n_321), .B(n_340), .Y(n_382) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
NAND3xp33_ASAP7_75t_SL g328 ( .A(n_329), .B(n_349), .C(n_362), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_333), .C(n_341), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g399 ( .A(n_336), .Y(n_399) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_338), .B(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_344), .C(n_345), .Y(n_341) );
INVx2_ASAP7_75t_SL g353 ( .A(n_343), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_344), .A2(n_355), .B1(n_357), .B2(n_358), .Y(n_354) );
OAI21xp33_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_366), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVxp33_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
NAND4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_391), .C(n_404), .D(n_409), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .C(n_387), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_385), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_381), .A2(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_388), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_420), .A2(n_434), .B(n_435), .Y(n_731) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_421), .Y(n_428) );
INVx1_ASAP7_75t_SL g729 ( .A(n_421), .Y(n_729) );
NOR2x2_ASAP7_75t_L g724 ( .A(n_422), .B(n_706), .Y(n_724) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g705 ( .A(n_423), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
CKINVDCx6p67_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_SL g727 ( .A(n_434), .B(n_436), .Y(n_727) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g715 ( .A(n_441), .Y(n_715) );
OR4x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_601), .C(n_660), .D(n_687), .Y(n_441) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_543), .C(n_568), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_475), .B(n_492), .C(n_519), .Y(n_443) );
AOI211xp5_ASAP7_75t_SL g691 ( .A1(n_444), .A2(n_692), .B(n_694), .C(n_697), .Y(n_691) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .Y(n_444) );
INVx1_ASAP7_75t_L g566 ( .A(n_445), .Y(n_566) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g541 ( .A(n_446), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g573 ( .A(n_446), .Y(n_573) );
AND2x2_ASAP7_75t_L g628 ( .A(n_446), .B(n_597), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_446), .B(n_490), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_446), .B(n_491), .Y(n_686) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g547 ( .A(n_447), .Y(n_547) );
AND2x2_ASAP7_75t_L g590 ( .A(n_447), .B(n_466), .Y(n_590) );
AND2x2_ASAP7_75t_L g608 ( .A(n_447), .B(n_491), .Y(n_608) );
INVx4_ASAP7_75t_L g540 ( .A(n_455), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_455), .A2(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g676 ( .A(n_455), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .Y(n_455) );
INVx1_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_491), .Y(n_545) );
OR2x2_ASAP7_75t_L g574 ( .A(n_456), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g588 ( .A(n_456), .Y(n_588) );
INVx3_ASAP7_75t_L g597 ( .A(n_456), .Y(n_597) );
AND2x2_ASAP7_75t_L g607 ( .A(n_456), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_456), .B(n_546), .Y(n_640) );
AND2x2_ASAP7_75t_L g664 ( .A(n_456), .B(n_620), .Y(n_664) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
AND2x2_ASAP7_75t_L g700 ( .A(n_466), .B(n_542), .Y(n_700) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_488), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_477), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_608), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_477), .B(n_597), .Y(n_682) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
AND2x2_ASAP7_75t_L g546 ( .A(n_478), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g587 ( .A(n_478), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_485), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_488), .B(n_583), .Y(n_605) );
INVx1_ASAP7_75t_L g644 ( .A(n_488), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_488), .B(n_571), .Y(n_688) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g551 ( .A(n_489), .B(n_546), .Y(n_551) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_491), .B(n_542), .Y(n_575) );
INVx1_ASAP7_75t_L g654 ( .A(n_491), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_492), .A2(n_593), .A3(n_653), .B1(n_679), .B2(n_681), .C1(n_683), .C2(n_685), .Y(n_678) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_493), .B(n_501), .Y(n_492) );
AND2x2_ASAP7_75t_L g533 ( .A(n_493), .B(n_511), .Y(n_533) );
INVx1_ASAP7_75t_SL g536 ( .A(n_493), .Y(n_536) );
AND2x2_ASAP7_75t_L g538 ( .A(n_493), .B(n_502), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_493), .B(n_555), .Y(n_561) );
INVx2_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_493), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g631 ( .A(n_493), .B(n_555), .Y(n_631) );
BUFx2_ASAP7_75t_L g648 ( .A(n_493), .Y(n_648) );
AND2x2_ASAP7_75t_L g662 ( .A(n_493), .B(n_522), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_501), .B(n_550), .Y(n_577) );
AND2x2_ASAP7_75t_L g704 ( .A(n_501), .B(n_580), .Y(n_704) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
OR2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g555 ( .A(n_502), .Y(n_555) );
AND2x2_ASAP7_75t_L g600 ( .A(n_502), .B(n_523), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_502), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_502), .Y(n_684) );
AND2x2_ASAP7_75t_L g535 ( .A(n_511), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g557 ( .A(n_511), .Y(n_557) );
BUFx2_ASAP7_75t_L g563 ( .A(n_511), .Y(n_563) );
AND2x2_ASAP7_75t_L g582 ( .A(n_511), .B(n_555), .Y(n_582) );
INVx3_ASAP7_75t_L g594 ( .A(n_511), .Y(n_594) );
OR2x2_ASAP7_75t_L g604 ( .A(n_511), .B(n_555), .Y(n_604) );
AOI31xp33_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_534), .A3(n_537), .B(n_539), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_521), .B(n_556), .Y(n_567) );
OR2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_561), .Y(n_591) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_522), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g612 ( .A(n_522), .B(n_604), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_522), .B(n_594), .Y(n_622) );
AND2x2_ASAP7_75t_L g629 ( .A(n_522), .B(n_630), .Y(n_629) );
NAND2x1_ASAP7_75t_L g657 ( .A(n_522), .B(n_593), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_522), .B(n_648), .Y(n_658) );
AND2x2_ASAP7_75t_L g670 ( .A(n_522), .B(n_555), .Y(n_670) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g550 ( .A(n_523), .Y(n_550) );
INVx1_ASAP7_75t_L g616 ( .A(n_533), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_533), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_535), .B(n_611), .Y(n_645) );
AND2x4_ASAP7_75t_L g556 ( .A(n_536), .B(n_557), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g635 ( .A(n_541), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_541), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g583 ( .A(n_542), .B(n_573), .Y(n_583) );
AND2x2_ASAP7_75t_L g677 ( .A(n_542), .B(n_547), .Y(n_677) );
INVx1_ASAP7_75t_L g702 ( .A(n_542), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_548), .B1(n_551), .B2(n_552), .C(n_558), .Y(n_543) );
CKINVDCx14_ASAP7_75t_R g564 ( .A(n_544), .Y(n_564) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_545), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_548), .B(n_599), .Y(n_618) );
INVx3_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g667 ( .A(n_549), .B(n_563), .Y(n_667) );
AND2x2_ASAP7_75t_L g581 ( .A(n_550), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g611 ( .A(n_550), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_550), .B(n_594), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_550), .B(n_651), .C(n_682), .Y(n_681) );
AOI211xp5_ASAP7_75t_SL g614 ( .A1(n_551), .A2(n_615), .B(n_617), .C(n_625), .Y(n_614) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_553), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_554), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_554), .B(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g696 ( .A(n_556), .B(n_670), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B1(n_565), .B2(n_567), .Y(n_558) );
NOR2xp33_ASAP7_75t_SL g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_562), .B(n_611), .Y(n_642) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_565), .A2(n_657), .B1(n_688), .B2(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_576), .B1(n_578), .B2(n_583), .C(n_584), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_574), .A2(n_585), .B1(n_591), .B2(n_592), .C(n_595), .Y(n_584) );
INVx1_ASAP7_75t_L g627 ( .A(n_575), .Y(n_627) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_SL g599 ( .A(n_580), .Y(n_599) );
OR2x2_ASAP7_75t_L g672 ( .A(n_580), .B(n_604), .Y(n_672) );
AND2x2_ASAP7_75t_L g674 ( .A(n_580), .B(n_582), .Y(n_674) );
INVx1_ASAP7_75t_L g613 ( .A(n_583), .Y(n_613) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_586), .A2(n_644), .B(n_645), .Y(n_643) );
OR2x2_ASAP7_75t_L g650 ( .A(n_586), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g624 ( .A(n_587), .B(n_608), .Y(n_624) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp33_ASAP7_75t_SL g641 ( .A(n_592), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_593), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_594), .B(n_630), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_597), .A2(n_610), .B(n_612), .C(n_613), .Y(n_609) );
NAND2x1_ASAP7_75t_SL g634 ( .A(n_597), .B(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_647), .B1(n_649), .B2(n_652), .Y(n_646) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_600), .B(n_690), .Y(n_689) );
NAND5xp2_ASAP7_75t_L g601 ( .A(n_602), .B(n_614), .C(n_632), .D(n_646), .E(n_655), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_609), .Y(n_602) );
INVx1_ASAP7_75t_L g659 ( .A(n_605), .Y(n_659) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_607), .A2(n_626), .B1(n_666), .B2(n_668), .C(n_671), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_608), .B(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_611), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_611), .B(n_677), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_621), .B2(n_623), .Y(n_617) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g699 ( .A(n_628), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_640), .B2(n_641), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g683 ( .A(n_638), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g690 ( .A(n_648), .Y(n_690) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_658), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_665), .C(n_678), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_663), .A2(n_688), .B(n_689), .C(n_691), .Y(n_687) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_667), .B(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B(n_703), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g717 ( .A(n_705), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_707), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_708), .Y(n_721) );
INVx1_ASAP7_75t_L g712 ( .A(n_709), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B1(n_718), .B2(n_719), .Y(n_714) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
NAND2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
endmodule