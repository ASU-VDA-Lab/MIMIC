module fake_ariane_1998_n_1394 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1394);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1394;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_163),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_162),
.B(n_42),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_213),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_158),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_153),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_63),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_70),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_211),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_209),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_92),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_95),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_237),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_111),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_152),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_200),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_52),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_86),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_107),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_118),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_182),
.B(n_5),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_273),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_130),
.B(n_119),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_279),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_120),
.B(n_161),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_185),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_93),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_25),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_156),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_271),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_131),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_328),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_98),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_189),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_30),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_125),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_64),
.B(n_50),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_154),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_194),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_170),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_145),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_116),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_266),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_91),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_72),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_226),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_260),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_212),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_303),
.B(n_278),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_308),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_26),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_183),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_70),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_242),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_29),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_270),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_148),
.B(n_252),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_199),
.B(n_236),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_53),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_206),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_291),
.B(n_180),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_123),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_43),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_171),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_151),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_128),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_172),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_198),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_173),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_338),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_62),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_147),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_201),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_191),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_344),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_197),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_106),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_346),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_32),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_14),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_277),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_60),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_195),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_30),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_310),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_274),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_51),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_38),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_48),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_221),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_0),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_347),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_210),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_18),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_132),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_240),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_7),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_103),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_55),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_290),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_165),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_129),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_141),
.B(n_321),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_230),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_17),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_269),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_202),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_13),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_176),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_224),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_13),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_133),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_51),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_207),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_77),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_104),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_34),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_302),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_336),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_135),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_174),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_20),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_166),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_218),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_251),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_287),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_317),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_208),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_155),
.B(n_267),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_216),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_311),
.B(n_84),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_259),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_127),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_18),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_43),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_301),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_80),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_50),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_222),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_298),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_83),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_312),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_367),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_371),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_367),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_367),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_361),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_361),
.B(n_0),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_403),
.B(n_1),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_400),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_513)
);

BUFx8_ASAP7_75t_L g514 ( 
.A(n_385),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_360),
.B(n_402),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_444),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_372),
.B(n_2),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_444),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_462),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_456),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_456),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_462),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_413),
.B(n_3),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_456),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_372),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_4),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_439),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_476),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_351),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_496),
.Y(n_533)
);

NOR2x1_ASAP7_75t_L g534 ( 
.A(n_355),
.B(n_121),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_407),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_363),
.B(n_10),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_373),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_352),
.B(n_11),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_382),
.Y(n_541)
);

AOI22x1_ASAP7_75t_R g542 ( 
.A1(n_388),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_390),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_360),
.A2(n_124),
.B(n_122),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_353),
.B(n_16),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_411),
.B(n_19),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_474),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_349),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_448),
.B(n_21),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_421),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_408),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_362),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_356),
.B(n_22),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_421),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_501),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_369),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_376),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_357),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_470),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_434),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_395),
.Y(n_566)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_364),
.A2(n_26),
.B(n_27),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_365),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_384),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_468),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_468),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

AND2x2_ASAP7_75t_SL g576 ( 
.A(n_440),
.B(n_27),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_374),
.Y(n_577)
);

OAI22x1_ASAP7_75t_R g578 ( 
.A1(n_381),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_463),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_472),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_420),
.A2(n_33),
.B1(n_28),
.B2(n_31),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_397),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_559),
.B(n_460),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_502),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_R g587 ( 
.A(n_504),
.B(n_412),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_515),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_583),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_535),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_538),
.B(n_368),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_538),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_512),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_511),
.B(n_536),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_535),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_530),
.B(n_359),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_554),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_568),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_511),
.B(n_359),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_536),
.B(n_405),
.Y(n_605)
);

BUFx6f_ASAP7_75t_SL g606 ( 
.A(n_576),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_570),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_577),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_551),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_579),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_552),
.B(n_475),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_581),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_561),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_515),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_551),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_404),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_503),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_517),
.A2(n_493),
.B1(n_494),
.B2(n_392),
.Y(n_621)
);

NOR2x1p5_ASAP7_75t_L g622 ( 
.A(n_519),
.B(n_416),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_553),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_553),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_561),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_552),
.A2(n_509),
.B1(n_545),
.B2(n_540),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_553),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_560),
.B(n_466),
.C(n_420),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_566),
.B(n_378),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_558),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_520),
.B(n_523),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_539),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_600),
.A2(n_576),
.B1(n_524),
.B2(n_527),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_SL g636 ( 
.A(n_600),
.B(n_529),
.C(n_513),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_503),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_621),
.A2(n_567),
.B1(n_509),
.B2(n_527),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_586),
.B(n_548),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_620),
.B(n_524),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_586),
.B(n_548),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_537),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_623),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_593),
.B(n_533),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_545),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_SL g646 ( 
.A(n_630),
.B(n_556),
.C(n_550),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_605),
.B(n_549),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_631),
.B(n_557),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_594),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_618),
.B(n_505),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_605),
.B(n_543),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_604),
.B(n_506),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_621),
.B(n_514),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_602),
.B(n_514),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_597),
.A2(n_560),
.B1(n_550),
.B2(n_556),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_633),
.B(n_526),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_508),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_602),
.B(n_591),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_529),
.C(n_513),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_592),
.B(n_547),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_591),
.B(n_436),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_629),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_591),
.B(n_452),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_585),
.B(n_555),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_582),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_612),
.B(n_516),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_629),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_619),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_625),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_612),
.B(n_531),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_607),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_612),
.B(n_609),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_622),
.B(n_354),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_611),
.B(n_518),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_608),
.Y(n_676)
);

NAND2x1_ASAP7_75t_L g677 ( 
.A(n_589),
.B(n_567),
.Y(n_677)
);

AND2x6_ASAP7_75t_SL g678 ( 
.A(n_613),
.B(n_578),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_599),
.B(n_455),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_614),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_626),
.B(n_521),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_626),
.B(n_632),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_626),
.B(n_522),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_632),
.B(n_525),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_634),
.B(n_532),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_606),
.A2(n_528),
.B1(n_423),
.B2(n_426),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_589),
.B(n_603),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_589),
.B(n_603),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_603),
.B(n_558),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_SL g690 ( 
.A(n_606),
.B(n_528),
.C(n_441),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_595),
.B(n_610),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_610),
.B(n_616),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_614),
.B(n_562),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_627),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_624),
.B(n_571),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_627),
.B(n_563),
.Y(n_696)
);

INVx8_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_640),
.B(n_391),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_676),
.B(n_569),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_640),
.B(n_660),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_657),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_647),
.B(n_569),
.Y(n_702)
);

AOI21x1_ASAP7_75t_L g703 ( 
.A1(n_677),
.A2(n_544),
.B(n_534),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_648),
.A2(n_480),
.B(n_405),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_660),
.B(n_422),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_687),
.A2(n_615),
.B(n_406),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_642),
.B(n_429),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_642),
.B(n_442),
.Y(n_708)
);

AO22x1_ASAP7_75t_L g709 ( 
.A1(n_659),
.A2(n_542),
.B1(n_358),
.B2(n_445),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_688),
.A2(n_615),
.B(n_406),
.Y(n_710)
);

INVx6_ASAP7_75t_L g711 ( 
.A(n_671),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_643),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_635),
.B(n_399),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_682),
.A2(n_377),
.B(n_380),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_658),
.B(n_427),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_651),
.B(n_432),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_639),
.A2(n_389),
.B(n_386),
.Y(n_717)
);

AND2x2_ASAP7_75t_SL g718 ( 
.A(n_686),
.B(n_488),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_641),
.A2(n_689),
.B(n_673),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_638),
.A2(n_655),
.B1(n_656),
.B2(n_649),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_651),
.B(n_464),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_664),
.B(n_478),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_685),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_697),
.A2(n_396),
.B(n_394),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_664),
.B(n_483),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_662),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_675),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_696),
.B(n_582),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_644),
.B(n_481),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_680),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_667),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_694),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_670),
.B(n_672),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_497),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_661),
.B(n_500),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_563),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_666),
.B(n_652),
.Y(n_738)
);

AO22x1_ASAP7_75t_L g739 ( 
.A1(n_659),
.A2(n_542),
.B1(n_587),
.B2(n_565),
.Y(n_739)
);

AO32x2_ASAP7_75t_L g740 ( 
.A1(n_636),
.A2(n_490),
.A3(n_375),
.B1(n_350),
.B2(n_587),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_668),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_669),
.Y(n_742)
);

BUFx4_ASAP7_75t_SL g743 ( 
.A(n_678),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_564),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_646),
.A2(n_417),
.B1(n_419),
.B2(n_409),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_681),
.A2(n_684),
.B(n_683),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_636),
.A2(n_418),
.B1(n_431),
.B2(n_430),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_679),
.B(n_387),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_691),
.Y(n_749)
);

BUFx12f_ASAP7_75t_L g750 ( 
.A(n_665),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_674),
.B(n_393),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_654),
.B(n_575),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_692),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_695),
.A2(n_450),
.B(n_447),
.Y(n_754)
);

AO32x1_ASAP7_75t_L g755 ( 
.A1(n_646),
.A2(n_453),
.A3(n_465),
.B1(n_458),
.B2(n_451),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_690),
.A2(n_471),
.B(n_467),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_665),
.B(n_580),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_665),
.B(n_473),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_635),
.A2(n_482),
.B1(n_484),
.B2(n_477),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_487),
.B1(n_491),
.B2(n_486),
.Y(n_760)
);

BUFx8_ASAP7_75t_SL g761 ( 
.A(n_680),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_647),
.B(n_492),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_680),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_645),
.A2(n_414),
.B(n_415),
.C(n_379),
.Y(n_764)
);

OR2x6_ASAP7_75t_SL g765 ( 
.A(n_680),
.B(n_425),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

BUFx2_ASAP7_75t_SL g767 ( 
.A(n_676),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_673),
.B(n_617),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_645),
.A2(n_370),
.B(n_499),
.C(n_479),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_635),
.A2(n_435),
.B1(n_438),
.B2(n_433),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_640),
.B(n_449),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_640),
.B(n_454),
.Y(n_772)
);

NOR2x1_ASAP7_75t_L g773 ( 
.A(n_658),
.B(n_366),
.Y(n_773)
);

BUFx8_ASAP7_75t_L g774 ( 
.A(n_676),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_671),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_657),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_676),
.B(n_33),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_676),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_657),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_657),
.Y(n_780)
);

INVx3_ASAP7_75t_SL g781 ( 
.A(n_680),
.Y(n_781)
);

AOI21xp33_ASAP7_75t_L g782 ( 
.A1(n_645),
.A2(n_424),
.B(n_383),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_657),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_640),
.B(n_489),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_671),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_637),
.A2(n_495),
.B(n_461),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_761),
.B(n_443),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_699),
.B(n_34),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_742),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_763),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_781),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_778),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_711),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_734),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_703),
.A2(n_468),
.B(n_126),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_767),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_729),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_774),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_702),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_731),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_729),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_SL g802 ( 
.A1(n_728),
.A2(n_35),
.B(n_36),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_762),
.A2(n_596),
.B1(n_588),
.B2(n_574),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_698),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_746),
.A2(n_710),
.B(n_706),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_733),
.B(n_596),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_760),
.A2(n_574),
.B(n_572),
.C(n_39),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_722),
.B(n_37),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_711),
.B(n_38),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_741),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_771),
.A2(n_136),
.B(n_134),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_714),
.A2(n_138),
.B(n_137),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_705),
.B(n_39),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_772),
.A2(n_140),
.B(n_139),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_784),
.A2(n_143),
.B(n_142),
.Y(n_815)
);

OAI21x1_ASAP7_75t_SL g816 ( 
.A1(n_720),
.A2(n_40),
.B(n_41),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_745),
.A2(n_44),
.B(n_40),
.C(n_42),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_725),
.B(n_44),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_716),
.B(n_707),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_708),
.B(n_45),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_713),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_712),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_SL g823 ( 
.A1(n_724),
.A2(n_146),
.B(n_144),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_749),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_704),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_701),
.B(n_54),
.Y(n_826)
);

AO32x2_ASAP7_75t_L g827 ( 
.A1(n_747),
.A2(n_56),
.A3(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_751),
.A2(n_150),
.B(n_149),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_752),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_775),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_753),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_765),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_758),
.A2(n_65),
.B(n_61),
.C(n_63),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_718),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_766),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_776),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_738),
.A2(n_735),
.B(n_786),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_775),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

CKINVDCx6p67_ASAP7_75t_R g840 ( 
.A(n_785),
.Y(n_840)
);

AO31x2_ASAP7_75t_L g841 ( 
.A1(n_756),
.A2(n_159),
.A3(n_160),
.B(n_157),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_779),
.B(n_67),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_730),
.A2(n_783),
.B(n_780),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_721),
.B(n_68),
.Y(n_844)
);

AO32x2_ASAP7_75t_L g845 ( 
.A1(n_770),
.A2(n_68),
.A3(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_727),
.B(n_73),
.Y(n_846)
);

BUFx10_ASAP7_75t_L g847 ( 
.A(n_715),
.Y(n_847)
);

AO32x2_ASAP7_75t_L g848 ( 
.A1(n_740),
.A2(n_74),
.A3(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_717),
.A2(n_167),
.B(n_164),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_769),
.A2(n_169),
.B(n_168),
.Y(n_851)
);

AO32x2_ASAP7_75t_L g852 ( 
.A1(n_740),
.A2(n_75),
.A3(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_736),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_853)
);

INVx8_ASAP7_75t_L g854 ( 
.A(n_750),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_768),
.A2(n_177),
.B(n_175),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_757),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_726),
.Y(n_857)
);

AOI22x1_ASAP7_75t_SL g858 ( 
.A1(n_743),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_785),
.Y(n_859)
);

BUFx4_ASAP7_75t_SL g860 ( 
.A(n_737),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_754),
.A2(n_179),
.B(n_178),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_785),
.B(n_81),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_748),
.A2(n_184),
.B(n_181),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_744),
.B(n_82),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_732),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_740),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_773),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_739),
.Y(n_868)
);

BUFx4_ASAP7_75t_R g869 ( 
.A(n_709),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_755),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_755),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_700),
.B(n_85),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_SL g873 ( 
.A1(n_720),
.A2(n_188),
.B(n_187),
.Y(n_873)
);

OAI22x1_ASAP7_75t_L g874 ( 
.A1(n_728),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_700),
.B(n_87),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_700),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_763),
.B(n_90),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_91),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_SL g879 ( 
.A(n_760),
.B(n_92),
.C(n_93),
.Y(n_879)
);

AOI221x1_ASAP7_75t_L g880 ( 
.A1(n_782),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_700),
.B(n_94),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_700),
.B(n_96),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_699),
.B(n_97),
.Y(n_883)
);

INVx3_ASAP7_75t_SL g884 ( 
.A(n_781),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_699),
.B(n_99),
.Y(n_885)
);

AOI221x1_ASAP7_75t_L g886 ( 
.A1(n_782),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.C(n_103),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_778),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_700),
.A2(n_192),
.B(n_190),
.Y(n_888)
);

INVx3_ASAP7_75t_SL g889 ( 
.A(n_781),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_700),
.A2(n_196),
.B(n_193),
.Y(n_890)
);

INVx3_ASAP7_75t_SL g891 ( 
.A(n_781),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_767),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_734),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_734),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_700),
.B(n_101),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_700),
.B(n_102),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_700),
.B(n_104),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_719),
.A2(n_205),
.B(n_204),
.Y(n_898)
);

AOI21x1_ASAP7_75t_SL g899 ( 
.A1(n_700),
.A2(n_105),
.B(n_106),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_699),
.B(n_105),
.Y(n_900)
);

AOI21x1_ASAP7_75t_SL g901 ( 
.A1(n_700),
.A2(n_107),
.B(n_108),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_734),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_699),
.B(n_108),
.Y(n_903)
);

AO32x2_ASAP7_75t_L g904 ( 
.A1(n_759),
.A2(n_109),
.A3(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_778),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_767),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_702),
.B(n_109),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_702),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_761),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_700),
.B(n_110),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_700),
.B(n_112),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_700),
.B(n_113),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_734),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_699),
.B(n_114),
.Y(n_914)
);

INVx6_ASAP7_75t_L g915 ( 
.A(n_774),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_699),
.B(n_114),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_700),
.B(n_115),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_734),
.Y(n_918)
);

AOI221xp5_ASAP7_75t_SL g919 ( 
.A1(n_759),
.A2(n_117),
.B1(n_118),
.B2(n_214),
.C(n_215),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_792),
.B(n_217),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_835),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_907),
.B(n_219),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_794),
.B(n_220),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_836),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_824),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_831),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_819),
.A2(n_223),
.B(n_225),
.Y(n_927)
);

AO21x2_ASAP7_75t_L g928 ( 
.A1(n_837),
.A2(n_227),
.B(n_228),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_849),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_872),
.A2(n_229),
.B(n_231),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_810),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_893),
.B(n_232),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_894),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_822),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_799),
.B(n_348),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_902),
.Y(n_936)
);

AO31x2_ASAP7_75t_L g937 ( 
.A1(n_871),
.A2(n_233),
.A3(n_234),
.B(n_235),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_793),
.B(n_238),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_791),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_875),
.A2(n_239),
.B(n_241),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_913),
.B(n_243),
.Y(n_941)
);

OA21x2_ASAP7_75t_L g942 ( 
.A1(n_805),
.A2(n_244),
.B(n_245),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_918),
.B(n_246),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_826),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_808),
.A2(n_247),
.B(n_248),
.C(n_249),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_865),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_878),
.A2(n_250),
.B(n_253),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_842),
.Y(n_948)
);

NOR2x1_ASAP7_75t_R g949 ( 
.A(n_915),
.B(n_254),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_846),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_816),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_881),
.A2(n_255),
.B(n_257),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_882),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_908),
.B(n_258),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_884),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_844),
.A2(n_261),
.B(n_262),
.C(n_263),
.Y(n_957)
);

AOI21xp33_ASAP7_75t_L g958 ( 
.A1(n_818),
.A2(n_264),
.B(n_265),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_905),
.Y(n_960)
);

AO31x2_ASAP7_75t_L g961 ( 
.A1(n_851),
.A2(n_272),
.A3(n_275),
.B(n_276),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_896),
.A2(n_280),
.B(n_281),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_897),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_788),
.B(n_343),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_910),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_885),
.B(n_282),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_898),
.A2(n_283),
.B(n_284),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_889),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_911),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_791),
.B(n_285),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_830),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_912),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_917),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_843),
.A2(n_286),
.B(n_288),
.C(n_289),
.Y(n_975)
);

BUFx2_ASAP7_75t_SL g976 ( 
.A(n_909),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_800),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_812),
.A2(n_293),
.B(n_294),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_829),
.B(n_295),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_838),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_915),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_820),
.A2(n_296),
.B(n_297),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_856),
.B(n_859),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_860),
.Y(n_984)
);

BUFx2_ASAP7_75t_R g985 ( 
.A(n_891),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_855),
.A2(n_299),
.B(n_300),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_797),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_840),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_813),
.A2(n_304),
.B(n_305),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_848),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_919),
.A2(n_306),
.B(n_309),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_848),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_790),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_313),
.B(n_314),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_864),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_852),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_868),
.Y(n_998)
);

AO21x2_ASAP7_75t_L g999 ( 
.A1(n_861),
.A2(n_315),
.B(n_316),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_883),
.B(n_318),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_834),
.A2(n_319),
.B(n_320),
.C(n_322),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_814),
.A2(n_323),
.B(n_324),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_821),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_815),
.A2(n_325),
.B(n_326),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_900),
.B(n_327),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_852),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_873),
.A2(n_330),
.B(n_331),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_879),
.A2(n_796),
.B1(n_906),
.B2(n_892),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_790),
.Y(n_1009)
);

OA21x2_ASAP7_75t_L g1010 ( 
.A1(n_828),
.A2(n_332),
.B(n_333),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_839),
.B(n_797),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_903),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_914),
.B(n_341),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_867),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_801),
.B(n_798),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_888),
.A2(n_890),
.B(n_899),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_901),
.A2(n_863),
.B(n_850),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_916),
.B(n_847),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_802),
.B(n_874),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_854),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_823),
.A2(n_803),
.B(n_853),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_870),
.A2(n_886),
.B(n_880),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_804),
.A2(n_825),
.B(n_876),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_817),
.A2(n_833),
.B(n_807),
.Y(n_1024)
);

OA21x2_ASAP7_75t_L g1025 ( 
.A1(n_841),
.A2(n_827),
.B(n_862),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_787),
.B(n_854),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_827),
.A2(n_845),
.B(n_904),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_809),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_904),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_809),
.B(n_877),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_845),
.A2(n_869),
.B(n_832),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_795),
.B(n_805),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_792),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_791),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_794),
.B(n_893),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_810),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_799),
.B(n_702),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_791),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_794),
.B(n_893),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_884),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_791),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_810),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_907),
.A2(n_762),
.B(n_702),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_792),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_810),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_789),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_799),
.B(n_702),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_871),
.A3(n_764),
.B(n_851),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_835),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_866),
.A2(n_871),
.A3(n_764),
.B(n_851),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_794),
.B(n_893),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_835),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1044),
.B(n_1037),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1033),
.B(n_955),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_921),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1047),
.B(n_996),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_977),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1035),
.B(n_1039),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1043),
.A2(n_1031),
.B1(n_1003),
.B2(n_1019),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_960),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_946),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_1038),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_988),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1051),
.B(n_933),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1046),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_931),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1048),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_924),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_1015),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_933),
.B(n_936),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_931),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_1011),
.B(n_998),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_934),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1015),
.B(n_983),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_939),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_956),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_946),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_924),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_1030),
.B(n_976),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_925),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_926),
.B(n_929),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_926),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_939),
.Y(n_1085)
);

INVxp33_ASAP7_75t_L g1086 ( 
.A(n_1018),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_983),
.B(n_981),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1030),
.B(n_1028),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1040),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_965),
.B(n_929),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1049),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1036),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1049),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1042),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1052),
.B(n_920),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1052),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1045),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_974),
.B(n_953),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_974),
.B(n_959),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_967),
.B(n_1013),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_964),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1048),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1014),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1050),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_1050),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_951),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_963),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_966),
.B(n_970),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_991),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1025),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_973),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_939),
.B(n_1034),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_972),
.B(n_980),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_944),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_994),
.B(n_1034),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_948),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_950),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_993),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_984),
.B(n_1008),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1034),
.B(n_1041),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_993),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_997),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1016),
.A2(n_1017),
.B(n_1027),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_972),
.B(n_980),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1020),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_997),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1006),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_969),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1026),
.B(n_987),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1020),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_987),
.B(n_935),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1024),
.A2(n_927),
.B(n_1021),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_938),
.B(n_985),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1006),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_928),
.Y(n_1135)
);

AO21x2_ASAP7_75t_L g1136 ( 
.A1(n_930),
.A2(n_940),
.B(n_999),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_923),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1023),
.A2(n_979),
.B(n_943),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_932),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_941),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_1029),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_971),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1000),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1005),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1009),
.B(n_989),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1022),
.B(n_1025),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1032),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_954),
.Y(n_1148)
);

INVx4_ASAP7_75t_L g1149 ( 
.A(n_1022),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_949),
.B(n_922),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_986),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1001),
.B(n_992),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_937),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_937),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_992),
.B(n_1012),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_957),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_937),
.Y(n_1157)
);

CKINVDCx14_ASAP7_75t_R g1158 ( 
.A(n_958),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_975),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_968),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1092),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1057),
.B(n_945),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1067),
.B(n_961),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1086),
.B(n_978),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1106),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1054),
.B(n_961),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1090),
.B(n_961),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1081),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1059),
.B(n_990),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1065),
.B(n_982),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1055),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1098),
.B(n_947),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1120),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_L g1174 ( 
.A(n_1150),
.B(n_952),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1106),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1092),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1088),
.B(n_942),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1094),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1076),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1067),
.B(n_962),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1095),
.B(n_968),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1076),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1060),
.A2(n_1007),
.B1(n_1002),
.B2(n_1010),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1075),
.B(n_1002),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1075),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1077),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1097),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1064),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1060),
.A2(n_995),
.B1(n_1004),
.B2(n_1158),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1074),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1099),
.B(n_1108),
.Y(n_1191)
);

AND2x4_ASAP7_75t_SL g1192 ( 
.A(n_1115),
.B(n_1081),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1061),
.B(n_1107),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1070),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1081),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1112),
.B(n_1061),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1086),
.B(n_1073),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1087),
.B(n_1133),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1115),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1111),
.B(n_1114),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1072),
.B(n_1083),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1123),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1156),
.B(n_1137),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1123),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1131),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1100),
.B(n_1072),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1053),
.B(n_1056),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1069),
.B(n_1079),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1080),
.B(n_1082),
.Y(n_1209)
);

INVx4_ASAP7_75t_R g1210 ( 
.A(n_1063),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1071),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1115),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1119),
.B(n_1085),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1084),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1058),
.B(n_1091),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1101),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1125),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1089),
.B(n_1145),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1131),
.B(n_1103),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1103),
.B(n_1113),
.Y(n_1223)
);

NOR2x1_ASAP7_75t_SL g1224 ( 
.A(n_1132),
.B(n_1142),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1113),
.B(n_1124),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1131),
.B(n_1124),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1062),
.B(n_1078),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1149),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1160),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1125),
.B(n_1062),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1078),
.B(n_1148),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1129),
.B(n_1063),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1130),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_L g1234 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1077),
.B(n_1128),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1128),
.B(n_1158),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1188),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1166),
.B(n_1146),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1191),
.B(n_1109),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1187),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1216),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1171),
.B(n_1134),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1165),
.B(n_1068),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1232),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1218),
.B(n_1118),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1197),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1212),
.B(n_1149),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1171),
.B(n_1121),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1205),
.B(n_1126),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1207),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1208),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1206),
.B(n_1122),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1180),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1181),
.B(n_1109),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1205),
.B(n_1147),
.Y(n_1256)
);

AND2x4_ASAP7_75t_SL g1257 ( 
.A(n_1185),
.B(n_1205),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1201),
.B(n_1193),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1175),
.B(n_1105),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1175),
.B(n_1105),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1186),
.B(n_1156),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1209),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1212),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1217),
.B(n_1141),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1161),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1188),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1176),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1177),
.B(n_1163),
.Y(n_1268)
);

INVxp67_ASAP7_75t_SL g1269 ( 
.A(n_1229),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1178),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1196),
.B(n_1141),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1228),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1163),
.B(n_1110),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1234),
.B(n_1066),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1214),
.B(n_1102),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1190),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1184),
.B(n_1104),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1203),
.B(n_1189),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1203),
.B(n_1151),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1200),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1202),
.B(n_1204),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1211),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1186),
.B(n_1159),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1264),
.B(n_1215),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1263),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1237),
.B(n_1266),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1242),
.Y(n_1287)
);

AOI21xp33_ASAP7_75t_L g1288 ( 
.A1(n_1278),
.A2(n_1174),
.B(n_1164),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1269),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1280),
.B(n_1220),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1256),
.B(n_1224),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1258),
.B(n_1173),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1256),
.B(n_1268),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1268),
.B(n_1238),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1243),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1282),
.B(n_1246),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1283),
.B(n_1162),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1279),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1241),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1238),
.B(n_1202),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1249),
.Y(n_1301)
);

NOR2x1_ASAP7_75t_L g1302 ( 
.A(n_1261),
.B(n_1236),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1257),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1255),
.B(n_1204),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1255),
.B(n_1164),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1278),
.B(n_1168),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1246),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1272),
.Y(n_1308)
);

AND3x2_ASAP7_75t_L g1309 ( 
.A(n_1247),
.B(n_1199),
.C(n_1198),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1279),
.B(n_1189),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1271),
.B(n_1233),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1240),
.B(n_1194),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1265),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1267),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1253),
.B(n_1194),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1270),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1276),
.Y(n_1317)
);

NAND2x1_ASAP7_75t_L g1318 ( 
.A(n_1272),
.B(n_1210),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1287),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1297),
.B(n_1248),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1294),
.B(n_1293),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1295),
.B(n_1251),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1289),
.B(n_1285),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1311),
.B(n_1233),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1300),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1299),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1286),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1294),
.B(n_1311),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1310),
.A2(n_1157),
.B1(n_1154),
.B2(n_1153),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1293),
.B(n_1259),
.Y(n_1331)
);

CKINVDCx16_ASAP7_75t_R g1332 ( 
.A(n_1293),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1300),
.B(n_1259),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1305),
.B(n_1260),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1305),
.B(n_1252),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1290),
.A2(n_1221),
.B(n_1235),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_R g1337 ( 
.A(n_1309),
.B(n_1281),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1291),
.B(n_1260),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1313),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1284),
.B(n_1244),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1292),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1312),
.B(n_1262),
.Y(n_1342)
);

AOI322xp5_ASAP7_75t_L g1343 ( 
.A1(n_1310),
.A2(n_1239),
.A3(n_1183),
.B1(n_1253),
.B2(n_1245),
.C1(n_1275),
.C2(n_1273),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1326),
.B(n_1307),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1319),
.Y(n_1345)
);

OA21x2_ASAP7_75t_SL g1346 ( 
.A1(n_1341),
.A2(n_1315),
.B(n_1291),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1327),
.Y(n_1347)
);

AOI322xp5_ASAP7_75t_L g1348 ( 
.A1(n_1320),
.A2(n_1288),
.A3(n_1302),
.B1(n_1239),
.B2(n_1183),
.C1(n_1304),
.C2(n_1301),
.Y(n_1348)
);

OAI32xp33_ASAP7_75t_L g1349 ( 
.A1(n_1337),
.A2(n_1332),
.A3(n_1326),
.B1(n_1329),
.B2(n_1306),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1337),
.A2(n_1320),
.B1(n_1330),
.B2(n_1342),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1339),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1324),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1328),
.A2(n_1306),
.B1(n_1318),
.B2(n_1298),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1330),
.A2(n_1273),
.B1(n_1275),
.B2(n_1277),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1335),
.A2(n_1317),
.B1(n_1316),
.B2(n_1314),
.C(n_1169),
.Y(n_1355)
);

OAI211xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1323),
.A2(n_1308),
.B(n_1231),
.C(n_1227),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1325),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1334),
.B(n_1308),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1338),
.A2(n_1291),
.B1(n_1277),
.B2(n_1250),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1336),
.A2(n_1298),
.B1(n_1303),
.B2(n_1225),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1340),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1350),
.B(n_1325),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1349),
.A2(n_1338),
.B(n_1322),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1304),
.B2(n_1170),
.C(n_1172),
.Y(n_1364)
);

AOI211xp5_ASAP7_75t_L g1365 ( 
.A1(n_1360),
.A2(n_1331),
.B(n_1281),
.C(n_1321),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1351),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1345),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1347),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1364),
.A2(n_1356),
.B1(n_1352),
.B2(n_1346),
.C(n_1354),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1367),
.B(n_1357),
.Y(n_1370)
);

NOR3xp33_ASAP7_75t_SL g1371 ( 
.A(n_1362),
.B(n_1353),
.C(n_1358),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1368),
.B(n_1366),
.Y(n_1372)
);

OAI21xp33_ASAP7_75t_L g1373 ( 
.A1(n_1365),
.A2(n_1348),
.B(n_1361),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1370),
.B(n_1363),
.C(n_1353),
.D(n_1343),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1371),
.B(n_1359),
.C(n_1344),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1372),
.Y(n_1376)
);

OAI211xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1373),
.A2(n_1223),
.B(n_1138),
.C(n_1152),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1213),
.Y(n_1378)
);

NAND4xp25_ASAP7_75t_L g1379 ( 
.A(n_1370),
.B(n_1230),
.C(n_1298),
.D(n_1195),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1376),
.Y(n_1380)
);

NOR4xp25_ASAP7_75t_L g1381 ( 
.A(n_1377),
.B(n_1179),
.C(n_1219),
.D(n_1182),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1378),
.B(n_1213),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1381),
.B(n_1374),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_L g1384 ( 
.A(n_1380),
.B(n_1375),
.C(n_1379),
.D(n_1222),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1383),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1385),
.B(n_1384),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1386),
.Y(n_1387)
);

AOI22x1_ASAP7_75t_L g1388 ( 
.A1(n_1386),
.A2(n_1385),
.B1(n_1382),
.B2(n_1182),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1387),
.A2(n_1155),
.B(n_1226),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1388),
.A2(n_1136),
.B1(n_1250),
.B2(n_1274),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1390),
.B(n_1254),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1389),
.B(n_1254),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1392),
.B(n_1192),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1393),
.A2(n_1391),
.B1(n_1136),
.B2(n_1135),
.Y(n_1394)
);


endmodule