module fake_jpeg_415_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_54),
.B1(n_51),
.B2(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_43),
.B1(n_48),
.B2(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_76),
.B1(n_64),
.B2(n_53),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_50),
.B1(n_53),
.B2(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_55),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_52),
.B1(n_62),
.B2(n_49),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_91),
.B1(n_79),
.B2(n_5),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_6),
.B(n_7),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_11),
.B(n_14),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_7),
.B(n_8),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_39),
.B(n_17),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_31),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_120),
.C(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_123),
.B1(n_107),
.B2(n_35),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_23),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_108),
.Y(n_129)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_24),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_26),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_134),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_37),
.B1(n_32),
.B2(n_36),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_113),
.B(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_141),
.B(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_124),
.B1(n_123),
.B2(n_111),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_143),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_142),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_146),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_124),
.B1(n_138),
.B2(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_148),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_132),
.B1(n_130),
.B2(n_129),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_132),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_117),
.Y(n_155)
);


endmodule