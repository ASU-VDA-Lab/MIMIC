module fake_jpeg_30496_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B(n_4),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_46),
.B1(n_39),
.B2(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_46),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_44),
.B(n_42),
.C(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

AO21x2_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_8),
.B(n_12),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_76),
.B1(n_81),
.B2(n_25),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_36),
.B1(n_20),
.B2(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_64),
.B1(n_58),
.B2(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_7),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_90),
.B(n_84),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_16),
.B(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_24),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_26),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.Y(n_108)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.C(n_95),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_90),
.B(n_92),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_84),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_96),
.B1(n_100),
.B2(n_97),
.C(n_93),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_95),
.C(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_108),
.C(n_88),
.Y(n_111)
);

AOI31xp67_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_110),
.A3(n_99),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_85),
.B1(n_29),
.B2(n_30),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_27),
.Y(n_115)
);


endmodule