module fake_jpeg_25263_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_17),
.B1(n_30),
.B2(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_17),
.B1(n_18),
.B2(n_15),
.Y(n_72)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_36),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_19),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_61),
.Y(n_92)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_16),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_18),
.B(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_78),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_33),
.B1(n_30),
.B2(n_17),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_36),
.B1(n_34),
.B2(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_63),
.B1(n_76),
.B2(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_77),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_29),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_36),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_87),
.B1(n_89),
.B2(n_98),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_14),
.C(n_12),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_15),
.B1(n_21),
.B2(n_36),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_34),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_90),
.B(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_21),
.B1(n_34),
.B2(n_22),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_20),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_45),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_73),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_87),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_106),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_109),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_70),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_112),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_70),
.B(n_20),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_121),
.Y(n_134)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_120),
.Y(n_123)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_60),
.B(n_67),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_118),
.B(n_101),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_0),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_89),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_110),
.C(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_132),
.C(n_105),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_81),
.B(n_88),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_133),
.B(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_99),
.C(n_88),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_81),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_81),
.B1(n_98),
.B2(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_138),
.B1(n_140),
.B2(n_114),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_100),
.B1(n_85),
.B2(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_84),
.B1(n_59),
.B2(n_82),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_120),
.C(n_115),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_152),
.C(n_127),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_109),
.B(n_118),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_107),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_153),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_46),
.Y(n_151)
);

XOR2x1_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_154),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_116),
.C(n_60),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_137),
.B1(n_136),
.B2(n_129),
.Y(n_153)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_123),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_161),
.C(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_134),
.C(n_139),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_165),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_125),
.C(n_129),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_124),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_175),
.B1(n_167),
.B2(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_174),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_153),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_156),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_126),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_180),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_151),
.B1(n_167),
.B2(n_142),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_182),
.C(n_141),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_141),
.B1(n_159),
.B2(n_60),
.Y(n_182)
);

AOI211xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_172),
.B(n_159),
.C(n_126),
.Y(n_185)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_186),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_2),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_182),
.B1(n_180),
.B2(n_4),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_190),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_5),
.C(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_7),
.B(n_8),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_196),
.Y(n_199)
);


endmodule