module fake_jpeg_1129_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_0),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_19),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_40),
.B1(n_44),
.B2(n_38),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_62),
.B1(n_57),
.B2(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_56),
.Y(n_76)
);

XNOR2x2_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_54),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_39),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_47),
.B1(n_37),
.B2(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_62),
.B1(n_47),
.B2(n_37),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_73),
.B1(n_21),
.B2(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_39),
.B1(n_73),
.B2(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_93),
.C(n_7),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_17),
.B(n_32),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_100),
.B1(n_16),
.B2(n_29),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_9),
.Y(n_113)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_8),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_106),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_13),
.B(n_28),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_6),
.B(n_7),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

AO221x1_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_94),
.B1(n_98),
.B2(n_26),
.C(n_27),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_90),
.C(n_95),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_107),
.C(n_108),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_121),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_102),
.B(n_24),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_119),
.B1(n_116),
.B2(n_115),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_11),
.C(n_34),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_123),
.Y(n_129)
);


endmodule