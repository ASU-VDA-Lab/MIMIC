module fake_jpeg_28622_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_0),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx2_ASAP7_75t_SL g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_50),
.B1(n_63),
.B2(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_81),
.B1(n_85),
.B2(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_91),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_50),
.B1(n_63),
.B2(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_77),
.B1(n_58),
.B2(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_69),
.B1(n_52),
.B2(n_65),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_64),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_108),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_1),
.B(n_2),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_113),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_61),
.B1(n_60),
.B2(n_59),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_3),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_122),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_7),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_28),
.A3(n_48),
.B1(n_43),
.B2(n_40),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_119),
.B1(n_133),
.B2(n_120),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_27),
.C(n_39),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_31),
.C(n_13),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_142),
.B1(n_150),
.B2(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_12),
.B1(n_14),
.B2(n_18),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_148),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_21),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_25),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_152),
.B1(n_135),
.B2(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_135),
.B1(n_121),
.B2(n_38),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_37),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_164),
.C(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_151),
.C(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_153),
.B1(n_136),
.B2(n_158),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_163),
.B(n_156),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_161),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_157),
.Y(n_173)
);


endmodule