module fake_jpeg_700_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_28),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_31),
.C(n_26),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.C(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_31),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_30),
.B2(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_37),
.B1(n_15),
.B2(n_16),
.Y(n_59)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_44),
.B(n_5),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_7),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_62),
.B(n_10),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_75),
.B(n_68),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_8),
.CI(n_11),
.CON(n_75),
.SN(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_71),
.B(n_72),
.Y(n_78)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_76),
.B(n_75),
.C(n_70),
.D(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_17),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_19),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_23),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_24),
.Y(n_83)
);


endmodule