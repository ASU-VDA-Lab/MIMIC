module fake_jpeg_30933_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

AOI22xp33_ASAP7_75t_L g5 ( 
.A1(n_0),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_5)
);

INVx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g7 ( 
.A1(n_5),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_7),
.A2(n_8),
.B(n_1),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_SL g8 ( 
.A1(n_5),
.A2(n_0),
.B(n_1),
.Y(n_8)
);

NOR3xp33_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_10),
.C(n_6),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_6),
.B(n_3),
.Y(n_10)
);


endmodule