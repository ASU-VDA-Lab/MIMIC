module fake_jpeg_8851_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

OA22x2_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_23),
.B1(n_29),
.B2(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_16),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_34),
.B1(n_31),
.B2(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_27),
.B(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_41),
.B1(n_24),
.B2(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_27),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_24),
.B1(n_33),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_24),
.B1(n_33),
.B2(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_83),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_88),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_17),
.B(n_20),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_19),
.C(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_106),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_60),
.B1(n_45),
.B2(n_52),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_108),
.B1(n_111),
.B2(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_100),
.B(n_105),
.Y(n_149)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_116),
.B(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_112),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_45),
.B1(n_20),
.B2(n_22),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_66),
.A2(n_75),
.B1(n_93),
.B2(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_119),
.B1(n_106),
.B2(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_17),
.B(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_28),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_71),
.B1(n_55),
.B2(n_48),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_141),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_130),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_82),
.B(n_76),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g176 ( 
.A(n_125),
.B(n_145),
.C(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_93),
.C(n_83),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_139),
.C(n_61),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_129),
.B1(n_150),
.B2(n_96),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_72),
.B1(n_74),
.B2(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_135),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_84),
.B1(n_85),
.B2(n_92),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_142),
.B1(n_119),
.B2(n_112),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_85),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_94),
.A2(n_71),
.B1(n_77),
.B2(n_56),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_120),
.B1(n_96),
.B2(n_87),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_73),
.B(n_17),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_89),
.B1(n_53),
.B2(n_67),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_28),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_114),
.Y(n_154)
);

OR2x4_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_19),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_115),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_89),
.B1(n_71),
.B2(n_19),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_154),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_168),
.B(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_21),
.Y(n_193)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_173),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_117),
.B(n_104),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_167),
.B(n_181),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_172),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_109),
.B(n_96),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_141),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_128),
.B1(n_121),
.B2(n_139),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_136),
.B1(n_132),
.B2(n_129),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_17),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_17),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_9),
.C(n_15),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_17),
.B(n_30),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_19),
.B(n_30),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_16),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_185),
.A2(n_191),
.B1(n_195),
.B2(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_121),
.B1(n_134),
.B2(n_144),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_134),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_199),
.C(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_21),
.B1(n_30),
.B2(n_87),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_154),
.B1(n_159),
.B2(n_176),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_9),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_156),
.B1(n_175),
.B2(n_170),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_16),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_181),
.C(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_159),
.B1(n_163),
.B2(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_193),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_220),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_230),
.C(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_152),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_165),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_232),
.B(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_162),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_227),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_198),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_186),
.B(n_168),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_203),
.B(n_196),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_198),
.B1(n_188),
.B2(n_186),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_253),
.B1(n_227),
.B2(n_214),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_242),
.B(n_254),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_188),
.B(n_187),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_202),
.C(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_252),
.C(n_230),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_200),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_182),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_163),
.C(n_4),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_14),
.B(n_12),
.Y(n_254)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_268),
.C(n_269),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_213),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_262),
.B(n_263),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_223),
.B1(n_212),
.B2(n_210),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_264),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_231),
.B1(n_252),
.B2(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_224),
.B1(n_210),
.B2(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_237),
.B(n_254),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_222),
.C(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_220),
.C(n_216),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_240),
.B(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_265),
.B1(n_257),
.B2(n_5),
.Y(n_291)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_241),
.B1(n_242),
.B2(n_239),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_269),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_250),
.B1(n_246),
.B2(n_238),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_245),
.B(n_11),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.C(n_281),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_10),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_286),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_271),
.C(n_5),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_265),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_3),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_272),
.B1(n_291),
.B2(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_296),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_271),
.B(n_281),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_285),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

AOI321xp33_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_6),
.A3(n_7),
.B1(n_294),
.B2(n_297),
.C(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_307),
.C(n_303),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_299),
.A2(n_289),
.B(n_288),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_309),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_308),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_313),
.Y(n_314)
);


endmodule