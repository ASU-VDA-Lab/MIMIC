module real_jpeg_26470_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_249;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_216;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_7),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_4),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_4),
.A2(n_41),
.B1(n_70),
.B2(n_71),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_26),
.C(n_29),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_27),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_48),
.C(n_51),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_4),
.B(n_67),
.C(n_70),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_4),
.B(n_100),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_4),
.B(n_60),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_19),
.B1(n_20),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_189)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_32),
.B1(n_70),
.B2(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_21),
.B1(n_51),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_21),
.B1(n_70),
.B2(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_75),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_73),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_35),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_35),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_38),
.B(n_39),
.Y(n_37)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_22),
.A2(n_27),
.B1(n_40),
.B2(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_24),
.B(n_185),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_29),
.B(n_219),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_36),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_36),
.B(n_289),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_42),
.CI(n_53),
.CON(n_36),
.SN(n_36)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_38),
.A2(n_39),
.B(n_56),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_45),
.A2(n_50),
.B(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_60),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_46),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_50),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_50),
.A2(n_104),
.B(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_51),
.B(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.C(n_61),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_54),
.B(n_123),
.C(n_130),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_54),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_54),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_54),
.A2(n_130),
.B1(n_131),
.B2(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_54),
.A2(n_102),
.B1(n_144),
.B2(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_54),
.B(n_102),
.C(n_182),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_61),
.B1(n_112),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_58),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_108),
.C(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_63),
.B(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_65),
.A2(n_90),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_69),
.A2(n_89),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_70),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_288),
.B(n_290),
.Y(n_75)
);

OAI211xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_132),
.B(n_146),
.C(n_287),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_117),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_117),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_95),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_97),
.C(n_106),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_91),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_91),
.B1(n_92),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_80),
.A2(n_87),
.B1(n_120),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_82),
.B(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_85),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_83),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_84),
.A2(n_125),
.B(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_87),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_107),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_98),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_102),
.B(n_203),
.C(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_102),
.A2(n_193),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_109),
.B1(n_140),
.B2(n_145),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_130),
.C(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_108),
.A2(n_109),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_108),
.A2(n_109),
.B1(n_164),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_156),
.C(n_164),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_109),
.B(n_136),
.C(n_140),
.Y(n_289)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_121),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_124),
.Y(n_278)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_127),
.A2(n_128),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_127),
.A2(n_128),
.B1(n_216),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_128),
.B(n_210),
.C(n_216),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_128),
.B(n_187),
.C(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_130),
.A2(n_131),
.B1(n_178),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_130),
.A2(n_131),
.B1(n_162),
.B2(n_175),
.Y(n_255)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_131),
.B(n_162),
.C(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_147),
.C(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_134),
.B(n_135),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_168),
.B(n_286),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_166),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_150),
.B(n_166),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_151),
.B(n_153),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_155),
.B(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_156),
.A2(n_157),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_162),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_189),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_162),
.A2(n_175),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_281),
.B(n_285),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_206),
.B(n_267),
.C(n_280),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_195),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_171),
.B(n_195),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_181),
.B2(n_194),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_180),
.C(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_186),
.A2(n_187),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_241),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_197),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_205),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_266),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_225),
.B(n_265),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_209),
.B(n_222),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_210),
.A2(n_211),
.B1(n_261),
.B2(n_263),
.Y(n_260)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_258),
.B(n_264),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_252),
.B(n_257),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_244),
.B(n_251),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_234),
.B(n_243),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_242),
.Y(n_234)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_277),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);


endmodule