module fake_netlist_6_3193_n_8072 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_8072);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_8072;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_6566;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_6872;
wire n_1351;
wire n_5254;
wire n_6441;
wire n_1212;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_7111;
wire n_6141;
wire n_3849;
wire n_7933;
wire n_7967;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_6960;
wire n_1061;
wire n_3089;
wire n_783;
wire n_7180;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_7190;
wire n_7504;
wire n_6126;
wire n_6725;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_8023;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_2179;
wire n_5963;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_4249;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_6999;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_7161;
wire n_3030;
wire n_830;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_7000;
wire n_7398;
wire n_2926;
wire n_1078;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_6882;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_6325;
wire n_4724;
wire n_945;
wire n_5598;
wire n_7983;
wire n_7389;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_8070;
wire n_4696;
wire n_6660;
wire n_4347;
wire n_5259;
wire n_6913;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_8022;
wire n_5930;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_7686;
wire n_1421;
wire n_3664;
wire n_6914;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_6374;
wire n_2843;
wire n_7651;
wire n_6628;
wire n_3760;
wire n_6015;
wire n_4262;
wire n_1560;
wire n_734;
wire n_1088;
wire n_6526;
wire n_1894;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_7196;
wire n_3347;
wire n_5136;
wire n_907;
wire n_8040;
wire n_5638;
wire n_4110;
wire n_6784;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_6323;
wire n_6110;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_6371;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_7256;
wire n_6404;
wire n_7331;
wire n_7774;
wire n_7856;
wire n_5680;
wire n_6674;
wire n_6148;
wire n_6951;
wire n_7625;
wire n_4102;
wire n_3871;
wire n_1641;
wire n_2735;
wire n_4662;
wire n_6989;
wire n_4671;
wire n_7863;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_6896;
wire n_7770;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_7147;
wire n_2770;
wire n_4507;
wire n_2101;
wire n_5902;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_6196;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_6485;
wire n_6107;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_1075;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_7564;
wire n_3859;
wire n_2692;
wire n_6768;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_7110;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_6431;
wire n_6990;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_7849;
wire n_4331;
wire n_7297;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_7533;
wire n_7221;
wire n_4375;
wire n_1701;
wire n_6575;
wire n_6055;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_5897;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_7569;
wire n_2641;
wire n_7734;
wire n_7062;
wire n_7823;
wire n_7861;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_7039;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_7077;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_5865;
wire n_6836;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_7905;
wire n_2092;
wire n_7753;
wire n_1654;
wire n_6771;
wire n_7950;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_6248;
wire n_6952;
wire n_6795;
wire n_5314;
wire n_1588;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_3968;
wire n_2096;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_5795;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_5226;
wire n_6715;
wire n_6714;
wire n_890;
wire n_7677;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_6584;
wire n_1709;
wire n_7009;
wire n_2393;
wire n_2657;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_6581;
wire n_2279;
wire n_6010;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_7013;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_7290;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_7488;
wire n_2558;
wire n_7315;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_6042;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_7438;
wire n_2145;
wire n_7268;
wire n_7337;
wire n_898;
wire n_4964;
wire n_5957;
wire n_6965;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_925;
wire n_1932;
wire n_1101;
wire n_6800;
wire n_4636;
wire n_7461;
wire n_4322;
wire n_3644;
wire n_6955;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_7278;
wire n_6509;
wire n_4576;
wire n_7454;
wire n_5929;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_6839;
wire n_7232;
wire n_4345;
wire n_7377;
wire n_996;
wire n_6646;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_7098;
wire n_7069;
wire n_7904;
wire n_6033;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_6097;
wire n_6369;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_3700;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_3104;
wire n_6809;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_7840;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_1432;
wire n_5212;
wire n_989;
wire n_7080;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_5811;
wire n_899;
wire n_7739;
wire n_6766;
wire n_1035;
wire n_4914;
wire n_7624;
wire n_4939;
wire n_7629;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_7003;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_5901;
wire n_6538;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_7010;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_6519;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_6530;
wire n_7219;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_7299;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_6402;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_7243;
wire n_6609;
wire n_7326;
wire n_5326;
wire n_7471;
wire n_7067;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_6748;
wire n_7741;
wire n_998;
wire n_5035;
wire n_717;
wire n_7790;
wire n_6149;
wire n_1383;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_1424;
wire n_6414;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_7528;
wire n_8026;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_7941;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_6902;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_5741;
wire n_2773;
wire n_6205;
wire n_6380;
wire n_7478;
wire n_7913;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_7939;
wire n_2788;
wire n_964;
wire n_4756;
wire n_6449;
wire n_2797;
wire n_6723;
wire n_7458;
wire n_6440;
wire n_7436;
wire n_4746;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_7435;
wire n_3441;
wire n_3534;
wire n_6997;
wire n_5952;
wire n_3964;
wire n_2416;
wire n_5947;
wire n_1877;
wire n_3944;
wire n_6124;
wire n_6736;
wire n_7685;
wire n_7363;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_5985;
wire n_2209;
wire n_3605;
wire n_6622;
wire n_1602;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_6528;
wire n_2274;
wire n_7532;
wire n_8051;
wire n_5761;
wire n_6773;
wire n_4618;
wire n_7375;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_6885;
wire n_2146;
wire n_6531;
wire n_2131;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_7912;
wire n_2575;
wire n_5100;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_7728;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_6339;
wire n_1917;
wire n_8024;
wire n_1580;
wire n_7730;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_7281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_7711;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_6763;
wire n_2049;
wire n_858;
wire n_5182;
wire n_7858;
wire n_956;
wire n_5534;
wire n_8003;
wire n_4880;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_3845;
wire n_1696;
wire n_6556;
wire n_1594;
wire n_1869;
wire n_6889;
wire n_7230;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_5196;
wire n_6199;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_6726;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_7011;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_2448;
wire n_5949;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_6478;
wire n_7952;
wire n_3406;
wire n_820;
wire n_951;
wire n_6100;
wire n_6516;
wire n_952;
wire n_3919;
wire n_6977;
wire n_7660;
wire n_6915;
wire n_2263;
wire n_7834;
wire n_5185;
wire n_6911;
wire n_6599;
wire n_974;
wire n_6522;
wire n_5023;
wire n_2656;
wire n_4952;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_7890;
wire n_3973;
wire n_2756;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_807;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_1275;
wire n_2884;
wire n_6808;
wire n_1510;
wire n_7620;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_6207;
wire n_6931;
wire n_7006;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_6963;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_7381;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_7837;
wire n_7717;
wire n_1037;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_7627;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_3195;
wire n_2526;
wire n_6346;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_7335;
wire n_4189;
wire n_3817;
wire n_7811;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_6059;
wire n_7499;
wire n_3042;
wire n_6065;
wire n_7292;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_6075;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_7977;
wire n_7211;
wire n_5618;
wire n_6861;
wire n_6781;
wire n_1586;
wire n_7847;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_6133;
wire n_3723;
wire n_1190;
wire n_7822;
wire n_6453;
wire n_4380;
wire n_5978;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_6127;
wire n_4398;
wire n_2498;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_7289;
wire n_4193;
wire n_3570;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_7354;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_7960;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_7482;
wire n_1043;
wire n_4090;
wire n_6115;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_6838;
wire n_6867;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_6139;
wire n_1361;
wire n_6256;
wire n_7965;
wire n_3262;
wire n_6613;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_6361;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_6085;
wire n_7474;
wire n_5731;
wire n_6329;
wire n_6678;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_7325;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_6370;
wire n_2518;
wire n_5883;
wire n_7166;
wire n_6554;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_3988;
wire n_6560;
wire n_1720;
wire n_3476;
wire n_7028;
wire n_4842;
wire n_7838;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_7873;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_6535;
wire n_942;
wire n_7518;
wire n_2798;
wire n_7414;
wire n_6147;
wire n_2852;
wire n_1524;
wire n_6448;
wire n_7791;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_3292;
wire n_1496;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_6643;
wire n_7146;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_6157;
wire n_4859;
wire n_2626;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_5218;
wire n_7052;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_5960;
wire n_4571;
wire n_3698;
wire n_7888;
wire n_5358;
wire n_6397;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_6073;
wire n_7502;
wire n_1484;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_7312;
wire n_7919;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_7085;
wire n_1373;
wire n_3958;
wire n_6939;
wire n_7848;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_6689;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_1385;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_7288;
wire n_1257;
wire n_7707;
wire n_3197;
wire n_7223;
wire n_7833;
wire n_4987;
wire n_5512;
wire n_7274;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_6206;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_3124;
wire n_1741;
wire n_7466;
wire n_1002;
wire n_6529;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_6290;
wire n_7429;
wire n_6025;
wire n_1337;
wire n_1477;
wire n_7277;
wire n_6455;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_7179;
wire n_7122;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_4376;
wire n_6203;
wire n_1001;
wire n_6408;
wire n_2241;
wire n_6555;
wire n_7683;
wire n_6150;
wire n_7630;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_6892;
wire n_4462;
wire n_7061;
wire n_6401;
wire n_7322;
wire n_1716;
wire n_6685;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_7051;
wire n_1976;
wire n_7880;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_6679;
wire n_749;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_6574;
wire n_6571;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_7824;
wire n_1074;
wire n_3569;
wire n_739;
wire n_7094;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8060;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_7036;
wire n_6392;
wire n_1810;
wire n_5915;
wire n_7351;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_7608;
wire n_5779;
wire n_2020;
wire n_1643;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_7909;
wire n_7413;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_6286;
wire n_7675;
wire n_4023;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_721;
wire n_1461;
wire n_742;
wire n_7175;
wire n_3617;
wire n_2076;
wire n_6019;
wire n_3567;
wire n_1598;
wire n_7524;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_6214;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_7783;
wire n_6692;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_6036;
wire n_4391;
wire n_946;
wire n_1303;
wire n_6552;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_7697;
wire n_1944;
wire n_6403;
wire n_7306;
wire n_1347;
wire n_7947;
wire n_795;
wire n_1221;
wire n_7547;
wire n_7470;
wire n_6013;
wire n_7733;
wire n_1245;
wire n_7693;
wire n_3215;
wire n_6491;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_6348;
wire n_6744;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_6982;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_6293;
wire n_6661;
wire n_5847;
wire n_7345;
wire n_6049;
wire n_1460;
wire n_911;
wire n_7385;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_6558;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_6136;
wire n_1058;
wire n_3378;
wire n_6855;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_6312;
wire n_2505;
wire n_4817;
wire n_6668;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_7653;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_6859;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_6388;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_6995;
wire n_4491;
wire n_5696;
wire n_7032;
wire n_4486;
wire n_6971;
wire n_1816;
wire n_6131;
wire n_5848;
wire n_3024;
wire n_7475;
wire n_4612;
wire n_6435;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_8018;
wire n_3936;
wire n_1349;
wire n_7937;
wire n_6829;
wire n_2723;
wire n_5485;
wire n_7819;
wire n_5823;
wire n_7305;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_7993;
wire n_7181;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_6822;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_7071;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_7391;
wire n_6617;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_7511;
wire n_6533;
wire n_849;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_1753;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_2471;
wire n_6983;
wire n_4412;
wire n_2807;
wire n_6801;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_6113;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_7321;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_3815;
wire n_3896;
wire n_6655;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_7584;
wire n_4457;
wire n_7537;
wire n_4093;
wire n_1616;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_6837;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_7486;
wire n_6756;
wire n_1027;
wire n_3266;
wire n_7023;
wire n_3574;
wire n_7496;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_7410;
wire n_6200;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_6670;
wire n_3741;
wire n_6373;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_7899;
wire n_4819;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_1708;
wire n_7131;
wire n_805;
wire n_6411;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_7302;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_7797;
wire n_3668;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_7582;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_6534;
wire n_3340;
wire n_5227;
wire n_7809;
wire n_873;
wire n_3946;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_7060;
wire n_7607;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_7867;
wire n_3275;
wire n_836;
wire n_6135;
wire n_7761;
wire n_8007;
wire n_3678;
wire n_6814;
wire n_3440;
wire n_8001;
wire n_2094;
wire n_7525;
wire n_1511;
wire n_7257;
wire n_2356;
wire n_7553;
wire n_1422;
wire n_7529;
wire n_1772;
wire n_4692;
wire n_6791;
wire n_3165;
wire n_1119;
wire n_6824;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_7650;
wire n_3316;
wire n_6903;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_6450;
wire n_3261;
wire n_7520;
wire n_4187;
wire n_6309;
wire n_940;
wire n_7903;
wire n_2058;
wire n_2660;
wire n_6733;
wire n_7384;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_3532;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_7639;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_6179;
wire n_6395;
wire n_976;
wire n_7054;
wire n_7605;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_7433;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_808;
wire n_5519;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_6654;
wire n_8019;
wire n_3791;
wire n_6083;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_4320;
wire n_7832;
wire n_3884;
wire n_5808;
wire n_7726;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_6120;
wire n_6068;
wire n_6933;
wire n_4141;
wire n_3438;
wire n_6547;
wire n_5193;
wire n_6423;
wire n_2850;
wire n_6342;
wire n_6641;
wire n_1481;
wire n_6984;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_7441;
wire n_7106;
wire n_7213;
wire n_3883;
wire n_5961;
wire n_5866;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_6687;
wire n_5822;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_7031;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_788;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_7133;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_1866;
wire n_7424;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_7523;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_6790;
wire n_5953;
wire n_3099;
wire n_7141;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6505;
wire n_1663;
wire n_6459;
wire n_4172;
wire n_3403;
wire n_7626;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_3686;
wire n_7669;
wire n_4502;
wire n_5958;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_7367;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_7323;
wire n_7189;
wire n_7301;
wire n_6258;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_6905;
wire n_3725;
wire n_6704;
wire n_3933;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_1175;
wire n_7244;
wire n_7368;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_903;
wire n_7633;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_8063;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_816;
wire n_6210;
wire n_6500;
wire n_8032;
wire n_1188;
wire n_7427;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_6163;
wire n_7628;
wire n_5972;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_1624;
wire n_1124;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_8039;
wire n_5757;
wire n_1515;
wire n_961;
wire n_7557;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_7128;
wire n_2377;
wire n_6849;
wire n_7594;
wire n_950;
wire n_7457;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_7788;
wire n_4361;
wire n_5488;
wire n_6760;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_7752;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_6825;
wire n_1987;
wire n_7586;
wire n_6452;
wire n_968;
wire n_7767;
wire n_2271;
wire n_1008;
wire n_6611;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_7207;
wire n_5843;
wire n_7744;
wire n_2078;
wire n_7021;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_7748;
wire n_3450;
wire n_6827;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_6227;
wire n_7215;
wire n_7485;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_5523;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_8016;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_6564;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_6468;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_6857;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_3293;
wire n_872;
wire n_3922;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_847;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_6871;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_6904;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_7017;
wire n_7777;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_7652;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_6499;
wire n_7830;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_7138;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_7966;
wire n_5059;
wire n_5887;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_6276;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_7208;
wire n_2119;
wire n_947;
wire n_1117;
wire n_7961;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_6893;
wire n_7406;
wire n_3223;
wire n_3140;
wire n_7807;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_7680;
wire n_926;
wire n_3654;
wire n_2848;
wire n_1849;
wire n_919;
wire n_1698;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_5937;
wire n_777;
wire n_6422;
wire n_1299;
wire n_6751;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_6040;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_4659;
wire n_3600;
wire n_6741;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_3324;
wire n_2338;
wire n_1178;
wire n_6160;
wire n_6650;
wire n_7066;
wire n_7183;
wire n_796;
wire n_1195;
wire n_7789;
wire n_7606;
wire n_6192;
wire n_1811;
wire n_6368;
wire n_7140;
wire n_7193;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_5721;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_6012;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_7344;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_6707;
wire n_4874;
wire n_4401;
wire n_889;
wire n_6064;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_6787;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_7710;
wire n_2389;
wire n_7892;
wire n_2132;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_1787;
wire n_6769;
wire n_1993;
wire n_2281;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_7206;
wire n_4223;
wire n_7538;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_6799;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_7716;
wire n_6487;
wire n_5121;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_6807;
wire n_7251;
wire n_4489;
wire n_4839;
wire n_7254;
wire n_2596;
wire n_3163;
wire n_7540;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_6563;
wire n_1531;
wire n_7882;
wire n_2828;
wire n_7554;
wire n_2384;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_6341;
wire n_6384;
wire n_1901;
wire n_3869;
wire n_7421;
wire n_2556;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_7991;
wire n_6233;
wire n_2227;
wire n_6377;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_6257;
wire n_2159;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_4955;
wire n_4149;
wire n_5936;
wire n_4355;
wire n_7646;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_6587;
wire n_1129;
wire n_6987;
wire n_7781;
wire n_7360;
wire n_2181;
wire n_6069;
wire n_2911;
wire n_7497;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_7665;
wire n_3429;
wire n_2379;
wire n_7793;
wire n_3554;
wire n_1593;
wire n_6991;
wire n_1202;
wire n_7101;
wire n_7671;
wire n_1635;
wire n_7530;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_7204;
wire n_6887;
wire n_7578;
wire n_3462;
wire n_7654;
wire n_2851;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_8059;
wire n_6633;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_6579;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_5875;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_732;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_7120;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_6789;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_6252;
wire n_1871;
wire n_4860;
wire n_6211;
wire n_845;
wire n_5844;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_6164;
wire n_768;
wire n_7576;
wire n_6173;
wire n_7786;
wire n_3651;
wire n_7313;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_6934;
wire n_6630;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_6737;
wire n_4488;
wire n_3767;
wire n_6612;
wire n_6606;
wire n_2544;
wire n_6695;
wire n_3550;
wire n_4211;
wire n_7779;
wire n_6189;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_750;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_3839;
wire n_2823;
wire n_6410;
wire n_6158;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_1057;
wire n_7419;
wire n_6506;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_6935;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_6688;
wire n_5980;
wire n_7818;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_6608;
wire n_3533;
wire n_1622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_6798;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_6753;
wire n_2171;
wire n_6527;
wire n_7341;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_6639;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_6430;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_7996;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_7517;
wire n_1152;
wire n_6627;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_6058;
wire n_711;
wire n_7745;
wire n_3105;
wire n_2872;
wire n_6666;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_6190;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_6249;
wire n_2738;
wire n_972;
wire n_5348;
wire n_6594;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_7095;
wire n_936;
wire n_3821;
wire n_3045;
wire n_6969;
wire n_885;
wire n_6615;
wire n_6161;
wire n_7459;
wire n_2970;
wire n_2167;
wire n_7294;
wire n_2342;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_7184;
wire n_6607;
wire n_6062;
wire n_7908;
wire n_1974;
wire n_4122;
wire n_7974;
wire n_7551;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_6482;
wire n_4128;
wire n_6294;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_5845;
wire n_5945;
wire n_804;
wire n_2390;
wire n_6246;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_7250;
wire n_1782;
wire n_5755;
wire n_5600;
wire n_8043;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_3208;
wire n_4944;
wire n_2195;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_4715;
wire n_6123;
wire n_6901;
wire n_4935;
wire n_4694;
wire n_6841;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_6922;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_1672;
wire n_6774;
wire n_6271;
wire n_6489;
wire n_1925;
wire n_4407;
wire n_7402;
wire n_737;
wire n_3517;
wire n_4045;
wire n_3893;
wire n_4598;
wire n_3061;
wire n_2945;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_5993;
wire n_8054;
wire n_6716;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_7914;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_7113;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_2840;
wire n_6779;
wire n_8010;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_7216;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_6762;
wire n_6178;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_7706;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_6458;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_7642;
wire n_6577;
wire n_6740;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_6315;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_7156;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_6910;
wire n_6262;
wire n_7604;
wire n_2827;
wire n_1177;
wire n_7703;
wire n_3515;
wire n_1150;
wire n_6319;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_6536;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_6978;
wire n_5351;
wire n_5909;
wire n_6093;
wire n_4543;
wire n_740;
wire n_7378;
wire n_4157;
wire n_6845;
wire n_6947;
wire n_4229;
wire n_5293;
wire n_6099;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_1401;
wire n_7498;
wire n_1516;
wire n_3846;
wire n_6321;
wire n_3512;
wire n_6819;
wire n_5201;
wire n_2029;
wire n_7501;
wire n_5890;
wire n_6415;
wire n_6465;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_7931;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_6899;
wire n_7549;
wire n_7373;
wire n_7895;
wire n_832;
wire n_6592;
wire n_3049;
wire n_6626;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_7740;
wire n_3679;
wire n_5891;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_4930;
wire n_5623;
wire n_6944;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_4593;
wire n_7238;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_7572;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_5990;
wire n_7043;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_7760;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_4231;
wire n_6281;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_6846;
wire n_6311;
wire n_930;
wire n_7590;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_7048;
wire n_6886;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_6593;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_7176;
wire n_7682;
wire n_990;
wire n_6231;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_6932;
wire n_6746;
wire n_7901;
wire n_870;
wire n_5395;
wire n_1253;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_1693;
wire n_6446;
wire n_7980;
wire n_3802;
wire n_3256;
wire n_6996;
wire n_7218;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_6749;
wire n_2188;
wire n_1989;
wire n_7005;
wire n_2802;
wire n_7732;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_2425;
wire n_6777;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_7405;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_7922;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_6310;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_6683;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_2047;
wire n_6229;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_6907;
wire n_3989;
wire n_7144;
wire n_2490;
wire n_7089;
wire n_7286;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_4254;
wire n_6177;
wire n_1996;
wire n_6332;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_5982;
wire n_1158;
wire n_2248;
wire n_7403;
wire n_5011;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_6696;
wire n_753;
wire n_3925;
wire n_3180;
wire n_7343;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_6116;
wire n_7859;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_7972;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_7916;
wire n_3717;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_6167;
wire n_1884;
wire n_8008;
wire n_6170;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_6307;
wire n_6094;
wire n_2038;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_6155;
wire n_7269;
wire n_6267;
wire n_7787;
wire n_1833;
wire n_3903;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_7507;
wire n_7159;
wire n_5378;
wire n_6028;
wire n_1417;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_4648;
wire n_3094;
wire n_6299;
wire n_6813;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_7425;
wire n_6669;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_1748;
wire n_8058;
wire n_3504;
wire n_6638;
wire n_7719;
wire n_4272;
wire n_5615;
wire n_6220;
wire n_1025;
wire n_7562;
wire n_2930;
wire n_3111;
wire n_6985;
wire n_7619;
wire n_7170;
wire n_1885;
wire n_7366;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_7935;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_6772;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_6318;
wire n_2353;
wire n_4099;
wire n_7918;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_6916;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_6651;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_7845;
wire n_5550;
wire n_3911;
wire n_7536;
wire n_7472;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_6604;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_5881;
wire n_1370;
wire n_7222;
wire n_1786;
wire n_7942;
wire n_6473;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_7725;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_6483;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_7647;
wire n_2645;
wire n_3904;
wire n_8036;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_7300;
wire n_6697;
wire n_7875;
wire n_6975;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_7643;
wire n_4733;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_5955;
wire n_7242;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_6076;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_7778;
wire n_758;
wire n_5851;
wire n_7073;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_6390;
wire n_5796;
wire n_772;
wire n_2806;
wire n_6665;
wire n_7224;
wire n_770;
wire n_3028;
wire n_7746;
wire n_3662;
wire n_2981;
wire n_6958;
wire n_3076;
wire n_886;
wire n_7563;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_6549;
wire n_6297;
wire n_6523;
wire n_6653;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_4687;
wire n_2836;
wire n_7531;
wire n_1404;
wire n_5492;
wire n_5995;
wire n_2378;
wire n_7721;
wire n_887;
wire n_7192;
wire n_5905;
wire n_2655;
wire n_4600;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_1467;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_8057;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_2370;
wire n_2612;
wire n_7527;
wire n_7417;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_6582;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_7388;
wire n_3568;
wire n_3850;
wire n_1230;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_7090;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_7227;
wire n_7415;
wire n_824;
wire n_6745;
wire n_6972;
wire n_4297;
wire n_8030;
wire n_6052;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_6240;
wire n_6347;
wire n_5020;
wire n_7689;
wire n_6511;
wire n_5297;
wire n_7121;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_1970;
wire n_6358;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_6603;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_7534;
wire n_1957;
wire n_4354;
wire n_6986;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_5959;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_8031;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_6396;
wire n_5642;
wire n_4581;
wire n_6890;
wire n_4377;
wire n_7827;
wire n_2143;
wire n_905;
wire n_6109;
wire n_4792;
wire n_7731;
wire n_3842;
wire n_1680;
wire n_993;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_6770;
wire n_2654;
wire n_3036;
wire n_7943;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_7081;
wire n_2711;
wire n_7132;
wire n_4199;
wire n_5885;
wire n_6663;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_7319;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_7828;
wire n_4773;
wire n_7940;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_6621;
wire n_7001;
wire n_4822;
wire n_1214;
wire n_850;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_6783;
wire n_825;
wire n_6066;
wire n_3785;
wire n_6897;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_7708;
wire n_4055;
wire n_2178;
wire n_5968;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_6497;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_7108;
wire n_6470;
wire n_1796;
wire n_7333;
wire n_2082;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_7371;
wire n_7463;
wire n_6573;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_6693;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_7285;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_6409;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_7954;
wire n_1465;
wire n_2622;
wire n_7951;
wire n_2658;
wire n_7552;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_6130;
wire n_4603;
wire n_7273;
wire n_1523;
wire n_7231;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_7449;
wire n_7772;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_7239;
wire n_1493;
wire n_5690;
wire n_7050;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_6623;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_7597;
wire n_5801;
wire n_6047;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_6652;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_6970;
wire n_6921;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_7674;
wire n_3171;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_4540;
wire n_6344;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_6624;
wire n_6956;
wire n_4284;
wire n_6305;
wire n_1005;
wire n_1947;
wire n_6209;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_7126;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_7329;
wire n_7408;
wire n_2650;
wire n_7107;
wire n_5652;
wire n_6457;
wire n_987;
wire n_7690;
wire n_7123;
wire n_5499;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_6950;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_6694;
wire n_3497;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_7229;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_1181;
wire n_7258;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_6856;
wire n_3996;
wire n_1049;
wire n_6466;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_7709;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_6820;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_2368;
wire n_8041;
wire n_4175;
wire n_6438;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_7332;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_7512;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_7766;
wire n_6469;
wire n_6700;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_6758;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_7955;
wire n_811;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_7287;
wire n_5497;
wire n_880;
wire n_6464;
wire n_6356;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_7637;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_7127;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_1382;
wire n_5408;
wire n_7801;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_7959;
wire n_7019;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_8071;
wire n_1427;
wire n_2745;
wire n_7735;
wire n_8004;
wire n_1080;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_5964;
wire n_6004;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_5234;
wire n_4431;
wire n_7546;
wire n_2421;
wire n_1136;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_6588;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_7575;
wire n_3571;
wire n_7083;
wire n_1775;
wire n_2410;
wire n_7720;
wire n_6222;
wire n_1093;
wire n_1783;
wire n_6268;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_6456;
wire n_7521;
wire n_3407;
wire n_5992;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_1185;
wire n_7187;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_6467;
wire n_5079;
wire n_6540;
wire n_6625;
wire n_1453;
wire n_6336;
wire n_6796;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_6541;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_7603;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_6757;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_8006;
wire n_7636;
wire n_2955;
wire n_5592;
wire n_6954;
wire n_2158;
wire n_6938;
wire n_4609;
wire n_7866;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_7205;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_7020;
wire n_7990;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_5157;
wire n_3525;
wire n_2100;
wire n_3314;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_6421;
wire n_1905;
wire n_7407;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_7148;
wire n_6328;
wire n_5956;
wire n_5287;
wire n_6236;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_3907;
wire n_1103;
wire n_2875;
wire n_6144;
wire n_3338;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_2219;
wire n_6835;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_7104;
wire n_7124;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_2304;
wire n_7799;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_7513;
wire n_3572;
wire n_6602;
wire n_3886;
wire n_6708;
wire n_6645;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_6242;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_7692;
wire n_5174;
wire n_4234;
wire n_7469;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_7560;
wire n_7645;
wire n_1397;
wire n_3236;
wire n_901;
wire n_3141;
wire n_2755;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_7082;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_5570;
wire n_6418;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5927;
wire n_7495;
wire n_7392;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_6400;
wire n_2607;
wire n_7666;
wire n_7945;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_6941;
wire n_1943;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_1320;
wire n_7543;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_7877;
wire n_7963;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_6398;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_7284;
wire n_1983;
wire n_7264;
wire n_5391;
wire n_1938;
wire n_7737;
wire n_6537;
wire n_2472;
wire n_7328;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_3957;
wire n_2894;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_7135;
wire n_6224;
wire n_6578;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_7024;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_1692;
wire n_1084;
wire n_6614;
wire n_5912;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_8035;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_7152;
wire n_2200;
wire n_6165;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_6567;
wire n_2670;
wire n_2700;
wire n_5910;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_3134;
wire n_5965;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_7240;
wire n_7570;
wire n_896;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_2084;
wire n_4875;
wire n_7817;
wire n_5682;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_8002;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_7237;
wire n_5681;
wire n_6877;
wire n_7423;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_4040;
wire n_1640;
wire n_2406;
wire n_7617;
wire n_806;
wire n_2141;
wire n_5316;
wire n_7718;
wire n_6940;
wire n_7396;
wire n_5703;
wire n_7835;
wire n_833;
wire n_6320;
wire n_7998;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_7561;
wire n_6810;
wire n_7842;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_6202;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_7163;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_7236;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_7130;
wire n_1241;
wire n_7201;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_7491;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_6792;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_5979;
wire n_3558;
wire n_7559;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_6044;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_4726;
wire n_7678;
wire n_1045;
wire n_5907;
wire n_786;
wire n_1559;
wire n_6045;
wire n_1872;
wire n_6731;
wire n_7526;
wire n_5040;
wire n_6063;
wire n_1325;
wire n_6504;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_7004;
wire n_7821;
wire n_1727;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_5977;
wire n_7879;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_7696;
wire n_6003;
wire n_6684;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_6600;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_6673;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_3621;
wire n_6031;
wire n_6962;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_7887;
wire n_7246;
wire n_4365;
wire n_6060;
wire n_1882;
wire n_7929;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_7270;
wire n_3758;
wire n_5417;
wire n_6967;
wire n_2587;
wire n_7550;
wire n_3199;
wire n_3339;
wire n_6742;
wire n_6853;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_6691;
wire n_7087;
wire n_1953;
wire n_6191;
wire n_4741;
wire n_6172;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_7851;
wire n_6894;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_6834;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_5842;
wire n_6817;
wire n_6927;
wire n_5814;
wire n_2814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_6215;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_6517;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_7862;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_5064;
wire n_7825;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_6966;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_6722;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_6035;
wire n_1994;
wire n_957;
wire n_7874;
wire n_7622;
wire n_2566;
wire n_6364;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_7102;
wire n_7420;
wire n_2906;
wire n_4342;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_6061;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_7831;
wire n_2914;
wire n_5786;
wire n_8065;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_6419;
wire n_1083;
wire n_7784;
wire n_5768;
wire n_3553;
wire n_2465;
wire n_7225;
wire n_2275;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_1721;
wire n_3494;
wire n_6244;
wire n_6900;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_1028;
wire n_6942;
wire n_7705;
wire n_2106;
wire n_2265;
wire n_7228;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_7932;
wire n_4409;
wire n_7509;
wire n_5872;
wire n_6862;
wire n_7058;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_708;
wire n_1973;
wire n_6840;
wire n_3181;
wire n_6338;
wire n_5700;
wire n_1500;
wire n_6037;
wire n_7981;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_5874;
wire n_6266;
wire n_6488;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_7164;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_7018;
wire n_5873;
wire n_7975;
wire n_1085;
wire n_2042;
wire n_771;
wire n_6317;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_7167;
wire n_6480;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_7865;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_2035;
wire n_7844;
wire n_7134;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_6875;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_7079;
wire n_981;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_2071;
wire n_1144;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_7267;
wire n_4599;
wire n_3233;
wire n_997;
wire n_4437;
wire n_5222;
wire n_7316;
wire n_7850;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_7812;
wire n_1198;
wire n_7103;
wire n_4061;
wire n_7460;
wire n_6176;
wire n_2174;
wire n_6367;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_7056;
wire n_6572;
wire n_1133;
wire n_4429;
wire n_7962;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_7813;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_6080;
wire n_4865;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_7473;
wire n_7200;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_7688;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_7795;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_7038;
wire n_2001;
wire n_7723;
wire n_4341;
wire n_1629;
wire n_7404;
wire n_5368;
wire n_4263;
wire n_1819;
wire n_1260;
wire n_3555;
wire n_7059;
wire n_7450;
wire n_915;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_812;
wire n_6145;
wire n_1131;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_1006;
wire n_3110;
wire n_7271;
wire n_1632;
wire n_7826;
wire n_5933;
wire n_1888;
wire n_6204;
wire n_1311;
wire n_7076;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_6842;
wire n_3467;
wire n_6866;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_6451;
wire n_3039;
wire n_1226;
wire n_6514;
wire n_3740;
wire n_5996;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_7105;
wire n_1958;
wire n_7049;
wire n_5903;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_6710;
wire n_4984;
wire n_2579;
wire n_6345;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_7535;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_7057;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_6957;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_7944;
wire n_7262;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_7016;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_6379;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_8044;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_6719;
wire n_7178;
wire n_1380;
wire n_2847;
wire n_7506;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_6232;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_2521;
wire n_1099;
wire n_8052;
wire n_4578;
wire n_2211;
wire n_6362;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_7142;
wire n_1285;
wire n_1985;
wire n_6326;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_1172;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_7241;
wire n_7247;
wire n_7172;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_7235;
wire n_2447;
wire n_6239;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_7340;
wire n_6974;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_6713;
wire n_8064;
wire n_7657;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_7096;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_1163;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_2495;
wire n_7999;
wire n_6087;
wire n_7593;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_8068;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_7764;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_5969;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_1211;
wire n_6454;
wire n_5022;
wire n_7041;
wire n_7307;
wire n_5670;
wire n_1280;
wire n_6041;
wire n_6918;
wire n_3296;
wire n_7350;
wire n_5276;
wire n_8012;
wire n_1445;
wire n_7672;
wire n_2551;
wire n_6664;
wire n_1526;
wire n_5047;
wire n_7318;
wire n_2985;
wire n_1978;
wire n_6472;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_5879;
wire n_8062;
wire n_4403;
wire n_5238;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_6375;
wire n_6352;
wire n_1054;
wire n_7063;
wire n_1956;
wire n_7047;
wire n_4139;
wire n_6632;
wire n_4549;
wire n_6238;
wire n_1986;
wire n_8038;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_6081;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_6724;
wire n_5429;
wire n_6545;
wire n_813;
wire n_6705;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_7074;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_6591;
wire n_2207;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_6946;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_6289;
wire n_7037;
wire n_3748;
wire n_3272;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_7599;
wire n_7928;
wire n_4393;
wire n_1162;
wire n_6532;
wire n_821;
wire n_4372;
wire n_1068;
wire n_7293;
wire n_982;
wire n_5640;
wire n_7600;
wire n_932;
wire n_2831;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3978;
wire n_3317;
wire n_6721;
wire n_5560;
wire n_6644;
wire n_2123;
wire n_1697;
wire n_6512;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_6108;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_7614;
wire n_2941;
wire n_1278;
wire n_7839;
wire n_5108;
wire n_7347;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_4337;
wire n_4130;
wire n_5941;
wire n_2009;
wire n_7759;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_6340;
wire n_3092;
wire n_1289;
wire n_6219;
wire n_3055;
wire n_6706;
wire n_7479;
wire n_3966;
wire n_2866;
wire n_7395;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_7078;
wire n_2580;
wire n_6761;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_3384;
wire n_1950;
wire n_6811;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_4478;
wire n_1662;
wire n_7372;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_6868;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_7174;
wire n_5202;
wire n_4965;
wire n_8021;
wire n_3346;
wire n_7803;
wire n_1896;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_6659;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_6011;
wire n_1886;
wire n_4371;
wire n_6225;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_7086;
wire n_728;
wire n_3415;
wire n_1063;
wire n_6648;
wire n_4607;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_3918;
wire n_5876;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_6601;
wire n_7920;
wire n_7810;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_7025;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_6826;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_5856;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_8014;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_7768;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_7982;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_6879;
wire n_1295;
wire n_7567;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_7684;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_7370;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_2151;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_6306;
wire n_6720;
wire n_6888;
wire n_826;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_1714;
wire n_718;
wire n_6095;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_5311;
wire n_6590;
wire n_2089;
wire n_7583;
wire n_3522;
wire n_6559;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_2148;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3975;
wire n_3018;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_1838;
wire n_6287;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_7353;
wire n_2002;
wire n_2138;
wire n_7758;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_5772;
wire n_7571;
wire n_4775;
wire n_2208;
wire n_5884;
wire n_6671;
wire n_6812;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_2134;
wire n_1176;
wire n_7792;
wire n_7510;
wire n_6662;
wire n_5603;
wire n_6525;
wire n_7422;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_7109;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5924;
wire n_1505;
wire n_7253;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_6702;
wire n_3620;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_2520;
wire n_7380;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_7749;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_7574;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_6005;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_6169;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_7713;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_6936;
wire n_2589;
wire n_4535;
wire n_7704;
wire n_7487;
wire n_755;
wire n_6302;
wire n_2442;
wire n_7641;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_7203;
wire n_1137;
wire n_7169;
wire n_7670;
wire n_3612;
wire n_4695;
wire n_6848;
wire n_2545;
wire n_3509;
wire n_5919;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_7439;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_6343;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_6850;
wire n_5005;
wire n_6098;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_6979;
wire n_7815;
wire n_7934;
wire n_723;
wire n_3144;
wire n_3244;
wire n_6865;
wire n_1141;
wire n_1268;
wire n_7276;
wire n_8056;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_6747;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_3640;
wire n_3481;
wire n_995;
wire n_1159;
wire n_6640;
wire n_2250;
wire n_3033;
wire n_6142;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_2374;
wire n_1681;
wire n_6034;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_7233;
wire n_7602;
wire n_7034;
wire n_5220;
wire n_1618;
wire n_7390;
wire n_4867;
wire n_6870;
wire n_6221;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_1653;
wire n_7881;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_6071;
wire n_2920;
wire n_773;
wire n_7598;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_6833;
wire n_6793;
wire n_1169;
wire n_6767;
wire n_6295;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_8053;
wire n_848;
wire n_6385;
wire n_7426;
wire n_4247;
wire n_7045;
wire n_3169;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_7984;
wire n_6788;
wire n_2023;
wire n_7014;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_7220;
wire n_1323;
wire n_6709;
wire n_2627;
wire n_4422;
wire n_960;
wire n_6550;
wire n_6712;
wire n_7416;
wire n_6143;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_6743;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_7465;
wire n_5967;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_2515;
wire n_7936;
wire n_6084;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_7738;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_5966;
wire n_2201;
wire n_725;
wire n_6634;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_7462;
wire n_4635;
wire n_994;
wire n_5735;
wire n_7490;
wire n_2278;
wire n_7545;
wire n_1020;
wire n_1273;
wire n_7160;
wire n_7464;
wire n_4214;
wire n_6919;
wire n_3448;
wire n_7805;
wire n_7115;
wire n_7295;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_7348;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_6681;
wire n_6104;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_1095;
wire n_6973;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_7453;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_7946;
wire n_1499;
wire n_1409;
wire n_5877;
wire n_7681;
wire n_6018;
wire n_6619;
wire n_5189;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_8042;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_7210;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_4155;
wire n_6854;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_1216;
wire n_2716;
wire n_6032;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_7855;
wire n_3043;
wire n_8050;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_6981;
wire n_2220;
wire n_7065;
wire n_2577;
wire n_1262;
wire n_3529;
wire n_3238;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_6122;
wire n_2790;
wire n_7911;
wire n_6765;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_7330;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_7336;
wire n_2373;
wire n_1472;
wire n_7446;
wire n_3628;
wire n_7854;
wire n_5454;
wire n_800;
wire n_4734;
wire n_7493;
wire n_7357;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_7923;
wire n_2244;
wire n_6439;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_7714;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_6406;
wire n_7440;
wire n_1102;
wire n_1963;
wire n_6945;
wire n_3790;
wire n_7029;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_6618;
wire n_6474;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_7317;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_6000;
wire n_2782;
wire n_3977;
wire n_8055;
wire n_6816;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_6425;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_6492;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_6046;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_4007;
wire n_4949;
wire n_6852;
wire n_2642;
wire n_4239;
wire n_7468;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_6251;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_6869;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_7621;
wire n_7359;
wire n_3321;
wire n_5809;
wire n_2567;
wire n_2322;
wire n_3377;
wire n_2727;
wire n_7924;
wire n_4782;
wire n_1321;
wire n_7659;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_7153;
wire n_1235;
wire n_2759;
wire n_7836;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_7280;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_7886;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_6631;
wire n_4469;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_6228;
wire n_6711;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_8017;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_7275;
wire n_2885;
wire n_7195;
wire n_6102;
wire n_6274;
wire n_3097;
wire n_7007;
wire n_2062;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_6072;
wire n_7610;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_7259;
wire n_1607;
wire n_1454;
wire n_6353;
wire n_4953;
wire n_6992;
wire n_2348;
wire n_2944;
wire n_6818;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_5932;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_7539;
wire n_841;
wire n_1476;
wire n_3391;
wire n_7616;
wire n_1800;
wire n_6498;
wire n_1463;
wire n_3458;
wire n_7775;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_7930;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_6976;
wire n_6304;
wire n_5236;
wire n_853;
wire n_7640;
wire n_875;
wire n_5012;
wire n_1678;
wire n_6864;
wire n_7969;
wire n_3787;
wire n_1256;
wire n_7548;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_5025;
wire n_933;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_3135;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_8000;
wire n_1217;
wire n_7197;
wire n_5645;
wire n_3990;
wire n_7393;
wire n_6917;
wire n_6937;
wire n_7591;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_7727;
wire n_7358;
wire n_988;
wire n_2796;
wire n_7324;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_6301;
wire n_1204;
wire n_1132;
wire n_6929;
wire n_1327;
wire n_955;
wire n_8045;
wire n_7729;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_7565;
wire n_1120;
wire n_6699;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_2290;
wire n_7382;
wire n_4811;
wire n_2048;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_2005;
wire n_4857;
wire n_7437;
wire n_6677;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_7618;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_6764;
wire n_863;
wire n_3774;
wire n_5733;
wire n_6780;
wire n_2910;
wire n_6620;
wire n_6597;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_866;
wire n_7282;
wire n_2287;
wire n_6586;
wire n_6333;
wire n_7139;
wire n_5791;
wire n_5727;
wire n_761;
wire n_5946;
wire n_5997;
wire n_2492;
wire n_7953;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_5975;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_6510;
wire n_3334;
wire n_5938;
wire n_6237;
wire n_5602;
wire n_5097;
wire n_844;
wire n_4985;
wire n_7751;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_7581;
wire n_888;
wire n_6360;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_7346;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_7579;
wire n_4025;
wire n_7428;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_7150;
wire n_7155;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_6475;
wire n_7015;
wire n_3982;
wire n_7283;
wire n_7699;
wire n_6314;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_7249;
wire n_3796;
wire n_6394;
wire n_6964;
wire n_3840;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_4246;
wire n_7432;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_6752;
wire n_1156;
wire n_6426;
wire n_2600;
wire n_984;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_7612;
wire n_7494;
wire n_868;
wire n_4353;
wire n_735;
wire n_6350;
wire n_4787;
wire n_7736;
wire n_5633;
wire n_1218;
wire n_5664;
wire n_7589;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_2429;
wire n_985;
wire n_2440;
wire n_6054;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_6235;
wire n_7843;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_7756;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_7700;
wire n_4451;
wire n_4332;
wire n_810;
wire n_7555;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_7988;
wire n_3563;
wire n_6513;
wire n_7500;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_5925;
wire n_2909;
wire n_754;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_6330;
wire n_3187;
wire n_3218;
wire n_6802;
wire n_861;
wire n_6909;
wire n_7157;
wire n_6908;
wire n_857;
wire n_7411;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_7266;
wire n_2221;
wire n_8046;
wire n_7871;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_4210;
wire n_1010;
wire n_4981;
wire n_6477;
wire n_6263;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_2709;
wire n_7198;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_7794;
wire n_2185;
wire n_6038;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_6605;
wire n_5032;
wire n_1899;
wire n_6313;
wire n_784;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_7145;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_2098;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_5920;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_7994;
wire n_1449;
wire n_4703;
wire n_7349;
wire n_7715;
wire n_2419;
wire n_6180;
wire n_5683;
wire n_6349;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_1742;
wire n_4030;

BUFx3_ASAP7_75t_L g708 ( 
.A(n_248),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_697),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_504),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_222),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_699),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_443),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_447),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_542),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_218),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_368),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_607),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_78),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_596),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_67),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_15),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_420),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_699),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_166),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_55),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_414),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_579),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_61),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_356),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_280),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_354),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_51),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_446),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_94),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_177),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_277),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_492),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_114),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_426),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_501),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_238),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_546),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_56),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_9),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_659),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_696),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_82),
.Y(n_748)
);

CKINVDCx14_ASAP7_75t_R g749 ( 
.A(n_228),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_371),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_290),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_637),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_133),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_283),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_693),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_176),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_281),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_245),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_320),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_434),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_511),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_84),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_701),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_20),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_106),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_625),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_163),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_582),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_502),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_549),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_340),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_617),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_210),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_565),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_467),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_9),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_552),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_252),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_492),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_491),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_692),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_461),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_128),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_625),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_605),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_131),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_438),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_380),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_34),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_209),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_707),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_449),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_270),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_112),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_695),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_258),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_606),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_389),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_80),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_470),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_267),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_22),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_413),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_195),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_377),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_21),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_116),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_707),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_24),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_387),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_443),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_619),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_688),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_143),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_585),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_302),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_318),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_334),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_343),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_549),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_140),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_461),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_594),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_250),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_98),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_692),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_512),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_475),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_446),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_79),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_69),
.Y(n_831)
);

CKINVDCx16_ASAP7_75t_R g832 ( 
.A(n_518),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_485),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_143),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_615),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_25),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_252),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_702),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_129),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_517),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_128),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_579),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_486),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_184),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_113),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_547),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_131),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_264),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_604),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_358),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_654),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_392),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_330),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_593),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_195),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_257),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_453),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_361),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_298),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_569),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_524),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_691),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_478),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_340),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_295),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_341),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_67),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_444),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_502),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_74),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_251),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_655),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_420),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_300),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_455),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_323),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_0),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_387),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_540),
.Y(n_879)
);

CKINVDCx14_ASAP7_75t_R g880 ( 
.A(n_683),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_36),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_619),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_411),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_536),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_390),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_497),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_25),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_266),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_164),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_306),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_380),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_651),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_576),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_480),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_140),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_671),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_412),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_481),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_466),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_332),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_467),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_528),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_33),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_46),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_177),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_276),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_559),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_650),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_175),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_278),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_347),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_7),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_687),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_156),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_173),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_370),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_64),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_200),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_343),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_504),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_578),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_188),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_661),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_522),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_49),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_172),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_436),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_602),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_522),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_636),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_42),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_635),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_319),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_433),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_543),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_348),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_201),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_154),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_167),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_69),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_563),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_432),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_541),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_388),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_78),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_45),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_463),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_519),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_685),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_159),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_341),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_686),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_61),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_56),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_18),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_274),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_386),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_267),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_572),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_568),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_638),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_690),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_654),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_474),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_370),
.Y(n_965)
);

BUFx8_ASAP7_75t_SL g966 ( 
.A(n_168),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_537),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_200),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_160),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_441),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_315),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_569),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_475),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_531),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_342),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_547),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_424),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_186),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_544),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_37),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_366),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_170),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_138),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_151),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_401),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_118),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_469),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_198),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_506),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_253),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_506),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_349),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_697),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_454),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_245),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_515),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_657),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_41),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_591),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_186),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_178),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_410),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_677),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_388),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_305),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_351),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_12),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_593),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_587),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_643),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_289),
.Y(n_1011)
);

BUFx5_ASAP7_75t_L g1012 ( 
.A(n_43),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_111),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_540),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_684),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_271),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_665),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_303),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_563),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_535),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_353),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_271),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_595),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_221),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_286),
.Y(n_1025)
);

BUFx5_ASAP7_75t_L g1026 ( 
.A(n_337),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_120),
.Y(n_1027)
);

CKINVDCx14_ASAP7_75t_R g1028 ( 
.A(n_325),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_643),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_257),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_192),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_576),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_614),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_418),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_442),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_689),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_630),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_641),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_489),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_SL g1040 ( 
.A(n_573),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_317),
.Y(n_1041)
);

BUFx2_ASAP7_75t_SL g1042 ( 
.A(n_305),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_354),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_375),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_529),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_89),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_73),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_426),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_611),
.Y(n_1049)
);

CKINVDCx16_ASAP7_75t_R g1050 ( 
.A(n_249),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_250),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_284),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_27),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_119),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_501),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_369),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_169),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_298),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_413),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_657),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_97),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_5),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_362),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_410),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_281),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_103),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_574),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_705),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_323),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_74),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_524),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_150),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_296),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_199),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_130),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_98),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_29),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_232),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_693),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_407),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_363),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_259),
.Y(n_1082)
);

CKINVDCx16_ASAP7_75t_R g1083 ( 
.A(n_489),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_517),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_399),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_460),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_405),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_535),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_342),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_508),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_507),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_34),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_335),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_411),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_163),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_24),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_134),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_670),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_311),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_25),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_543),
.Y(n_1101)
);

BUFx5_ASAP7_75t_L g1102 ( 
.A(n_19),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_108),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_690),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_326),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_55),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_316),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_164),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_122),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_599),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_203),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_75),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_586),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_285),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_642),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_337),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_302),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_339),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_32),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_191),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_132),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_424),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_181),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_552),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_49),
.Y(n_1125)
);

BUFx8_ASAP7_75t_SL g1126 ( 
.A(n_453),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_92),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_384),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_405),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_3),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_278),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_133),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_694),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_597),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_590),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_470),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_316),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_583),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_373),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_520),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_347),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_279),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_677),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_471),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_482),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_41),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_233),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_647),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_435),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_541),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_490),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_119),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_627),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_518),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_32),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_202),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_402),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_557),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_355),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_393),
.Y(n_1160)
);

CKINVDCx16_ASAP7_75t_R g1161 ( 
.A(n_241),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_95),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_412),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_236),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_612),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_221),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_678),
.Y(n_1167)
);

CKINVDCx16_ASAP7_75t_R g1168 ( 
.A(n_310),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_401),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_105),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_610),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_157),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_651),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_646),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_180),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_486),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_166),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_270),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_448),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_615),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_505),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_452),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_568),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_389),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_351),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_594),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_621),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_269),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_30),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_335),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_333),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_37),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_372),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_637),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_495),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_240),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_689),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_287),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_635),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_645),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_38),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_365),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_515),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_91),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_274),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_174),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_14),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_676),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_398),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_275),
.Y(n_1210)
);

BUFx8_ASAP7_75t_SL g1211 ( 
.A(n_403),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_631),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_251),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_686),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_240),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_670),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_105),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_659),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_326),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_529),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_406),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_698),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_661),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_468),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_449),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_121),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_630),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_169),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_220),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_458),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_588),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_586),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_107),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_94),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_671),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_237),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_22),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_87),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_403),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_436),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_37),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_575),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_649),
.Y(n_1243)
);

CKINVDCx14_ASAP7_75t_R g1244 ( 
.A(n_369),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_107),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_308),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_293),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_679),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_641),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_249),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_452),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_137),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_966),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1012),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_966),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1126),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1126),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1012),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1211),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1211),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_733),
.B(n_0),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_887),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1012),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_749),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1012),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_749),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_880),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_880),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1028),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1012),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1028),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1244),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1012),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1244),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1012),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1012),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_740),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_722),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1012),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1012),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_764),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1102),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1102),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1102),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1102),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_741),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1102),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_776),
.Y(n_1289)
);

BUFx10_ASAP7_75t_L g1290 ( 
.A(n_887),
.Y(n_1290)
);

INVx4_ASAP7_75t_R g1291 ( 
.A(n_1040),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_789),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_806),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_809),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1102),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1102),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_881),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1102),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1102),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1102),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_903),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1026),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_912),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1026),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_751),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_821),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_931),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_946),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_954),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_980),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1026),
.Y(n_1311)
);

CKINVDCx16_ASAP7_75t_R g1312 ( 
.A(n_832),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1125),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_925),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_887),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1026),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1026),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1146),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_751),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1026),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1237),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_708),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_887),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_896),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1250),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1026),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_832),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1026),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1026),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1252),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_887),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1026),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_816),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_982),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_910),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_887),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_712),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_712),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_712),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_712),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_709),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_712),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_712),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_712),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_895),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_895),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_895),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_887),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_713),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_714),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_717),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_895),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_895),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_725),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_727),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_895),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_728),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_895),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1001),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_729),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1001),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1001),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1001),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_731),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1092),
.B(n_0),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1021),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1092),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_734),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_735),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1001),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1092),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_736),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1001),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1001),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1092),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1092),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_737),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_739),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_715),
.Y(n_1379)
);

CKINVDCx16_ASAP7_75t_R g1380 ( 
.A(n_910),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_742),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1170),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1092),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_743),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1092),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1201),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_746),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1174),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1201),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_752),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_753),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_754),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_755),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_1009),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1201),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1201),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_756),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_757),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_760),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_761),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1201),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1245),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_762),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1201),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_763),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1201),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_745),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_816),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_745),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_745),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1009),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_765),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_836),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_715),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_836),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_766),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_767),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_836),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_768),
.Y(n_1419)
);

CKINVDCx14_ASAP7_75t_R g1420 ( 
.A(n_850),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_708),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_781),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_769),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_772),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_747),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_747),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_747),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1253),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_774),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_775),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1253),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_778),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_779),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_779),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_779),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_780),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_708),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_799),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_799),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1253),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_799),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1022),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_783),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1022),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_781),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_804),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1050),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_784),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_850),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_804),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_804),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_785),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_786),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_787),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_811),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_811),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_811),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_720),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_813),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_791),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_813),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_795),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_813),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_889),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_889),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1050),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_864),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_796),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_720),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_889),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_893),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_798),
.Y(n_1472)
);

CKINVDCx14_ASAP7_75t_R g1473 ( 
.A(n_864),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_720),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_1083),
.Y(n_1475)
);

XNOR2xp5_ASAP7_75t_L g1476 ( 
.A(n_925),
.B(n_1),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_800),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_893),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_801),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_893),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_803),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_908),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_875),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_875),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1083),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1161),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_908),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_807),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_908),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1161),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_917),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_810),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1203),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1029),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_917),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_917),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_812),
.Y(n_1497)
);

CKINVDCx16_ASAP7_75t_R g1498 ( 
.A(n_1168),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_943),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_943),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1029),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_943),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_967),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_909),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_817),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_822),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1168),
.Y(n_1507)
);

INVxp33_ASAP7_75t_SL g1508 ( 
.A(n_1203),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_967),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_823),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_909),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_827),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_967),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_970),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1227),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_970),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_828),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_970),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_972),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_830),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_831),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_833),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_972),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_972),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_1040),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_978),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_834),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_978),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_838),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_978),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_987),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_987),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_987),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_839),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_841),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_843),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_845),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_848),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_721),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_994),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_994),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_852),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_994),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_996),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_853),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_996),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_854),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_759),
.B(n_1),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_996),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1058),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_856),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1058),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1058),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_SL g1554 ( 
.A(n_711),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1065),
.Y(n_1555)
);

BUFx5_ASAP7_75t_L g1556 ( 
.A(n_1029),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1065),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1065),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_876),
.B(n_2),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1076),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_860),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1076),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1076),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_721),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_862),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_777),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_711),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_863),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_865),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1195),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1045),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1195),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_872),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1195),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1212),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1212),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1227),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1212),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1045),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_777),
.Y(n_1580)
);

BUFx2_ASAP7_75t_SL g1581 ( 
.A(n_750),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_794),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1045),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_733),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_802),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_873),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_711),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_802),
.Y(n_1588)
);

CKINVDCx16_ASAP7_75t_R g1589 ( 
.A(n_711),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_874),
.Y(n_1590)
);

BUFx2_ASAP7_75t_SL g1591 ( 
.A(n_750),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_877),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_878),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_877),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_955),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_955),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_884),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_998),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_998),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1007),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1007),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_885),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_748),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1053),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_886),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1053),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1062),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1062),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1077),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1077),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1096),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_890),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1096),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_891),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_892),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1100),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1155),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1100),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_894),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_897),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_L g1621 ( 
.A(n_759),
.B(n_2),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_902),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_905),
.Y(n_1623)
);

CKINVDCx16_ASAP7_75t_R g1624 ( 
.A(n_748),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1106),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_911),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1155),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1106),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1119),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1119),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_794),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1130),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1130),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1192),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1192),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1207),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_913),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1207),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1241),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1241),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_710),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_915),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_916),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_918),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_710),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_716),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_744),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_716),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_718),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_718),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_719),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_719),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_920),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_921),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1189),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_922),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_723),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_723),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_724),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_724),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_923),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_730),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1042),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_924),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_926),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_840),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_730),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_927),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_732),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_732),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_928),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_929),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_738),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_930),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_932),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_933),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_936),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_937),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_738),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_770),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_940),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_941),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_942),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_945),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_770),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1189),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_771),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_947),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_771),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_773),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_948),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_951),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_748),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_773),
.Y(n_1694)
);

INVxp33_ASAP7_75t_L g1695 ( 
.A(n_788),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_788),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_953),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_956),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_792),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_792),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_958),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_793),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_793),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_962),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_963),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_797),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_964),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_797),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_814),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_814),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1583),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1583),
.Y(n_1712)
);

INVxp33_ASAP7_75t_L g1713 ( 
.A(n_1511),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1611),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1539),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1647),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1525),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1577),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1579),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1579),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1375),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1375),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1385),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1385),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1386),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1386),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1325),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1389),
.Y(n_1728)
);

CKINVDCx20_ASAP7_75t_R g1729 ( 
.A(n_1564),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1566),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1389),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1395),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1259),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1330),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1395),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1396),
.Y(n_1736)
);

INVxp33_ASAP7_75t_SL g1737 ( 
.A(n_1265),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1341),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1396),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1349),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1401),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1350),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1580),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1582),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1525),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1401),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1404),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1404),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1351),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1406),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1406),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1365),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1354),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1421),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1421),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1355),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1631),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1437),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1357),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1437),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1474),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1474),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1360),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1494),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1494),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1501),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1666),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_1278),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1364),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1501),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1331),
.Y(n_1771)
);

CKINVDCx20_ASAP7_75t_R g1772 ( 
.A(n_1287),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1331),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1368),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1626),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1371),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1371),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1255),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1255),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1259),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1369),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1264),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1336),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1264),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1266),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1266),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1336),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1271),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1271),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1306),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1274),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1372),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1274),
.Y(n_1793)
);

INVxp33_ASAP7_75t_L g1794 ( 
.A(n_1684),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1276),
.Y(n_1795)
);

INVxp33_ASAP7_75t_SL g1796 ( 
.A(n_1267),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1276),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1277),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1663),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1377),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1277),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1280),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1280),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1281),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1281),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_SL g1806 ( 
.A(n_1603),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1284),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1284),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1286),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1286),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1324),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1378),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1381),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1384),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1288),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1288),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1295),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1387),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1295),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1296),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1296),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1298),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1603),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1298),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1299),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1299),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1337),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1337),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1334),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1338),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1338),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1339),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1366),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1382),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1339),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1390),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1693),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1340),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1704),
.Y(n_1839)
);

CKINVDCx16_ASAP7_75t_R g1840 ( 
.A(n_1312),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1340),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1312),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1342),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1391),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1342),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1392),
.Y(n_1846)
);

CKINVDCx16_ASAP7_75t_R g1847 ( 
.A(n_1335),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1393),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1388),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1397),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1402),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1343),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1693),
.Y(n_1853)
);

CKINVDCx20_ASAP7_75t_R g1854 ( 
.A(n_1275),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1398),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1343),
.Y(n_1856)
);

CKINVDCx20_ASAP7_75t_R g1857 ( 
.A(n_1314),
.Y(n_1857)
);

CKINVDCx16_ASAP7_75t_R g1858 ( 
.A(n_1335),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1344),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1344),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1345),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1315),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1556),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1345),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1346),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1399),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1346),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1400),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1347),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1403),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1405),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1347),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1352),
.Y(n_1873)
);

INVxp33_ASAP7_75t_SL g1874 ( 
.A(n_1268),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1352),
.Y(n_1875)
);

INVxp67_ASAP7_75t_SL g1876 ( 
.A(n_1322),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1353),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1353),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1356),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1348),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1356),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1412),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1587),
.Y(n_1883)
);

CKINVDCx16_ASAP7_75t_R g1884 ( 
.A(n_1380),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1348),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1411),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1315),
.Y(n_1887)
);

CKINVDCx20_ASAP7_75t_R g1888 ( 
.A(n_1442),
.Y(n_1888)
);

CKINVDCx20_ASAP7_75t_R g1889 ( 
.A(n_1444),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1322),
.Y(n_1890)
);

CKINVDCx14_ASAP7_75t_R g1891 ( 
.A(n_1420),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1416),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1358),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1417),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1419),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1587),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1305),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1556),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1358),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1423),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1367),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1424),
.Y(n_1902)
);

INVxp33_ASAP7_75t_SL g1903 ( 
.A(n_1269),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1458),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1359),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1359),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1362),
.Y(n_1907)
);

INVxp33_ASAP7_75t_L g1908 ( 
.A(n_1445),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1362),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1363),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1429),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1447),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1363),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1370),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1430),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1458),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1466),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1370),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1373),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1373),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1374),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1432),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1436),
.Y(n_1923)
);

INVxp67_ASAP7_75t_SL g1924 ( 
.A(n_1469),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1374),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1367),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1439),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1556),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1485),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1439),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1439),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1443),
.Y(n_1932)
);

INVxp33_ASAP7_75t_SL g1933 ( 
.A(n_1270),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1448),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1439),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1305),
.Y(n_1936)
);

CKINVDCx20_ASAP7_75t_R g1937 ( 
.A(n_1486),
.Y(n_1937)
);

INVxp33_ASAP7_75t_L g1938 ( 
.A(n_1408),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1439),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1480),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1480),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1480),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1452),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1315),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1480),
.Y(n_1945)
);

CKINVDCx20_ASAP7_75t_R g1946 ( 
.A(n_1490),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1469),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1480),
.Y(n_1948)
);

INVxp67_ASAP7_75t_SL g1949 ( 
.A(n_1571),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1563),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1408),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1563),
.Y(n_1952)
);

CKINVDCx16_ASAP7_75t_R g1953 ( 
.A(n_1380),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1563),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1507),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1563),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1453),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1563),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1572),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1572),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1572),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1394),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1572),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1572),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1315),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1394),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1454),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1610),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1610),
.Y(n_1969)
);

CKINVDCx16_ASAP7_75t_R g1970 ( 
.A(n_1475),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1315),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1376),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1460),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1610),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1610),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1475),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1462),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1610),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1327),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1633),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1633),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1633),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1633),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1449),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1633),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_1498),
.Y(n_1986)
);

INVxp67_ASAP7_75t_SL g1987 ( 
.A(n_1571),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1703),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1468),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1472),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1703),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1703),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1449),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1477),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1376),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1567),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1567),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1703),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1479),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1703),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1376),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1361),
.Y(n_2002)
);

INVxp33_ASAP7_75t_SL g2003 ( 
.A(n_1272),
.Y(n_2003)
);

INVxp33_ASAP7_75t_L g2004 ( 
.A(n_1515),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1376),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1589),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1361),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1481),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1361),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1488),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1589),
.Y(n_2011)
);

CKINVDCx20_ASAP7_75t_R g2012 ( 
.A(n_1473),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1302),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1302),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1317),
.Y(n_2015)
);

INVxp33_ASAP7_75t_L g2016 ( 
.A(n_1515),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1317),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1320),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1320),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1326),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1617),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1326),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1332),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1332),
.Y(n_2024)
);

INVxp33_ASAP7_75t_SL g2025 ( 
.A(n_1273),
.Y(n_2025)
);

INVxp33_ASAP7_75t_L g2026 ( 
.A(n_1559),
.Y(n_2026)
);

INVxp33_ASAP7_75t_L g2027 ( 
.A(n_1617),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1492),
.Y(n_2028)
);

CKINVDCx16_ASAP7_75t_R g2029 ( 
.A(n_1624),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1627),
.Y(n_2030)
);

INVxp67_ASAP7_75t_L g2031 ( 
.A(n_1319),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1556),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1556),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1556),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1556),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1556),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1627),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1556),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1497),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_SL g2040 ( 
.A(n_1263),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1376),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1655),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1584),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1655),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1584),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1588),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_1383),
.Y(n_2047)
);

CKINVDCx16_ASAP7_75t_R g2048 ( 
.A(n_1554),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_1686),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1505),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1506),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1588),
.Y(n_2052)
);

INVxp67_ASAP7_75t_SL g2053 ( 
.A(n_1383),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1592),
.Y(n_2054)
);

INVxp67_ASAP7_75t_L g2055 ( 
.A(n_1333),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_1467),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1592),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_1554),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1594),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1483),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1594),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1510),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1595),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1595),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1596),
.Y(n_2065)
);

CKINVDCx20_ASAP7_75t_R g2066 ( 
.A(n_1254),
.Y(n_2066)
);

CKINVDCx16_ASAP7_75t_R g2067 ( 
.A(n_1554),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1596),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1599),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1599),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1600),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1512),
.Y(n_2072)
);

CKINVDCx20_ASAP7_75t_R g2073 ( 
.A(n_1256),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_1484),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1517),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_1263),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1600),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1520),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1601),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1601),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1607),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1607),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1383),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1609),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1609),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1613),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1727),
.Y(n_2087)
);

AOI22x1_ASAP7_75t_SL g2088 ( 
.A1(n_2021),
.A2(n_846),
.B1(n_899),
.B2(n_840),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1771),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1734),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1752),
.B(n_1581),
.Y(n_2091)
);

INVx2_ASAP7_75t_SL g2092 ( 
.A(n_1716),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1719),
.B(n_1581),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2026),
.B(n_1883),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_2032),
.A2(n_1285),
.B(n_1283),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1887),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1783),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1887),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1738),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1783),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1887),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2026),
.A2(n_1508),
.B1(n_846),
.B2(n_959),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_1773),
.B(n_1425),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1776),
.Y(n_2104)
);

BUFx6f_ASAP7_75t_L g2105 ( 
.A(n_1887),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1777),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1720),
.B(n_1425),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1897),
.A2(n_899),
.B1(n_989),
.B2(n_959),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_2031),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1944),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2055),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1754),
.B(n_1591),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_1799),
.A2(n_1282),
.B1(n_1289),
.B2(n_1279),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1778),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1755),
.B(n_1591),
.Y(n_2115)
);

INVxp33_ASAP7_75t_SL g2116 ( 
.A(n_2049),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1944),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1787),
.Y(n_2118)
);

NOR2x1_ASAP7_75t_L g2119 ( 
.A(n_2076),
.B(n_1262),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1779),
.Y(n_2120)
);

BUFx8_ASAP7_75t_L g2121 ( 
.A(n_1886),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1782),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1936),
.A2(n_999),
.B1(n_1027),
.B2(n_989),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1896),
.B(n_1698),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1784),
.Y(n_2125)
);

OAI22x1_ASAP7_75t_SL g2126 ( 
.A1(n_2021),
.A2(n_1027),
.B1(n_1036),
.B2(n_999),
.Y(n_2126)
);

AND2x2_ASAP7_75t_SL g2127 ( 
.A(n_1717),
.B(n_1262),
.Y(n_2127)
);

INVx5_ASAP7_75t_L g2128 ( 
.A(n_1944),
.Y(n_2128)
);

CKINVDCx8_ASAP7_75t_R g2129 ( 
.A(n_1840),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1944),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1787),
.Y(n_2131)
);

OA21x2_ASAP7_75t_L g2132 ( 
.A1(n_2002),
.A2(n_1285),
.B(n_1283),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1880),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1785),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1880),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_2001),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2056),
.B(n_1504),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1758),
.B(n_1407),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1786),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1788),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1789),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_2076),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_2001),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1885),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1760),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_2001),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1791),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1733),
.B(n_1780),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1885),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2060),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1793),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1795),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1775),
.B(n_1707),
.Y(n_2153)
);

BUFx3_ASAP7_75t_L g2154 ( 
.A(n_1761),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1797),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_2001),
.Y(n_2156)
);

AND2x2_ASAP7_75t_SL g2157 ( 
.A(n_1842),
.B(n_815),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_2074),
.Y(n_2158)
);

INVx6_ASAP7_75t_L g2159 ( 
.A(n_1863),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1901),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1951),
.A2(n_1057),
.B1(n_1060),
.B2(n_1036),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1901),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1762),
.B(n_1407),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1839),
.B(n_1521),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1926),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_1764),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_2048),
.B(n_1522),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1931),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1876),
.B(n_1527),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1798),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_2033),
.A2(n_1300),
.B(n_1304),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1890),
.B(n_1529),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1765),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1931),
.Y(n_2174)
);

OAI22x1_ASAP7_75t_L g2175 ( 
.A1(n_1984),
.A2(n_1476),
.B1(n_1414),
.B2(n_1422),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1801),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1802),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1904),
.B(n_1534),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1993),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1803),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1766),
.B(n_1438),
.Y(n_2181)
);

BUFx8_ASAP7_75t_L g2182 ( 
.A(n_1806),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_2058),
.B(n_1697),
.Y(n_2183)
);

AND2x6_ASAP7_75t_L g2184 ( 
.A(n_1863),
.B(n_1300),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1804),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1948),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1862),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2067),
.B(n_1535),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_1770),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1948),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1952),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1862),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1862),
.Y(n_2193)
);

AOI22x1_ASAP7_75t_SL g2194 ( 
.A1(n_2030),
.A2(n_1060),
.B1(n_1073),
.B2(n_1057),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_1965),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1965),
.Y(n_2196)
);

BUFx2_ASAP7_75t_L g2197 ( 
.A(n_1962),
.Y(n_2197)
);

INVx4_ASAP7_75t_L g2198 ( 
.A(n_1898),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1952),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1971),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1721),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1722),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_1711),
.B(n_1438),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1805),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1723),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1807),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1714),
.B(n_1536),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1808),
.Y(n_2208)
);

INVx6_ASAP7_75t_L g2209 ( 
.A(n_1898),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_1971),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1712),
.B(n_1409),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2043),
.B(n_1450),
.Y(n_2212)
);

CKINVDCx20_ASAP7_75t_R g2213 ( 
.A(n_1768),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1809),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_1847),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2086),
.B(n_1450),
.Y(n_2216)
);

BUFx8_ASAP7_75t_SL g2217 ( 
.A(n_1857),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1810),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_2085),
.B(n_1455),
.Y(n_2219)
);

CKINVDCx11_ASAP7_75t_R g2220 ( 
.A(n_1857),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_1858),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_1823),
.A2(n_1293),
.B1(n_1294),
.B2(n_1292),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1740),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1972),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1815),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_1742),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1916),
.B(n_1409),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_1745),
.A2(n_1097),
.B1(n_1166),
.B2(n_1073),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1972),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_2034),
.A2(n_1311),
.B(n_1304),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1995),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_1995),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1724),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2005),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1725),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1816),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1726),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1817),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1884),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1924),
.B(n_1537),
.Y(n_2240)
);

BUFx12f_ASAP7_75t_L g2241 ( 
.A(n_1745),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1947),
.B(n_1701),
.Y(n_2242)
);

OA21x2_ASAP7_75t_L g2243 ( 
.A1(n_2007),
.A2(n_1316),
.B(n_1311),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_2005),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_2041),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1728),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_1769),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_1953),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1731),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1732),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1800),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1949),
.B(n_1410),
.Y(n_2252)
);

OAI21x1_ASAP7_75t_L g2253 ( 
.A1(n_2035),
.A2(n_1328),
.B(n_1316),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1735),
.Y(n_2254)
);

CKINVDCx8_ASAP7_75t_R g2255 ( 
.A(n_1970),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_1781),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1736),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1819),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_2045),
.B(n_1455),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1820),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_1792),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_2041),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1821),
.Y(n_2263)
);

BUFx6f_ASAP7_75t_L g2264 ( 
.A(n_2083),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1822),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1812),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1824),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_1962),
.Y(n_2268)
);

INVx4_ASAP7_75t_L g2269 ( 
.A(n_1928),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1825),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1826),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1739),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_SL g2273 ( 
.A1(n_2030),
.A2(n_1476),
.B1(n_1166),
.B2(n_1204),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2013),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_2083),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_1928),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1741),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1746),
.Y(n_2278)
);

BUFx2_ASAP7_75t_L g2279 ( 
.A(n_1966),
.Y(n_2279)
);

OA21x2_ASAP7_75t_L g2280 ( 
.A1(n_2009),
.A2(n_1329),
.B(n_1328),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_1891),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1747),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_1848),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1748),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2084),
.B(n_2046),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1827),
.Y(n_2286)
);

BUFx12f_ASAP7_75t_L g2287 ( 
.A(n_1749),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_1828),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2014),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_1830),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2015),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1987),
.B(n_1538),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1831),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2052),
.B(n_1461),
.Y(n_2294)
);

INVxp67_ASAP7_75t_L g2295 ( 
.A(n_1871),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2027),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1832),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1835),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2017),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2018),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_2019),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2020),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1750),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2082),
.B(n_1461),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1751),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_SL g2306 ( 
.A1(n_2037),
.A2(n_1204),
.B1(n_1220),
.B2(n_1097),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_2022),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_1794),
.B(n_1542),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2023),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_2024),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1838),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1813),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1841),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1843),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_1845),
.A2(n_1329),
.B(n_1502),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_1852),
.Y(n_2316)
);

BUFx6f_ASAP7_75t_L g2317 ( 
.A(n_1856),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1859),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2054),
.B(n_1410),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1860),
.Y(n_2320)
);

INVx5_ASAP7_75t_L g2321 ( 
.A(n_2040),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1861),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1864),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1865),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_1867),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2047),
.B(n_1545),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2057),
.B(n_1413),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_1938),
.A2(n_1225),
.B1(n_1228),
.B2(n_1220),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_1927),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1869),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1872),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_1892),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1873),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1875),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1877),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_1966),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1878),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2081),
.B(n_1502),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2059),
.B(n_1413),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2061),
.B(n_1415),
.Y(n_2340)
);

OA21x2_ASAP7_75t_L g2341 ( 
.A1(n_1879),
.A2(n_1893),
.B(n_1881),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1899),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_1930),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_2027),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1905),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2053),
.B(n_1547),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1906),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_1935),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1907),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_1909),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1794),
.B(n_1705),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_1939),
.Y(n_2352)
);

AOI22xp5_ASAP7_75t_L g2353 ( 
.A1(n_1938),
.A2(n_1228),
.B1(n_1231),
.B2(n_1225),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1910),
.Y(n_2354)
);

INVx5_ASAP7_75t_L g2355 ( 
.A(n_2040),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1913),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_1914),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_1837),
.B(n_1551),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1918),
.Y(n_2359)
);

BUFx8_ASAP7_75t_L g2360 ( 
.A(n_1806),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1919),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1920),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1921),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2063),
.B(n_1415),
.Y(n_2364)
);

AND2x6_ASAP7_75t_L g2365 ( 
.A(n_2036),
.B(n_815),
.Y(n_2365)
);

OA21x2_ASAP7_75t_L g2366 ( 
.A1(n_1925),
.A2(n_1523),
.B(n_1509),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1968),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_1940),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2064),
.B(n_1418),
.Y(n_2369)
);

OAI22xp5_ASAP7_75t_SL g2370 ( 
.A1(n_2037),
.A2(n_1246),
.B1(n_1231),
.B2(n_904),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1969),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_1853),
.A2(n_1301),
.B1(n_1303),
.B2(n_1297),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1941),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2065),
.B(n_1418),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2042),
.A2(n_1246),
.B1(n_904),
.B2(n_726),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_1814),
.B(n_1692),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1942),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_1945),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1950),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1974),
.Y(n_2380)
);

OAI21x1_ASAP7_75t_L g2381 ( 
.A1(n_2038),
.A2(n_1523),
.B(n_1509),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1954),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1975),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_1976),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1956),
.B(n_1561),
.Y(n_2385)
);

OAI21x1_ASAP7_75t_L g2386 ( 
.A1(n_1958),
.A2(n_1543),
.B(n_1533),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1959),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1960),
.Y(n_2388)
);

INVx4_ASAP7_75t_L g2389 ( 
.A(n_2040),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_1818),
.B(n_1565),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1978),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1980),
.Y(n_2392)
);

AND2x6_ASAP7_75t_L g2393 ( 
.A(n_1961),
.B(n_818),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_SL g2394 ( 
.A1(n_2042),
.A2(n_876),
.B1(n_1248),
.B2(n_726),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_1963),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1836),
.B(n_1568),
.Y(n_2396)
);

BUFx3_ASAP7_75t_L g2397 ( 
.A(n_1964),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1981),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1982),
.B(n_1569),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1983),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_1976),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1985),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1988),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_1991),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_1992),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1998),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2000),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2068),
.Y(n_2408)
);

BUFx3_ASAP7_75t_L g2409 ( 
.A(n_2069),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2070),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2071),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2004),
.A2(n_1308),
.B1(n_1309),
.B2(n_1307),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2077),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2079),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2080),
.B(n_1573),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_1806),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2004),
.B(n_1426),
.Y(n_2417)
);

INVx5_ASAP7_75t_L g2418 ( 
.A(n_2029),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_1844),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1973),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2039),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1846),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_1850),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_1855),
.B(n_1533),
.Y(n_2424)
);

BUFx12f_ASAP7_75t_L g2425 ( 
.A(n_1749),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_1866),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_1713),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1868),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_1870),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2016),
.A2(n_1313),
.B1(n_1318),
.B2(n_1310),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1882),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1894),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1895),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2010),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2028),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2050),
.Y(n_2436)
);

BUFx2_ASAP7_75t_L g2437 ( 
.A(n_1979),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2051),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2062),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2072),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_1753),
.B(n_1586),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1753),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_1713),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_SL g2444 ( 
.A1(n_2044),
.A2(n_1248),
.B1(n_790),
.B2(n_805),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1756),
.Y(n_2445)
);

OAI22x1_ASAP7_75t_SL g2446 ( 
.A1(n_2044),
.A2(n_1258),
.B1(n_1260),
.B2(n_1257),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_1756),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_1759),
.B(n_1543),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1759),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_1979),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2016),
.B(n_1426),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_1763),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1763),
.Y(n_2453)
);

OAI21x1_ASAP7_75t_L g2454 ( 
.A1(n_1737),
.A2(n_1558),
.B(n_1553),
.Y(n_2454)
);

CKINVDCx20_ASAP7_75t_R g2455 ( 
.A(n_1768),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1774),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1774),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_1900),
.A2(n_1621),
.B1(n_1548),
.B2(n_1493),
.Y(n_2458)
);

CKINVDCx8_ASAP7_75t_R g2459 ( 
.A(n_1900),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_1908),
.B(n_1427),
.Y(n_2460)
);

INVx4_ASAP7_75t_L g2461 ( 
.A(n_2078),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_1902),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_1902),
.Y(n_2463)
);

AND2x4_ASAP7_75t_L g2464 ( 
.A(n_1911),
.B(n_1553),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_1911),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1915),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1915),
.Y(n_2467)
);

CKINVDCx16_ASAP7_75t_R g2468 ( 
.A(n_2012),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1922),
.B(n_1590),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_1922),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_1923),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2078),
.B(n_1593),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1923),
.Y(n_2473)
);

AND2x4_ASAP7_75t_L g2474 ( 
.A(n_2075),
.B(n_1558),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_1737),
.B(n_1691),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_1932),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_1932),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_1934),
.A2(n_1574),
.B(n_1428),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_1934),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_1796),
.A2(n_1321),
.B1(n_1379),
.B2(n_1597),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_1943),
.B(n_1602),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1943),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_1957),
.Y(n_2483)
);

HB1xp67_ASAP7_75t_L g2484 ( 
.A(n_1718),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_1957),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_1967),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_1967),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_1977),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_1977),
.A2(n_790),
.B1(n_805),
.B2(n_782),
.Y(n_2489)
);

OAI22xp5_ASAP7_75t_SL g2490 ( 
.A1(n_1888),
.A2(n_808),
.B1(n_824),
.B2(n_782),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_1718),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_1989),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_1986),
.Y(n_2493)
);

OA21x2_ASAP7_75t_L g2494 ( 
.A1(n_1989),
.A2(n_1574),
.B(n_1428),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_1990),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_1986),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_1990),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_1994),
.Y(n_2498)
);

AOI22x1_ASAP7_75t_SL g2499 ( 
.A1(n_1715),
.A2(n_824),
.B1(n_883),
.B2(n_808),
.Y(n_2499)
);

AND2x4_ASAP7_75t_L g2500 ( 
.A(n_1994),
.B(n_1427),
.Y(n_2500)
);

AOI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_1999),
.A2(n_883),
.B1(n_1008),
.B2(n_935),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_1999),
.Y(n_2502)
);

CKINVDCx6p67_ASAP7_75t_R g2503 ( 
.A(n_2012),
.Y(n_2503)
);

OA21x2_ASAP7_75t_L g2504 ( 
.A1(n_2008),
.A2(n_1433),
.B(n_1431),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2008),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2075),
.B(n_1605),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_1908),
.B(n_1431),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_1996),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_1996),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_1997),
.Y(n_2510)
);

INVx2_ASAP7_75t_SL g2511 ( 
.A(n_1772),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_1796),
.Y(n_2512)
);

BUFx3_ASAP7_75t_L g2513 ( 
.A(n_1874),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_1997),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2006),
.B(n_1433),
.Y(n_2515)
);

INVx5_ASAP7_75t_L g2516 ( 
.A(n_1874),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_1903),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2006),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_1903),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_1933),
.B(n_1612),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2011),
.B(n_1434),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_1772),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1933),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2381),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2381),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2366),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2366),
.Y(n_2527)
);

INVxp67_ASAP7_75t_L g2528 ( 
.A(n_2137),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2386),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2366),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2366),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2386),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2095),
.Y(n_2533)
);

HB1xp67_ASAP7_75t_L g2534 ( 
.A(n_2092),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2092),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2109),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2109),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2095),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2171),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2315),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2171),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2230),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2150),
.Y(n_2543)
);

NOR2x1_ASAP7_75t_L g2544 ( 
.A(n_2389),
.B(n_2441),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2145),
.B(n_1585),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2230),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2253),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2253),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2116),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2091),
.B(n_1614),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_2315),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2315),
.Y(n_2552)
);

NAND3xp33_ASAP7_75t_L g2553 ( 
.A(n_2094),
.B(n_2207),
.C(n_2458),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2315),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2145),
.B(n_1585),
.Y(n_2555)
);

XOR2xp5_ASAP7_75t_L g2556 ( 
.A(n_2126),
.B(n_1790),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2132),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2145),
.B(n_1598),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2132),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2091),
.B(n_1615),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2103),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2103),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2103),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2103),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2137),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2132),
.Y(n_2566)
);

BUFx2_ASAP7_75t_L g2567 ( 
.A(n_2150),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2132),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2133),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2133),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2135),
.Y(n_2571)
);

INVx6_ASAP7_75t_L g2572 ( 
.A(n_2159),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2158),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2135),
.Y(n_2574)
);

CKINVDCx20_ASAP7_75t_R g2575 ( 
.A(n_2213),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2144),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2243),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2243),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2460),
.B(n_1619),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2144),
.Y(n_2580)
);

BUFx2_ASAP7_75t_L g2581 ( 
.A(n_2158),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2149),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2149),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2111),
.Y(n_2584)
);

NAND2xp33_ASAP7_75t_SL g2585 ( 
.A(n_2332),
.B(n_1261),
.Y(n_2585)
);

CKINVDCx8_ASAP7_75t_R g2586 ( 
.A(n_2468),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2243),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2160),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2160),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2243),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2162),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2162),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2280),
.Y(n_2593)
);

INVxp67_ASAP7_75t_L g2594 ( 
.A(n_2427),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2280),
.Y(n_2595)
);

INVx1_ASAP7_75t_SL g2596 ( 
.A(n_2443),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2280),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2460),
.B(n_1620),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2280),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2154),
.B(n_1598),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2148),
.B(n_1622),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2484),
.Y(n_2602)
);

AND2x6_ASAP7_75t_L g2603 ( 
.A(n_2416),
.B(n_818),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2341),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2454),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2119),
.A2(n_2025),
.B1(n_2003),
.B2(n_1637),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2097),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2341),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2097),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2341),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2114),
.B(n_1623),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2454),
.Y(n_2612)
);

INVxp67_ASAP7_75t_L g2613 ( 
.A(n_2491),
.Y(n_2613)
);

OA21x2_ASAP7_75t_L g2614 ( 
.A1(n_2263),
.A2(n_1435),
.B(n_1434),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2276),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2341),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2114),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2507),
.B(n_1642),
.Y(n_2618)
);

INVxp67_ASAP7_75t_L g2619 ( 
.A(n_2296),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2120),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2120),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2154),
.B(n_1604),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2122),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2122),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2097),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2154),
.B(n_1604),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2125),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2344),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2125),
.B(n_1643),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2100),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2134),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2134),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2196),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2100),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2100),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2507),
.B(n_1644),
.Y(n_2636)
);

INVx1_ASAP7_75t_SL g2637 ( 
.A(n_2455),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2139),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2139),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2276),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2140),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2140),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2141),
.B(n_1653),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2118),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2141),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2147),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2118),
.Y(n_2647)
);

XNOR2xp5_ASAP7_75t_L g2648 ( 
.A(n_2306),
.B(n_1715),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2147),
.B(n_1654),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2151),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2196),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2151),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2276),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2152),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2152),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2118),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2515),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2276),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2131),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2417),
.B(n_1656),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2417),
.B(n_1661),
.Y(n_2661)
);

OAI22xp5_ASAP7_75t_SL g2662 ( 
.A1(n_2273),
.A2(n_1889),
.B1(n_1912),
.B2(n_1888),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2155),
.Y(n_2663)
);

BUFx2_ASAP7_75t_L g2664 ( 
.A(n_2521),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2155),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2196),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2276),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2170),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2170),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2131),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2131),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2176),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2159),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_L g2674 ( 
.A(n_2159),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2173),
.B(n_1606),
.Y(n_2675)
);

BUFx8_ASAP7_75t_L g2676 ( 
.A(n_2437),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2176),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2177),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2177),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2180),
.Y(n_2680)
);

OAI21x1_ASAP7_75t_L g2681 ( 
.A1(n_2348),
.A2(n_1451),
.B(n_1441),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2180),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2515),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2451),
.B(n_1664),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2185),
.B(n_1665),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2185),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2204),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2521),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2217),
.Y(n_2689)
);

INVx3_ASAP7_75t_L g2690 ( 
.A(n_2196),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2204),
.B(n_1668),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2206),
.B(n_1671),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2451),
.B(n_1672),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2206),
.B(n_1674),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_2521),
.Y(n_2695)
);

XOR2xp5_ASAP7_75t_L g2696 ( 
.A(n_2126),
.B(n_1790),
.Y(n_2696)
);

XOR2xp5_ASAP7_75t_L g2697 ( 
.A(n_2273),
.B(n_1811),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2208),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2208),
.B(n_1675),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2220),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2521),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2214),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2203),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2196),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2159),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2203),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2173),
.B(n_1606),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2214),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2218),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2209),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2173),
.B(n_2285),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2231),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2218),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2225),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2424),
.B(n_2003),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2225),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2203),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2209),
.Y(n_2718)
);

OAI21x1_ASAP7_75t_L g2719 ( 
.A1(n_2348),
.A2(n_1451),
.B(n_1441),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2285),
.B(n_1608),
.Y(n_2720)
);

CKINVDCx8_ASAP7_75t_R g2721 ( 
.A(n_2468),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2203),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2236),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2236),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2238),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2209),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2238),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2168),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2258),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2168),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2424),
.B(n_2448),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_2209),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2174),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2258),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2260),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2424),
.B(n_2025),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2260),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2265),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2265),
.Y(n_2739)
);

BUFx2_ASAP7_75t_L g2740 ( 
.A(n_2179),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_2424),
.B(n_1676),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2301),
.Y(n_2742)
);

OA21x2_ASAP7_75t_L g2743 ( 
.A1(n_2263),
.A2(n_1440),
.B(n_1435),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2227),
.B(n_1677),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2301),
.Y(n_2745)
);

INVxp67_ASAP7_75t_L g2746 ( 
.A(n_2308),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2270),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2242),
.B(n_1678),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2270),
.Y(n_2749)
);

HB1xp67_ASAP7_75t_L g2750 ( 
.A(n_2448),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2174),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2271),
.B(n_1681),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2221),
.Y(n_2753)
);

INVx1_ASAP7_75t_SL g2754 ( 
.A(n_2437),
.Y(n_2754)
);

AND2x6_ASAP7_75t_L g2755 ( 
.A(n_2416),
.B(n_819),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2271),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2274),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2274),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2289),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2301),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_2239),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2289),
.B(n_1682),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2186),
.Y(n_2763)
);

BUFx6f_ASAP7_75t_L g2764 ( 
.A(n_2307),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2186),
.Y(n_2765)
);

HB1xp67_ASAP7_75t_L g2766 ( 
.A(n_2448),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2190),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2190),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2291),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2291),
.B(n_1683),
.Y(n_2770)
);

NAND2xp33_ASAP7_75t_L g2771 ( 
.A(n_2365),
.B(n_1688),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2299),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2448),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2153),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2299),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2231),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2464),
.B(n_1291),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2300),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2450),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2300),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2191),
.Y(n_2781)
);

HB1xp67_ASAP7_75t_L g2782 ( 
.A(n_2464),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2191),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2302),
.B(n_1383),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2500),
.A2(n_2011),
.B1(n_2073),
.B2(n_2066),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2285),
.B(n_1608),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2307),
.Y(n_2787)
);

HB1xp67_ASAP7_75t_L g2788 ( 
.A(n_2464),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2302),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2309),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2199),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2309),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2408),
.B(n_1383),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2408),
.B(n_1263),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2199),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2227),
.B(n_2252),
.Y(n_2796)
);

XOR2xp5_ASAP7_75t_L g2797 ( 
.A(n_2306),
.B(n_1811),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2478),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2285),
.B(n_1616),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_SL g2800 ( 
.A(n_2461),
.B(n_2066),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2142),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2165),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2409),
.B(n_2142),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2415),
.B(n_1889),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2307),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2478),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2478),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2478),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2248),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2165),
.Y(n_2810)
);

CKINVDCx8_ASAP7_75t_R g2811 ( 
.A(n_2418),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2494),
.Y(n_2812)
);

CKINVDCx20_ASAP7_75t_R g2813 ( 
.A(n_2087),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2494),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2231),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2231),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2494),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2263),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2267),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2231),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2142),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2267),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2287),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2464),
.B(n_968),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2494),
.Y(n_2825)
);

AOI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2500),
.A2(n_2073),
.B1(n_1937),
.B2(n_1946),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2511),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2267),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2184),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2244),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2408),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2408),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2272),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2164),
.B(n_1912),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_2184),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2272),
.Y(n_2836)
);

BUFx8_ASAP7_75t_L g2837 ( 
.A(n_2450),
.Y(n_2837)
);

INVxp67_ASAP7_75t_L g2838 ( 
.A(n_2474),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_SL g2839 ( 
.A(n_2461),
.B(n_1854),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2272),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2277),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2138),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2252),
.B(n_1263),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2093),
.B(n_2112),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2277),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2277),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2278),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2278),
.Y(n_2848)
);

OA21x2_ASAP7_75t_L g2849 ( 
.A1(n_2278),
.A2(n_1446),
.B(n_1440),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2282),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2282),
.Y(n_2851)
);

BUFx8_ASAP7_75t_L g2852 ( 
.A(n_2493),
.Y(n_2852)
);

NOR2xp33_ASAP7_75t_L g2853 ( 
.A(n_2469),
.B(n_1917),
.Y(n_2853)
);

CKINVDCx8_ASAP7_75t_R g2854 ( 
.A(n_2418),
.Y(n_2854)
);

HB1xp67_ASAP7_75t_L g2855 ( 
.A(n_2474),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2184),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2244),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2282),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2409),
.B(n_1616),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2348),
.A2(n_1451),
.B(n_1441),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2287),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2284),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2244),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2284),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2112),
.B(n_1695),
.Y(n_2865)
);

INVx3_ASAP7_75t_L g2866 ( 
.A(n_2244),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2093),
.B(n_1290),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2284),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2472),
.B(n_1917),
.Y(n_2869)
);

BUFx6f_ASAP7_75t_L g2870 ( 
.A(n_2184),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2303),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2409),
.B(n_1628),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2115),
.B(n_1628),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2474),
.B(n_969),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2244),
.Y(n_2875)
);

OAI21x1_ASAP7_75t_L g2876 ( 
.A1(n_2348),
.A2(n_1540),
.B(n_1478),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2511),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2303),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2102),
.B(n_935),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2303),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2305),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2522),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2184),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2305),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2305),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2211),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2211),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2212),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2115),
.B(n_1290),
.Y(n_2889)
);

BUFx6f_ASAP7_75t_L g2890 ( 
.A(n_2184),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2245),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2245),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2410),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2089),
.B(n_1290),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2410),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2089),
.B(n_1290),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2522),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2474),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2184),
.Y(n_2899)
);

XOR2xp5_ASAP7_75t_L g2900 ( 
.A(n_2088),
.B(n_1829),
.Y(n_2900)
);

BUFx6f_ASAP7_75t_L g2901 ( 
.A(n_2245),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2212),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2212),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2212),
.Y(n_2904)
);

INVxp67_ASAP7_75t_L g2905 ( 
.A(n_2475),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2216),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2520),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2481),
.B(n_1929),
.Y(n_2908)
);

HB1xp67_ASAP7_75t_L g2909 ( 
.A(n_2500),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_2425),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2216),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2216),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2411),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2245),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2411),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2138),
.B(n_1629),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2413),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2413),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2163),
.B(n_1629),
.Y(n_2919)
);

AND2x4_ASAP7_75t_L g2920 ( 
.A(n_2163),
.B(n_1634),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2414),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2216),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2219),
.Y(n_2923)
);

BUFx6f_ASAP7_75t_L g2924 ( 
.A(n_2245),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2500),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2219),
.Y(n_2926)
);

BUFx6f_ASAP7_75t_L g2927 ( 
.A(n_2262),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2262),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2414),
.Y(n_2929)
);

BUFx6f_ASAP7_75t_L g2930 ( 
.A(n_2262),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_2119),
.A2(n_1937),
.B1(n_1946),
.B2(n_1929),
.Y(n_2931)
);

OA21x2_ASAP7_75t_L g2932 ( 
.A1(n_2367),
.A2(n_1456),
.B(n_1446),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2311),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2319),
.B(n_1634),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2311),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2313),
.Y(n_2936)
);

BUFx6f_ASAP7_75t_L g2937 ( 
.A(n_2262),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2219),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2313),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2322),
.Y(n_2940)
);

INVx3_ASAP7_75t_L g2941 ( 
.A(n_2262),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2322),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2323),
.Y(n_2943)
);

OA21x2_ASAP7_75t_L g2944 ( 
.A1(n_2367),
.A2(n_1457),
.B(n_1456),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2323),
.Y(n_2945)
);

BUFx3_ASAP7_75t_L g2946 ( 
.A(n_2365),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2324),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2319),
.B(n_1635),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2324),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2219),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2259),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2330),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2330),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2333),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2365),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2104),
.B(n_1323),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2333),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2327),
.B(n_1635),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2345),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2345),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2259),
.Y(n_2961)
);

HB1xp67_ASAP7_75t_L g2962 ( 
.A(n_2215),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2259),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2259),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2349),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_SL g2966 ( 
.A(n_2461),
.B(n_1854),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2294),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2349),
.Y(n_2968)
);

BUFx6f_ASAP7_75t_L g2969 ( 
.A(n_2264),
.Y(n_2969)
);

AND2x6_ASAP7_75t_L g2970 ( 
.A(n_2416),
.B(n_819),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_SL g2971 ( 
.A(n_2516),
.B(n_973),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2294),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2361),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2294),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2104),
.B(n_1323),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2294),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2304),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2304),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2774),
.B(n_2905),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2818),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2614),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2550),
.B(n_2447),
.Y(n_2982)
);

INVx5_ASAP7_75t_L g2983 ( 
.A(n_2829),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_2550),
.B(n_2447),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2711),
.B(n_2106),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2907),
.B(n_2746),
.Y(n_2986)
);

INVx5_ASAP7_75t_L g2987 ( 
.A(n_2829),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2844),
.B(n_2504),
.Y(n_2988)
);

BUFx3_ASAP7_75t_L g2989 ( 
.A(n_2801),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2818),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2796),
.B(n_2504),
.Y(n_2991)
);

OAI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2553),
.A2(n_2470),
.B1(n_2486),
.B2(n_2479),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2796),
.A2(n_2365),
.B1(n_2504),
.B2(n_2393),
.Y(n_2993)
);

INVx2_ASAP7_75t_SL g2994 ( 
.A(n_2534),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_2689),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2819),
.Y(n_2996)
);

INVx2_ASAP7_75t_SL g2997 ( 
.A(n_2535),
.Y(n_2997)
);

BUFx3_ASAP7_75t_L g2998 ( 
.A(n_2801),
.Y(n_2998)
);

INVx3_ASAP7_75t_L g2999 ( 
.A(n_2533),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2560),
.B(n_2447),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2614),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2560),
.B(n_2447),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2614),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2614),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2743),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2829),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2720),
.A2(n_2365),
.B1(n_2504),
.B2(n_2393),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2819),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2748),
.B(n_2528),
.Y(n_3009)
);

CKINVDCx16_ASAP7_75t_R g3010 ( 
.A(n_2575),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2873),
.B(n_2169),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2822),
.Y(n_3012)
);

AOI22xp33_ASAP7_75t_SL g3013 ( 
.A1(n_2839),
.A2(n_2127),
.B1(n_2157),
.B2(n_2447),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2743),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2743),
.Y(n_3015)
);

OAI21xp33_ASAP7_75t_SL g3016 ( 
.A1(n_2617),
.A2(n_2621),
.B(n_2620),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_SL g3017 ( 
.A1(n_2966),
.A2(n_2127),
.B1(n_2800),
.B2(n_2157),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2743),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2849),
.Y(n_3019)
);

INVx4_ASAP7_75t_L g3020 ( 
.A(n_2615),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2873),
.B(n_2865),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2849),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2822),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2849),
.Y(n_3024)
);

OR2x2_ASAP7_75t_L g3025 ( 
.A(n_2543),
.B(n_2657),
.Y(n_3025)
);

NOR2x1p5_ASAP7_75t_L g3026 ( 
.A(n_2879),
.B(n_2519),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2828),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2849),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2828),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2865),
.B(n_2172),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2833),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2720),
.A2(n_2786),
.B1(n_2799),
.B2(n_2888),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2565),
.B(n_2376),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2833),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2607),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2536),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2925),
.B(n_2452),
.Y(n_3037)
);

NAND2xp33_ASAP7_75t_SL g3038 ( 
.A(n_2909),
.B(n_2452),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2617),
.B(n_2620),
.Y(n_3039)
);

BUFx3_ASAP7_75t_L g3040 ( 
.A(n_2821),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2621),
.B(n_2623),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2836),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2623),
.B(n_2178),
.Y(n_3043)
);

INVx8_ASAP7_75t_L g3044 ( 
.A(n_2603),
.Y(n_3044)
);

INVxp67_ASAP7_75t_SL g3045 ( 
.A(n_2615),
.Y(n_3045)
);

OR2x6_ASAP7_75t_L g3046 ( 
.A(n_2731),
.B(n_2419),
.Y(n_3046)
);

OR2x6_ASAP7_75t_L g3047 ( 
.A(n_2711),
.B(n_2419),
.Y(n_3047)
);

INVx3_ASAP7_75t_L g3048 ( 
.A(n_2533),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2594),
.B(n_2390),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2836),
.Y(n_3050)
);

INVx5_ASAP7_75t_L g3051 ( 
.A(n_2829),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2607),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2624),
.B(n_2240),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2609),
.Y(n_3054)
);

AND3x2_ASAP7_75t_L g3055 ( 
.A(n_2536),
.B(n_2281),
.C(n_2493),
.Y(n_3055)
);

INVx2_ASAP7_75t_SL g3056 ( 
.A(n_2567),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2609),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2840),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2625),
.Y(n_3059)
);

INVxp33_ASAP7_75t_SL g3060 ( 
.A(n_2689),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2840),
.Y(n_3061)
);

HB1xp67_ASAP7_75t_L g3062 ( 
.A(n_2567),
.Y(n_3062)
);

AOI22xp33_ASAP7_75t_L g3063 ( 
.A1(n_2720),
.A2(n_2365),
.B1(n_2393),
.B2(n_2310),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2711),
.B(n_2452),
.Y(n_3064)
);

INVx3_ASAP7_75t_L g3065 ( 
.A(n_2533),
.Y(n_3065)
);

BUFx10_ASAP7_75t_L g3066 ( 
.A(n_2853),
.Y(n_3066)
);

HB1xp67_ASAP7_75t_L g3067 ( 
.A(n_2581),
.Y(n_3067)
);

INVx8_ASAP7_75t_L g3068 ( 
.A(n_2603),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2624),
.B(n_2292),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2841),
.Y(n_3070)
);

INVx2_ASAP7_75t_SL g3071 ( 
.A(n_2581),
.Y(n_3071)
);

INVx4_ASAP7_75t_L g3072 ( 
.A(n_2615),
.Y(n_3072)
);

CKINVDCx20_ASAP7_75t_R g3073 ( 
.A(n_2813),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2886),
.B(n_2487),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2625),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2533),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2630),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2630),
.Y(n_3078)
);

INVx1_ASAP7_75t_SL g3079 ( 
.A(n_2537),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2744),
.B(n_2452),
.Y(n_3080)
);

INVxp33_ASAP7_75t_L g3081 ( 
.A(n_2573),
.Y(n_3081)
);

INVx3_ASAP7_75t_L g3082 ( 
.A(n_2533),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2634),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2841),
.Y(n_3084)
);

INVx3_ASAP7_75t_L g3085 ( 
.A(n_2542),
.Y(n_3085)
);

BUFx3_ASAP7_75t_L g3086 ( 
.A(n_2821),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2845),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_2700),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2634),
.Y(n_3089)
);

INVxp33_ASAP7_75t_SL g3090 ( 
.A(n_2662),
.Y(n_3090)
);

BUFx2_ASAP7_75t_L g3091 ( 
.A(n_2753),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2627),
.B(n_2326),
.Y(n_3092)
);

NAND2xp33_ASAP7_75t_L g3093 ( 
.A(n_2829),
.B(n_2452),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2786),
.A2(n_2365),
.B1(n_2393),
.B2(n_2310),
.Y(n_3094)
);

INVx2_ASAP7_75t_SL g3095 ( 
.A(n_2628),
.Y(n_3095)
);

AO22x2_ASAP7_75t_L g3096 ( 
.A1(n_2879),
.A2(n_2194),
.B1(n_2088),
.B2(n_2499),
.Y(n_3096)
);

INVx5_ASAP7_75t_L g3097 ( 
.A(n_2835),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2845),
.Y(n_3098)
);

BUFx3_ASAP7_75t_L g3099 ( 
.A(n_2803),
.Y(n_3099)
);

INVx2_ASAP7_75t_SL g3100 ( 
.A(n_2628),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2635),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2846),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2613),
.B(n_2396),
.Y(n_3103)
);

BUFx2_ASAP7_75t_L g3104 ( 
.A(n_2753),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2846),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2858),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2858),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2862),
.Y(n_3108)
);

CKINVDCx6p67_ASAP7_75t_R g3109 ( 
.A(n_2549),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2602),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2635),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_2700),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_2619),
.B(n_2506),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2644),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2627),
.B(n_2346),
.Y(n_3115)
);

OAI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2838),
.A2(n_2479),
.B1(n_2486),
.B2(n_2470),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2862),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2631),
.B(n_2106),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2803),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2868),
.Y(n_3120)
);

INVx2_ASAP7_75t_SL g3121 ( 
.A(n_2934),
.Y(n_3121)
);

BUFx10_ASAP7_75t_L g3122 ( 
.A(n_2869),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_2835),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2644),
.Y(n_3124)
);

CKINVDCx20_ASAP7_75t_R g3125 ( 
.A(n_2586),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2868),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2880),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_2596),
.B(n_2487),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2647),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2601),
.B(n_2487),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2880),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2647),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2881),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2656),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2881),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_2835),
.Y(n_3136)
);

NOR3xp33_ASAP7_75t_L g3137 ( 
.A(n_2834),
.B(n_2430),
.C(n_2412),
.Y(n_3137)
);

CKINVDCx20_ASAP7_75t_R g3138 ( 
.A(n_2586),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2631),
.B(n_2361),
.Y(n_3139)
);

HB1xp67_ASAP7_75t_L g3140 ( 
.A(n_2740),
.Y(n_3140)
);

BUFx10_ASAP7_75t_L g3141 ( 
.A(n_2908),
.Y(n_3141)
);

INVx3_ASAP7_75t_L g3142 ( 
.A(n_2542),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2656),
.Y(n_3143)
);

INVx2_ASAP7_75t_SL g3144 ( 
.A(n_2934),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2847),
.Y(n_3145)
);

BUFx4f_ASAP7_75t_L g3146 ( 
.A(n_2742),
.Y(n_3146)
);

INVx4_ASAP7_75t_L g3147 ( 
.A(n_2615),
.Y(n_3147)
);

NAND2x1p5_ASAP7_75t_L g3148 ( 
.A(n_2835),
.B(n_2198),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2632),
.B(n_2638),
.Y(n_3149)
);

INVxp33_ASAP7_75t_SL g3150 ( 
.A(n_2697),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2744),
.B(n_2462),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2847),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2659),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2659),
.Y(n_3154)
);

OAI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2750),
.A2(n_2470),
.B1(n_2486),
.B2(n_2479),
.Y(n_3155)
);

AND3x2_ASAP7_75t_L g3156 ( 
.A(n_2761),
.B(n_2496),
.C(n_2336),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2848),
.Y(n_3157)
);

BUFx6f_ASAP7_75t_SL g3158 ( 
.A(n_2549),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2660),
.B(n_2462),
.Y(n_3159)
);

OAI22x1_ASAP7_75t_L g3160 ( 
.A1(n_2797),
.A2(n_2353),
.B1(n_2328),
.B2(n_2108),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2670),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2848),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2670),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2671),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2632),
.B(n_2358),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_2835),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2671),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_2660),
.B(n_2462),
.Y(n_3168)
);

INVx2_ASAP7_75t_SL g3169 ( 
.A(n_2948),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2850),
.Y(n_3170)
);

INVx2_ASAP7_75t_SL g3171 ( 
.A(n_2948),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2850),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2851),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2851),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2864),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2864),
.Y(n_3176)
);

INVx4_ASAP7_75t_L g3177 ( 
.A(n_2615),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2871),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2871),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2878),
.Y(n_3180)
);

INVx1_ASAP7_75t_SL g3181 ( 
.A(n_2740),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2878),
.Y(n_3182)
);

AOI21x1_ASAP7_75t_L g3183 ( 
.A1(n_2552),
.A2(n_2380),
.B(n_2371),
.Y(n_3183)
);

BUFx10_ASAP7_75t_L g3184 ( 
.A(n_2804),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2638),
.B(n_2310),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2884),
.Y(n_3186)
);

AOI21x1_ASAP7_75t_L g3187 ( 
.A1(n_2552),
.A2(n_2380),
.B(n_2371),
.Y(n_3187)
);

INVx2_ASAP7_75t_SL g3188 ( 
.A(n_2958),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_L g3189 ( 
.A(n_2661),
.B(n_2487),
.Y(n_3189)
);

INVx1_ASAP7_75t_SL g3190 ( 
.A(n_2761),
.Y(n_3190)
);

INVx2_ASAP7_75t_SL g3191 ( 
.A(n_2958),
.Y(n_3191)
);

BUFx3_ASAP7_75t_L g3192 ( 
.A(n_2803),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_2661),
.B(n_2462),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_2684),
.B(n_2462),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2884),
.Y(n_3195)
);

INVx4_ASAP7_75t_L g3196 ( 
.A(n_2640),
.Y(n_3196)
);

OR2x6_ASAP7_75t_L g3197 ( 
.A(n_2664),
.B(n_2419),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2885),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2809),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2885),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2569),
.Y(n_3201)
);

INVx3_ASAP7_75t_L g3202 ( 
.A(n_2542),
.Y(n_3202)
);

XOR2x2_ASAP7_75t_SL g3203 ( 
.A(n_2826),
.B(n_2328),
.Y(n_3203)
);

AOI22x1_ASAP7_75t_L g3204 ( 
.A1(n_2605),
.A2(n_2310),
.B1(n_2202),
.B2(n_2205),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_2557),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_2886),
.B(n_2127),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_2684),
.B(n_2476),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2557),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2693),
.B(n_2476),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2809),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2559),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2542),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2639),
.B(n_2385),
.Y(n_3213)
);

CKINVDCx6p67_ASAP7_75t_R g3214 ( 
.A(n_2637),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2569),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2639),
.B(n_2399),
.Y(n_3216)
);

OAI22xp33_ASAP7_75t_SL g3217 ( 
.A1(n_2641),
.A2(n_991),
.B1(n_1024),
.B2(n_857),
.Y(n_3217)
);

INVxp67_ASAP7_75t_SL g3218 ( 
.A(n_2640),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2693),
.B(n_2495),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_2579),
.B(n_2476),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2579),
.B(n_2495),
.Y(n_3221)
);

CKINVDCx6p67_ASAP7_75t_R g3222 ( 
.A(n_2754),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2570),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2570),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2571),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2641),
.B(n_2201),
.Y(n_3226)
);

AOI21x1_ASAP7_75t_L g3227 ( 
.A1(n_2566),
.A2(n_2391),
.B(n_2383),
.Y(n_3227)
);

AND2x2_ASAP7_75t_SL g3228 ( 
.A(n_2798),
.B(n_2157),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2571),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_2916),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2574),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_2856),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2559),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2574),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_2664),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2576),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2576),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2642),
.B(n_2201),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2568),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2568),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2580),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2578),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2542),
.Y(n_3243)
);

BUFx2_ASAP7_75t_L g3244 ( 
.A(n_2683),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2580),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2582),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2582),
.Y(n_3247)
);

OR2x2_ASAP7_75t_L g3248 ( 
.A(n_2779),
.B(n_2102),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2583),
.Y(n_3249)
);

INVx3_ASAP7_75t_L g3250 ( 
.A(n_2548),
.Y(n_3250)
);

BUFx8_ASAP7_75t_SL g3251 ( 
.A(n_2823),
.Y(n_3251)
);

NAND2xp33_ASAP7_75t_L g3252 ( 
.A(n_2856),
.B(n_2476),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2887),
.B(n_2495),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_2548),
.Y(n_3254)
);

INVx4_ASAP7_75t_L g3255 ( 
.A(n_2640),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2578),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2583),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_2823),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2588),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_2856),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2587),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2588),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_2598),
.B(n_2476),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2642),
.B(n_2202),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_2786),
.A2(n_2393),
.B1(n_2205),
.B2(n_2235),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2587),
.Y(n_3266)
);

OR2x6_ASAP7_75t_L g3267 ( 
.A(n_2856),
.B(n_2419),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2645),
.B(n_2233),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_2590),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2590),
.Y(n_3270)
);

AOI22x1_ASAP7_75t_L g3271 ( 
.A1(n_2605),
.A2(n_2612),
.B1(n_2525),
.B2(n_2524),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_2799),
.A2(n_2393),
.B1(n_2233),
.B2(n_2237),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2589),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_L g3274 ( 
.A(n_2598),
.B(n_2498),
.Y(n_3274)
);

CKINVDCx16_ASAP7_75t_R g3275 ( 
.A(n_2931),
.Y(n_3275)
);

NAND2xp33_ASAP7_75t_SL g3276 ( 
.A(n_2766),
.B(n_2477),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2589),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_2916),
.Y(n_3278)
);

INVx4_ASAP7_75t_L g3279 ( 
.A(n_2640),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2595),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2591),
.Y(n_3281)
);

NOR2x1p5_ASAP7_75t_L g3282 ( 
.A(n_2611),
.B(n_2519),
.Y(n_3282)
);

NAND2xp33_ASAP7_75t_SL g3283 ( 
.A(n_2773),
.B(n_2477),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2591),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_SL g3285 ( 
.A(n_2618),
.B(n_2477),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2645),
.B(n_2235),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2592),
.Y(n_3287)
);

INVx4_ASAP7_75t_L g3288 ( 
.A(n_2640),
.Y(n_3288)
);

AND3x2_ASAP7_75t_L g3289 ( 
.A(n_2962),
.B(n_2496),
.C(n_2197),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2592),
.Y(n_3290)
);

AND2x6_ASAP7_75t_L g3291 ( 
.A(n_2798),
.B(n_2416),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2595),
.Y(n_3292)
);

NAND2xp33_ASAP7_75t_L g3293 ( 
.A(n_2856),
.B(n_2477),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2599),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2795),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2795),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_2618),
.B(n_2477),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2831),
.Y(n_3298)
);

INVx5_ASAP7_75t_L g3299 ( 
.A(n_2870),
.Y(n_3299)
);

AO21x2_ASAP7_75t_L g3300 ( 
.A1(n_2806),
.A2(n_2391),
.B(n_2383),
.Y(n_3300)
);

INVx2_ASAP7_75t_SL g3301 ( 
.A(n_2919),
.Y(n_3301)
);

AOI21x1_ASAP7_75t_L g3302 ( 
.A1(n_2566),
.A2(n_2398),
.B(n_2392),
.Y(n_3302)
);

NAND3xp33_ASAP7_75t_L g3303 ( 
.A(n_2646),
.B(n_2458),
.C(n_2246),
.Y(n_3303)
);

INVx5_ASAP7_75t_L g3304 ( 
.A(n_2870),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_2636),
.B(n_2498),
.Y(n_3305)
);

NAND2xp33_ASAP7_75t_L g3306 ( 
.A(n_2870),
.B(n_2485),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_2599),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_2636),
.B(n_2498),
.Y(n_3308)
);

INVxp33_ASAP7_75t_L g3309 ( 
.A(n_2584),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_2742),
.Y(n_3310)
);

OR2x2_ASAP7_75t_L g3311 ( 
.A(n_2688),
.B(n_2518),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_2526),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_2782),
.B(n_2485),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2526),
.Y(n_3314)
);

AND3x2_ASAP7_75t_L g3315 ( 
.A(n_2827),
.B(n_2197),
.C(n_2268),
.Y(n_3315)
);

BUFx6f_ASAP7_75t_L g3316 ( 
.A(n_2870),
.Y(n_3316)
);

BUFx6f_ASAP7_75t_L g3317 ( 
.A(n_2870),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2530),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_2919),
.Y(n_3319)
);

AOI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_2799),
.A2(n_2393),
.B1(n_2237),
.B2(n_2249),
.Y(n_3320)
);

NAND2xp33_ASAP7_75t_SL g3321 ( 
.A(n_2788),
.B(n_2485),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2831),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2646),
.B(n_2246),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2855),
.B(n_2485),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2650),
.B(n_2249),
.Y(n_3325)
);

AND2x4_ASAP7_75t_L g3326 ( 
.A(n_2561),
.B(n_2422),
.Y(n_3326)
);

INVxp67_ASAP7_75t_SL g3327 ( 
.A(n_2653),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2530),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2832),
.Y(n_3329)
);

INVx2_ASAP7_75t_SL g3330 ( 
.A(n_2859),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2531),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2898),
.B(n_2502),
.Y(n_3332)
);

INVxp33_ASAP7_75t_L g3333 ( 
.A(n_2648),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_2531),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_2629),
.B(n_2502),
.Y(n_3335)
);

INVx1_ASAP7_75t_SL g3336 ( 
.A(n_2827),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_2561),
.B(n_2422),
.Y(n_3337)
);

BUFx10_ASAP7_75t_L g3338 ( 
.A(n_2883),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_R g3339 ( 
.A(n_2861),
.B(n_2090),
.Y(n_3339)
);

INVx3_ASAP7_75t_L g3340 ( 
.A(n_2548),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2540),
.Y(n_3341)
);

INVx2_ASAP7_75t_SL g3342 ( 
.A(n_2859),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_2643),
.B(n_2485),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_2887),
.B(n_2502),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_2649),
.B(n_2488),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2685),
.B(n_2442),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2650),
.B(n_2652),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2540),
.Y(n_3348)
);

BUFx3_ASAP7_75t_L g3349 ( 
.A(n_2742),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_2888),
.A2(n_2250),
.B1(n_2257),
.B2(n_2254),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_2883),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_2691),
.B(n_2488),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_2902),
.A2(n_2250),
.B1(n_2257),
.B2(n_2254),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2832),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2728),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2728),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2730),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2554),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2554),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_2902),
.A2(n_2974),
.B1(n_2976),
.B2(n_2972),
.Y(n_3360)
);

INVx3_ASAP7_75t_L g3361 ( 
.A(n_2548),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2652),
.B(n_2318),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2730),
.Y(n_3363)
);

INVx8_ASAP7_75t_L g3364 ( 
.A(n_2603),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_2842),
.B(n_2488),
.Y(n_3365)
);

INVx3_ASAP7_75t_L g3366 ( 
.A(n_2548),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_2903),
.A2(n_2320),
.B1(n_2331),
.B2(n_2318),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_2883),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_2733),
.Y(n_3369)
);

INVx4_ASAP7_75t_L g3370 ( 
.A(n_2653),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2733),
.Y(n_3371)
);

INVx5_ASAP7_75t_L g3372 ( 
.A(n_2883),
.Y(n_3372)
);

INVx5_ASAP7_75t_L g3373 ( 
.A(n_2890),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2751),
.Y(n_3374)
);

AO21x2_ASAP7_75t_L g3375 ( 
.A1(n_2806),
.A2(n_2398),
.B(n_2392),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2751),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_SL g3377 ( 
.A(n_2692),
.B(n_2488),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_2694),
.B(n_2488),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2763),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_2763),
.Y(n_3380)
);

OR2x6_ASAP7_75t_L g3381 ( 
.A(n_2890),
.B(n_2419),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_2742),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2765),
.Y(n_3383)
);

CKINVDCx5p33_ASAP7_75t_R g3384 ( 
.A(n_2861),
.Y(n_3384)
);

OAI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_2654),
.A2(n_2492),
.B1(n_2449),
.B2(n_2465),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_2654),
.B(n_2320),
.Y(n_3386)
);

BUFx6f_ASAP7_75t_L g3387 ( 
.A(n_2890),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2765),
.Y(n_3388)
);

INVx4_ASAP7_75t_L g3389 ( 
.A(n_2653),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2767),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2767),
.Y(n_3391)
);

INVx2_ASAP7_75t_SL g3392 ( 
.A(n_2859),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2768),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2768),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2781),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2781),
.Y(n_3396)
);

INVx1_ASAP7_75t_SL g3397 ( 
.A(n_2877),
.Y(n_3397)
);

NAND2xp33_ASAP7_75t_SL g3398 ( 
.A(n_2695),
.B(n_2492),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_2783),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_2890),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2783),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2655),
.B(n_2331),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2791),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2791),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_2890),
.Y(n_3405)
);

INVx3_ASAP7_75t_L g3406 ( 
.A(n_2899),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_2538),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2802),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_L g3409 ( 
.A1(n_2903),
.A2(n_2334),
.B1(n_2337),
.B2(n_2335),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2802),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_2699),
.B(n_2492),
.Y(n_3411)
);

INVx1_ASAP7_75t_SL g3412 ( 
.A(n_2877),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_2538),
.Y(n_3413)
);

INVx2_ASAP7_75t_SL g3414 ( 
.A(n_2872),
.Y(n_3414)
);

NAND3xp33_ASAP7_75t_L g3415 ( 
.A(n_2655),
.B(n_2335),
.C(n_2334),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_2539),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_2752),
.B(n_2492),
.Y(n_3417)
);

AO21x2_ASAP7_75t_L g3418 ( 
.A1(n_2807),
.A2(n_2403),
.B(n_2400),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2663),
.B(n_2337),
.Y(n_3419)
);

AOI21x1_ASAP7_75t_L g3420 ( 
.A1(n_2593),
.A2(n_2403),
.B(n_2400),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_2899),
.Y(n_3421)
);

INVx4_ASAP7_75t_L g3422 ( 
.A(n_2653),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_2762),
.B(n_2492),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2663),
.B(n_2347),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_2539),
.Y(n_3425)
);

BUFx4f_ASAP7_75t_L g3426 ( 
.A(n_2742),
.Y(n_3426)
);

BUFx3_ASAP7_75t_L g3427 ( 
.A(n_2745),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_2872),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_2541),
.Y(n_3429)
);

OAI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_2665),
.A2(n_2973),
.B1(n_2968),
.B2(n_2669),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2665),
.B(n_2347),
.Y(n_3431)
);

INVx1_ASAP7_75t_SL g3432 ( 
.A(n_2882),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2541),
.Y(n_3433)
);

AND2x6_ASAP7_75t_L g3434 ( 
.A(n_2807),
.B(n_2423),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_L g3435 ( 
.A(n_2770),
.B(n_2442),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_SL g3436 ( 
.A(n_2745),
.B(n_2423),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_2668),
.B(n_2354),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2546),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_2668),
.B(n_2426),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2810),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_2546),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_2745),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_2547),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_2606),
.B(n_2449),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_2547),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_2932),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_2932),
.Y(n_3447)
);

AOI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_2669),
.A2(n_2354),
.B1(n_2359),
.B2(n_2357),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_2672),
.B(n_2426),
.Y(n_3449)
);

BUFx6f_ASAP7_75t_L g3450 ( 
.A(n_2899),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_2932),
.Y(n_3451)
);

INVxp67_ASAP7_75t_L g3452 ( 
.A(n_2882),
.Y(n_3452)
);

CKINVDCx20_ASAP7_75t_R g3453 ( 
.A(n_2721),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3298),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3172),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3206),
.B(n_2465),
.Y(n_3456)
);

CKINVDCx16_ASAP7_75t_R g3457 ( 
.A(n_3339),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_2979),
.B(n_2099),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3298),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3011),
.A2(n_3115),
.B(n_3092),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3322),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_3099),
.B(n_2701),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3021),
.B(n_2672),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3322),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3206),
.B(n_2467),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_2986),
.B(n_2223),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_3099),
.B(n_2920),
.Y(n_3467)
);

NAND2x1p5_ASAP7_75t_L g3468 ( 
.A(n_3146),
.B(n_2745),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3329),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3219),
.B(n_2467),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3009),
.B(n_2251),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3030),
.B(n_2677),
.Y(n_3472)
);

INVxp67_ASAP7_75t_SL g3473 ( 
.A(n_3205),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3329),
.Y(n_3474)
);

BUFx3_ASAP7_75t_L g3475 ( 
.A(n_3091),
.Y(n_3475)
);

NOR2xp33_ASAP7_75t_L g3476 ( 
.A(n_3033),
.B(n_2266),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3354),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3221),
.B(n_3274),
.Y(n_3478)
);

INVx4_ASAP7_75t_L g3479 ( 
.A(n_3047),
.Y(n_3479)
);

CKINVDCx20_ASAP7_75t_R g3480 ( 
.A(n_3073),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3354),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_3305),
.B(n_3308),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_3099),
.B(n_2920),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3049),
.B(n_2332),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2980),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_2980),
.Y(n_3486)
);

INVxp67_ASAP7_75t_L g3487 ( 
.A(n_3140),
.Y(n_3487)
);

AND2x2_ASAP7_75t_SL g3488 ( 
.A(n_3137),
.B(n_3010),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3172),
.Y(n_3489)
);

NAND2xp33_ASAP7_75t_SL g3490 ( 
.A(n_3026),
.B(n_2423),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3103),
.B(n_2421),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3119),
.B(n_2920),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_2990),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3248),
.B(n_2312),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2990),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3248),
.B(n_2461),
.Y(n_3496)
);

XOR2xp5_ASAP7_75t_L g3497 ( 
.A(n_3010),
.B(n_1829),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3175),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_2996),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_2996),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3008),
.Y(n_3501)
);

CKINVDCx5p33_ASAP7_75t_R g3502 ( 
.A(n_3251),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3008),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3012),
.Y(n_3504)
);

XOR2xp5_ASAP7_75t_L g3505 ( 
.A(n_3060),
.B(n_1833),
.Y(n_3505)
);

BUFx8_ASAP7_75t_L g3506 ( 
.A(n_3158),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_3119),
.B(n_2545),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3012),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3023),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3128),
.B(n_2421),
.Y(n_3510)
);

INVxp33_ASAP7_75t_L g3511 ( 
.A(n_3062),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3023),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_2989),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3027),
.Y(n_3514)
);

INVx1_ASAP7_75t_SL g3515 ( 
.A(n_3036),
.Y(n_3515)
);

BUFx2_ASAP7_75t_L g3516 ( 
.A(n_3091),
.Y(n_3516)
);

NAND2xp33_ASAP7_75t_SL g3517 ( 
.A(n_3026),
.B(n_2423),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3027),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3029),
.Y(n_3519)
);

INVx2_ASAP7_75t_SL g3520 ( 
.A(n_3104),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3029),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3031),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3031),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3335),
.B(n_2426),
.Y(n_3524)
);

OR2x6_ASAP7_75t_L g3525 ( 
.A(n_3197),
.B(n_2425),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3121),
.B(n_2497),
.Y(n_3526)
);

OAI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3016),
.A2(n_2719),
.B(n_2681),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_SL g3528 ( 
.A(n_3228),
.B(n_2459),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3175),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3034),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3034),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3042),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3042),
.Y(n_3533)
);

XNOR2x2_ASAP7_75t_L g3534 ( 
.A(n_3160),
.B(n_2228),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3050),
.Y(n_3535)
);

INVxp33_ASAP7_75t_SL g3536 ( 
.A(n_2995),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3050),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_2989),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3058),
.Y(n_3539)
);

INVx3_ASAP7_75t_R g3540 ( 
.A(n_3104),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3058),
.Y(n_3541)
);

HB1xp67_ASAP7_75t_L g3542 ( 
.A(n_3036),
.Y(n_3542)
);

BUFx6f_ASAP7_75t_L g3543 ( 
.A(n_2989),
.Y(n_3543)
);

BUFx6f_ASAP7_75t_L g3544 ( 
.A(n_2998),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3043),
.A2(n_2269),
.B(n_2198),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3121),
.B(n_2497),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3061),
.Y(n_3547)
);

INVxp33_ASAP7_75t_L g3548 ( 
.A(n_3067),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3061),
.Y(n_3549)
);

XNOR2xp5_ASAP7_75t_L g3550 ( 
.A(n_3125),
.B(n_1833),
.Y(n_3550)
);

BUFx8_ASAP7_75t_L g3551 ( 
.A(n_3158),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3070),
.Y(n_3552)
);

XOR2x2_ASAP7_75t_L g3553 ( 
.A(n_3203),
.B(n_2648),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3346),
.B(n_3435),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3070),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3084),
.Y(n_3556)
);

NAND2xp33_ASAP7_75t_SL g3557 ( 
.A(n_3158),
.B(n_2423),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3053),
.B(n_2677),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3084),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3069),
.B(n_2426),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3087),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3087),
.Y(n_3562)
);

XNOR2xp5_ASAP7_75t_L g3563 ( 
.A(n_3138),
.B(n_1834),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3098),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3098),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_L g3566 ( 
.A(n_3113),
.B(n_2429),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3102),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3102),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3105),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3105),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3106),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3176),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3189),
.B(n_2429),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3144),
.B(n_2497),
.Y(n_3574)
);

INVxp67_ASAP7_75t_SL g3575 ( 
.A(n_3205),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3106),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3165),
.B(n_3130),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3107),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_L g3579 ( 
.A(n_3444),
.B(n_2429),
.Y(n_3579)
);

CKINVDCx5p33_ASAP7_75t_R g3580 ( 
.A(n_2995),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3107),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3108),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3108),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3117),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3117),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3120),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3176),
.Y(n_3587)
);

BUFx6f_ASAP7_75t_L g3588 ( 
.A(n_2998),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3120),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3126),
.Y(n_3590)
);

NOR2xp67_ASAP7_75t_L g3591 ( 
.A(n_3258),
.B(n_2418),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3126),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2991),
.B(n_2678),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3127),
.Y(n_3594)
);

OR2x2_ASAP7_75t_L g3595 ( 
.A(n_3025),
.B(n_2268),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3127),
.Y(n_3596)
);

OR2x2_ASAP7_75t_L g3597 ( 
.A(n_3025),
.B(n_2279),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3131),
.Y(n_3598)
);

BUFx6f_ASAP7_75t_L g3599 ( 
.A(n_2998),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3131),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3133),
.Y(n_3601)
);

AND2x6_ASAP7_75t_L g3602 ( 
.A(n_3006),
.B(n_2604),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3119),
.B(n_2545),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3013),
.B(n_2434),
.Y(n_3604)
);

XNOR2x2_ASAP7_75t_L g3605 ( 
.A(n_3160),
.B(n_2228),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_3088),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3133),
.Y(n_3607)
);

INVx2_ASAP7_75t_SL g3608 ( 
.A(n_3199),
.Y(n_3608)
);

INVxp67_ASAP7_75t_SL g3609 ( 
.A(n_3208),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_L g3610 ( 
.A(n_3244),
.B(n_2429),
.Y(n_3610)
);

INVxp33_ASAP7_75t_SL g3611 ( 
.A(n_3088),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3135),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_3199),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3135),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3201),
.Y(n_3615)
);

XOR2xp5_ASAP7_75t_L g3616 ( 
.A(n_3060),
.B(n_1834),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3201),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3215),
.Y(n_3618)
);

XNOR2xp5_ASAP7_75t_L g3619 ( 
.A(n_3453),
.B(n_1849),
.Y(n_3619)
);

INVx1_ASAP7_75t_SL g3620 ( 
.A(n_3190),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3144),
.B(n_2678),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_SL g3622 ( 
.A(n_3228),
.B(n_2459),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3215),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3223),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3223),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3224),
.Y(n_3626)
);

CKINVDCx20_ASAP7_75t_R g3627 ( 
.A(n_3214),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3169),
.B(n_2679),
.Y(n_3628)
);

NOR2xp33_ASAP7_75t_L g3629 ( 
.A(n_3244),
.B(n_2445),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3224),
.Y(n_3630)
);

AOI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3183),
.A2(n_2525),
.B(n_2524),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3225),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3225),
.Y(n_3633)
);

INVx4_ASAP7_75t_L g3634 ( 
.A(n_3047),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3229),
.Y(n_3635)
);

XOR2xp5_ASAP7_75t_L g3636 ( 
.A(n_3112),
.B(n_1849),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3229),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3169),
.B(n_2679),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3231),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3231),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3171),
.B(n_2519),
.Y(n_3641)
);

NOR2xp67_ASAP7_75t_L g3642 ( 
.A(n_3258),
.B(n_2418),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3171),
.B(n_2519),
.Y(n_3643)
);

NOR2xp33_ASAP7_75t_SL g3644 ( 
.A(n_3228),
.B(n_2811),
.Y(n_3644)
);

NAND2xp33_ASAP7_75t_R g3645 ( 
.A(n_3150),
.B(n_2279),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3234),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3234),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3188),
.B(n_2680),
.Y(n_3648)
);

XOR2xp5_ASAP7_75t_L g3649 ( 
.A(n_3112),
.B(n_1851),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3236),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_2992),
.B(n_2445),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_3214),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3188),
.B(n_2453),
.Y(n_3653)
);

NAND2x1p5_ASAP7_75t_L g3654 ( 
.A(n_3146),
.B(n_2745),
.Y(n_3654)
);

AND2x6_ASAP7_75t_L g3655 ( 
.A(n_3006),
.B(n_2604),
.Y(n_3655)
);

OR2x2_ASAP7_75t_L g3656 ( 
.A(n_3181),
.B(n_2336),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3236),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3237),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3237),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3191),
.B(n_2680),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3191),
.B(n_2453),
.Y(n_3661)
);

OR2x2_ASAP7_75t_L g3662 ( 
.A(n_3079),
.B(n_2508),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_3040),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3182),
.Y(n_3664)
);

AND2x6_ASAP7_75t_L g3665 ( 
.A(n_3006),
.B(n_2608),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3017),
.B(n_2434),
.Y(n_3666)
);

CKINVDCx5p33_ASAP7_75t_R g3667 ( 
.A(n_3384),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3241),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3332),
.B(n_2456),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3241),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3245),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3245),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3246),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3246),
.Y(n_3674)
);

INVxp67_ASAP7_75t_SL g3675 ( 
.A(n_3208),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3247),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3247),
.Y(n_3677)
);

NAND2xp33_ASAP7_75t_R g3678 ( 
.A(n_3150),
.B(n_2897),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3249),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3249),
.Y(n_3680)
);

INVxp33_ASAP7_75t_L g3681 ( 
.A(n_3081),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3257),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3257),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3182),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3259),
.Y(n_3685)
);

CKINVDCx5p33_ASAP7_75t_R g3686 ( 
.A(n_3384),
.Y(n_3686)
);

INVxp67_ASAP7_75t_L g3687 ( 
.A(n_3056),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3186),
.Y(n_3688)
);

INVx2_ASAP7_75t_SL g3689 ( 
.A(n_3095),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3259),
.Y(n_3690)
);

INVxp33_ASAP7_75t_L g3691 ( 
.A(n_3309),
.Y(n_3691)
);

XOR2xp5_ASAP7_75t_L g3692 ( 
.A(n_3333),
.B(n_1851),
.Y(n_3692)
);

INVxp33_ASAP7_75t_L g3693 ( 
.A(n_3311),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3262),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3262),
.Y(n_3695)
);

CKINVDCx5p33_ASAP7_75t_R g3696 ( 
.A(n_3109),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3273),
.Y(n_3697)
);

XOR2xp5_ASAP7_75t_L g3698 ( 
.A(n_3275),
.B(n_1729),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3273),
.Y(n_3699)
);

CKINVDCx20_ASAP7_75t_R g3700 ( 
.A(n_3109),
.Y(n_3700)
);

AND2x2_ASAP7_75t_SL g3701 ( 
.A(n_3275),
.B(n_2434),
.Y(n_3701)
);

INVxp67_ASAP7_75t_SL g3702 ( 
.A(n_3211),
.Y(n_3702)
);

BUFx6f_ASAP7_75t_L g3703 ( 
.A(n_3040),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3277),
.Y(n_3704)
);

OAI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3016),
.A2(n_2988),
.B(n_3303),
.Y(n_3705)
);

OR2x2_ASAP7_75t_L g3706 ( 
.A(n_3079),
.B(n_2508),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3186),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_L g3708 ( 
.A(n_3452),
.B(n_2456),
.Y(n_3708)
);

XOR2x2_ASAP7_75t_L g3709 ( 
.A(n_3203),
.B(n_2797),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3277),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3281),
.Y(n_3711)
);

NAND2x1p5_ASAP7_75t_L g3712 ( 
.A(n_3146),
.B(n_2760),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3230),
.B(n_2457),
.Y(n_3713)
);

BUFx6f_ASAP7_75t_L g3714 ( 
.A(n_3040),
.Y(n_3714)
);

NAND2x1p5_ASAP7_75t_L g3715 ( 
.A(n_3426),
.B(n_2760),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3281),
.Y(n_3716)
);

NOR2xp33_ASAP7_75t_L g3717 ( 
.A(n_3336),
.B(n_2457),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3284),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3284),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3287),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3287),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3290),
.Y(n_3722)
);

XOR2x2_ASAP7_75t_L g3723 ( 
.A(n_3090),
.B(n_2697),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3290),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_3397),
.B(n_2463),
.Y(n_3725)
);

CKINVDCx5p33_ASAP7_75t_R g3726 ( 
.A(n_3222),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3195),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3295),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3295),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3195),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3296),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3230),
.B(n_2463),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_L g3733 ( 
.A(n_3412),
.B(n_2466),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3278),
.B(n_2466),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3296),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3095),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3408),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3408),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3410),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3410),
.Y(n_3740)
);

CKINVDCx5p33_ASAP7_75t_R g3741 ( 
.A(n_3222),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3210),
.Y(n_3742)
);

AND2x4_ASAP7_75t_L g3743 ( 
.A(n_3192),
.B(n_2545),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3440),
.Y(n_3744)
);

AND2x6_ASAP7_75t_L g3745 ( 
.A(n_3006),
.B(n_2608),
.Y(n_3745)
);

AND2x6_ASAP7_75t_L g3746 ( 
.A(n_3006),
.B(n_2610),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3440),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3145),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3363),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3278),
.B(n_2471),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3145),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_SL g3752 ( 
.A(n_3090),
.B(n_2811),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3301),
.B(n_2471),
.Y(n_3753)
);

CKINVDCx20_ASAP7_75t_R g3754 ( 
.A(n_3066),
.Y(n_3754)
);

CKINVDCx20_ASAP7_75t_R g3755 ( 
.A(n_3066),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3152),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3363),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3152),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3157),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3432),
.B(n_2473),
.Y(n_3760)
);

CKINVDCx5p33_ASAP7_75t_R g3761 ( 
.A(n_3066),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3157),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3162),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3162),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3170),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3170),
.Y(n_3766)
);

NOR2xp33_ASAP7_75t_L g3767 ( 
.A(n_3213),
.B(n_3216),
.Y(n_3767)
);

NOR2xp67_ASAP7_75t_L g3768 ( 
.A(n_3110),
.B(n_2418),
.Y(n_3768)
);

XOR2x2_ASAP7_75t_L g3769 ( 
.A(n_3156),
.B(n_2556),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_3235),
.B(n_2473),
.Y(n_3770)
);

INVx2_ASAP7_75t_SL g3771 ( 
.A(n_3100),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3301),
.B(n_2482),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3173),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3100),
.Y(n_3774)
);

INVxp67_ASAP7_75t_SL g3775 ( 
.A(n_3211),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3184),
.B(n_2482),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3235),
.B(n_2483),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3173),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3174),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3174),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_3093),
.A2(n_3293),
.B(n_3252),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3319),
.B(n_2483),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3178),
.Y(n_3783)
);

BUFx3_ASAP7_75t_L g3784 ( 
.A(n_3056),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3178),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3179),
.Y(n_3786)
);

NOR2xp33_ASAP7_75t_SL g3787 ( 
.A(n_3197),
.B(n_2854),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3369),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3179),
.Y(n_3789)
);

CKINVDCx20_ASAP7_75t_R g3790 ( 
.A(n_3066),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3180),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3180),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3198),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3198),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3200),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3200),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3369),
.Y(n_3797)
);

CKINVDCx5p33_ASAP7_75t_R g3798 ( 
.A(n_3122),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3355),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3319),
.B(n_3071),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3253),
.B(n_2505),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3355),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3356),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3356),
.Y(n_3804)
);

CKINVDCx20_ASAP7_75t_R g3805 ( 
.A(n_3122),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3357),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3253),
.B(n_2505),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_L g3808 ( 
.A(n_3071),
.B(n_2226),
.Y(n_3808)
);

AND2x4_ASAP7_75t_L g3809 ( 
.A(n_3192),
.B(n_2555),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3357),
.Y(n_3810)
);

XOR2x2_ASAP7_75t_L g3811 ( 
.A(n_3315),
.B(n_2556),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3371),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3192),
.B(n_2555),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3039),
.B(n_2682),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3311),
.B(n_2247),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3344),
.B(n_2434),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3374),
.Y(n_3817)
);

XNOR2xp5_ASAP7_75t_L g3818 ( 
.A(n_3289),
.B(n_2696),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3371),
.Y(n_3819)
);

XNOR2x2_ASAP7_75t_L g3820 ( 
.A(n_3096),
.B(n_2353),
.Y(n_3820)
);

INVxp33_ASAP7_75t_L g3821 ( 
.A(n_3365),
.Y(n_3821)
);

XOR2xp5_ASAP7_75t_L g3822 ( 
.A(n_3096),
.B(n_1729),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3041),
.B(n_2682),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3376),
.Y(n_3824)
);

XOR2xp5_ASAP7_75t_L g3825 ( 
.A(n_3096),
.B(n_1730),
.Y(n_3825)
);

INVx2_ASAP7_75t_SL g3826 ( 
.A(n_3110),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3184),
.B(n_2256),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3376),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3374),
.Y(n_3829)
);

XOR2xp5_ASAP7_75t_L g3830 ( 
.A(n_3096),
.B(n_1730),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3383),
.Y(n_3831)
);

XNOR2x2_ASAP7_75t_L g3832 ( 
.A(n_3080),
.B(n_2108),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3383),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3390),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3390),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3379),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3344),
.B(n_2434),
.Y(n_3837)
);

XNOR2xp5_ASAP7_75t_L g3838 ( 
.A(n_3055),
.B(n_2696),
.Y(n_3838)
);

INVxp67_ASAP7_75t_L g3839 ( 
.A(n_3365),
.Y(n_3839)
);

INVxp33_ASAP7_75t_L g3840 ( 
.A(n_3151),
.Y(n_3840)
);

BUFx6f_ASAP7_75t_L g3841 ( 
.A(n_3086),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3379),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3391),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3184),
.B(n_2435),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3391),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3380),
.Y(n_3846)
);

CKINVDCx20_ASAP7_75t_R g3847 ( 
.A(n_3122),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3393),
.Y(n_3848)
);

OAI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3303),
.A2(n_2719),
.B(n_2681),
.Y(n_3849)
);

CKINVDCx5p33_ASAP7_75t_R g3850 ( 
.A(n_3122),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3393),
.Y(n_3851)
);

OR2x2_ASAP7_75t_L g3852 ( 
.A(n_2994),
.B(n_2508),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3396),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3455),
.Y(n_3854)
);

AOI22xp5_ASAP7_75t_L g3855 ( 
.A1(n_3476),
.A2(n_2984),
.B1(n_3000),
.B2(n_2982),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_L g3856 ( 
.A(n_3554),
.B(n_3184),
.Y(n_3856)
);

NAND3xp33_ASAP7_75t_L g3857 ( 
.A(n_3554),
.B(n_2480),
.C(n_2523),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3482),
.B(n_3074),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_SL g3859 ( 
.A(n_3566),
.B(n_2435),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_3566),
.B(n_2435),
.Y(n_3860)
);

NOR3xp33_ASAP7_75t_L g3861 ( 
.A(n_3476),
.B(n_3168),
.C(n_3159),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_3669),
.B(n_3141),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_3669),
.B(n_3471),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3489),
.Y(n_3864)
);

INVxp67_ASAP7_75t_L g3865 ( 
.A(n_3542),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3494),
.B(n_2435),
.Y(n_3866)
);

BUFx6f_ASAP7_75t_L g3867 ( 
.A(n_3513),
.Y(n_3867)
);

NOR2xp33_ASAP7_75t_L g3868 ( 
.A(n_3471),
.B(n_1743),
.Y(n_3868)
);

O2A1O1Ixp5_ASAP7_75t_L g3869 ( 
.A1(n_3524),
.A2(n_3579),
.B(n_3604),
.C(n_3573),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3482),
.A2(n_3197),
.B1(n_3032),
.B2(n_3385),
.Y(n_3870)
);

OR2x6_ASAP7_75t_L g3871 ( 
.A(n_3525),
.B(n_3197),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3781),
.A2(n_3306),
.B(n_3426),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3767),
.B(n_3074),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3767),
.B(n_3439),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3478),
.B(n_3439),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3577),
.B(n_3449),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3491),
.B(n_3141),
.Y(n_3877)
);

NAND2xp33_ASAP7_75t_L g3878 ( 
.A(n_3577),
.B(n_2435),
.Y(n_3878)
);

INVx3_ASAP7_75t_L g3879 ( 
.A(n_3479),
.Y(n_3879)
);

INVx3_ASAP7_75t_L g3880 ( 
.A(n_3479),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3470),
.B(n_3449),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3460),
.B(n_3141),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3460),
.B(n_3141),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3524),
.B(n_3193),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_L g3885 ( 
.A(n_3458),
.B(n_3194),
.Y(n_3885)
);

AOI22xp33_ASAP7_75t_L g3886 ( 
.A1(n_3534),
.A2(n_3605),
.B1(n_3553),
.B2(n_3709),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3456),
.B(n_3207),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3484),
.B(n_2994),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3465),
.B(n_3209),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3498),
.Y(n_3890)
);

A2O1A1Ixp33_ASAP7_75t_L g3891 ( 
.A1(n_3579),
.A2(n_3002),
.B(n_3263),
.C(n_3220),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3513),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3615),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3472),
.B(n_3285),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_L g3895 ( 
.A(n_3458),
.B(n_3297),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3529),
.Y(n_3896)
);

INVx2_ASAP7_75t_SL g3897 ( 
.A(n_3475),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3472),
.B(n_3149),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3801),
.B(n_3347),
.Y(n_3899)
);

OAI22xp5_ASAP7_75t_L g3900 ( 
.A1(n_3560),
.A2(n_3197),
.B1(n_3047),
.B2(n_3046),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_L g3901 ( 
.A(n_3466),
.B(n_2997),
.Y(n_3901)
);

INVx2_ASAP7_75t_SL g3902 ( 
.A(n_3742),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3807),
.B(n_3496),
.Y(n_3903)
);

INVx3_ASAP7_75t_L g3904 ( 
.A(n_3634),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3494),
.B(n_2512),
.Y(n_3905)
);

AOI22xp5_ASAP7_75t_L g3906 ( 
.A1(n_3466),
.A2(n_2510),
.B1(n_2514),
.B2(n_2509),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3617),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3496),
.B(n_3326),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3572),
.Y(n_3909)
);

NOR2xp33_ASAP7_75t_L g3910 ( 
.A(n_3691),
.B(n_1743),
.Y(n_3910)
);

AND2x4_ASAP7_75t_L g3911 ( 
.A(n_3467),
.B(n_3483),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3560),
.B(n_3326),
.Y(n_3912)
);

INVx3_ASAP7_75t_L g3913 ( 
.A(n_3634),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3558),
.B(n_3326),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3558),
.B(n_3326),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3618),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3681),
.B(n_1744),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3623),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3624),
.Y(n_3919)
);

INVx4_ASAP7_75t_L g3920 ( 
.A(n_3513),
.Y(n_3920)
);

INVx4_ASAP7_75t_L g3921 ( 
.A(n_3538),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3587),
.Y(n_3922)
);

OR2x2_ASAP7_75t_L g3923 ( 
.A(n_3595),
.B(n_2509),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3625),
.Y(n_3924)
);

BUFx5_ASAP7_75t_L g3925 ( 
.A(n_3602),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3626),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3630),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3510),
.B(n_3337),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3620),
.B(n_1744),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3781),
.A2(n_3426),
.B(n_3345),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3664),
.Y(n_3931)
);

OAI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3573),
.A2(n_3047),
.B1(n_3046),
.B2(n_3267),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3632),
.Y(n_3933)
);

CKINVDCx5p33_ASAP7_75t_R g3934 ( 
.A(n_3480),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_L g3935 ( 
.A(n_3620),
.B(n_1757),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_3717),
.B(n_2512),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3684),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3463),
.B(n_3337),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_SL g3939 ( 
.A1(n_3820),
.A2(n_2370),
.B1(n_2375),
.B2(n_2394),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3463),
.B(n_3337),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3816),
.B(n_3337),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3717),
.B(n_2512),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_3725),
.B(n_2512),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3688),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3707),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3727),
.Y(n_3946)
);

A2O1A1Ixp33_ASAP7_75t_L g3947 ( 
.A1(n_3651),
.A2(n_3282),
.B(n_3352),
.C(n_3343),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_3725),
.B(n_2512),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3837),
.B(n_3139),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3653),
.B(n_2436),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3730),
.Y(n_3951)
);

AOI22xp5_ASAP7_75t_L g3952 ( 
.A1(n_3528),
.A2(n_2510),
.B1(n_2514),
.B2(n_2509),
.Y(n_3952)
);

BUFx6f_ASAP7_75t_SL g3953 ( 
.A(n_3784),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_3468),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3633),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3693),
.B(n_3815),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3661),
.B(n_3713),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_L g3958 ( 
.A(n_3511),
.B(n_1757),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3749),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3732),
.B(n_2436),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3757),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_3548),
.B(n_1767),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3733),
.B(n_2517),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3734),
.B(n_2438),
.Y(n_3964)
);

NAND2xp33_ASAP7_75t_L g3965 ( 
.A(n_3557),
.B(n_2517),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3750),
.B(n_2438),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3753),
.B(n_3772),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3635),
.Y(n_3968)
);

OR2x2_ASAP7_75t_L g3969 ( 
.A(n_3597),
.B(n_2510),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3821),
.B(n_2997),
.Y(n_3970)
);

OAI22xp33_ASAP7_75t_L g3971 ( 
.A1(n_3787),
.A2(n_2501),
.B1(n_2489),
.B2(n_2161),
.Y(n_3971)
);

AO22x1_ASAP7_75t_L g3972 ( 
.A1(n_3726),
.A2(n_2837),
.B1(n_2852),
.B2(n_2676),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3637),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3545),
.A2(n_3378),
.B(n_3377),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3782),
.B(n_2439),
.Y(n_3975)
);

INVx1_ASAP7_75t_SL g3976 ( 
.A(n_3515),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3815),
.B(n_2439),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3515),
.B(n_2261),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3814),
.B(n_2686),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3542),
.B(n_2283),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3639),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3788),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3814),
.B(n_3823),
.Y(n_3983)
);

INVxp67_ASAP7_75t_L g3984 ( 
.A(n_3662),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3545),
.A2(n_3417),
.B(n_3411),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3528),
.A2(n_2514),
.B1(n_2518),
.B2(n_2295),
.Y(n_3986)
);

O2A1O1Ixp33_ASAP7_75t_L g3987 ( 
.A1(n_3651),
.A2(n_3155),
.B(n_3116),
.C(n_3217),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3823),
.B(n_3526),
.Y(n_3988)
);

O2A1O1Ixp5_ASAP7_75t_L g3989 ( 
.A1(n_3666),
.A2(n_3423),
.B(n_3037),
.C(n_3436),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3832),
.A2(n_3217),
.B1(n_2686),
.B2(n_2698),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3733),
.B(n_2517),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3640),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3797),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3701),
.B(n_2420),
.Y(n_3994)
);

INVxp33_ASAP7_75t_L g3995 ( 
.A(n_3656),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3817),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3646),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3647),
.Y(n_3998)
);

NOR2xp33_ASAP7_75t_SL g3999 ( 
.A(n_3536),
.B(n_3611),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3760),
.B(n_2517),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3760),
.B(n_2517),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3650),
.Y(n_4002)
);

INVxp67_ASAP7_75t_SL g4003 ( 
.A(n_3473),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3657),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3488),
.A2(n_2687),
.B1(n_2702),
.B2(n_2698),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_3752),
.B(n_2428),
.Y(n_4006)
);

AOI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_3622),
.A2(n_2518),
.B1(n_1955),
.B2(n_2715),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3829),
.Y(n_4008)
);

AOI22xp33_ASAP7_75t_L g4009 ( 
.A1(n_3622),
.A2(n_2687),
.B1(n_2708),
.B2(n_2702),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3836),
.Y(n_4010)
);

INVx4_ASAP7_75t_L g4011 ( 
.A(n_3538),
.Y(n_4011)
);

INVxp33_ASAP7_75t_L g4012 ( 
.A(n_3550),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3658),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3546),
.B(n_3574),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3842),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3659),
.Y(n_4016)
);

NAND3xp33_ASAP7_75t_L g4017 ( 
.A(n_3776),
.B(n_2523),
.C(n_2431),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3839),
.B(n_2708),
.Y(n_4018)
);

INVxp67_ASAP7_75t_SL g4019 ( 
.A(n_3473),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3668),
.Y(n_4020)
);

BUFx6f_ASAP7_75t_L g4021 ( 
.A(n_3538),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3839),
.B(n_2709),
.Y(n_4022)
);

OAI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3610),
.A2(n_3047),
.B1(n_3046),
.B2(n_3267),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3670),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3641),
.B(n_2709),
.Y(n_4025)
);

OAI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3610),
.A2(n_3046),
.B1(n_3381),
.B2(n_3267),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_L g4027 ( 
.A(n_3643),
.B(n_2713),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3671),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3672),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3621),
.B(n_3628),
.Y(n_4030)
);

HB1xp67_ASAP7_75t_L g4031 ( 
.A(n_3516),
.Y(n_4031)
);

AOI22xp5_ASAP7_75t_L g4032 ( 
.A1(n_3645),
.A2(n_3678),
.B1(n_1955),
.B2(n_3827),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_SL g4033 ( 
.A(n_3520),
.B(n_2516),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3846),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3621),
.B(n_2713),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_SL g4036 ( 
.A(n_3608),
.B(n_2516),
.Y(n_4036)
);

NAND2x1p5_ASAP7_75t_L g4037 ( 
.A(n_3543),
.B(n_3442),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3673),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3613),
.B(n_2516),
.Y(n_4039)
);

OAI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3787),
.A2(n_2501),
.B1(n_2489),
.B2(n_2123),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3826),
.B(n_2516),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3674),
.Y(n_4042)
);

NOR2xp33_ASAP7_75t_L g4043 ( 
.A(n_3827),
.B(n_1767),
.Y(n_4043)
);

INVx2_ASAP7_75t_SL g4044 ( 
.A(n_3706),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_L g4045 ( 
.A(n_3487),
.B(n_2428),
.Y(n_4045)
);

NOR2xp67_ASAP7_75t_L g4046 ( 
.A(n_3667),
.B(n_2418),
.Y(n_4046)
);

INVx4_ASAP7_75t_L g4047 ( 
.A(n_3543),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_SL g4048 ( 
.A(n_3808),
.B(n_2516),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3770),
.B(n_2420),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3628),
.B(n_2714),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_3808),
.B(n_2431),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3638),
.B(n_2714),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3638),
.B(n_2716),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_L g4054 ( 
.A(n_3487),
.B(n_2432),
.Y(n_4054)
);

AOI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_3752),
.A2(n_2736),
.B1(n_2215),
.B2(n_2785),
.Y(n_4055)
);

AND2x4_ASAP7_75t_L g4056 ( 
.A(n_3467),
.B(n_3086),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3648),
.B(n_3660),
.Y(n_4057)
);

AND2x4_ASAP7_75t_L g4058 ( 
.A(n_3483),
.B(n_3086),
.Y(n_4058)
);

NOR2xp33_ASAP7_75t_L g4059 ( 
.A(n_3708),
.B(n_2432),
.Y(n_4059)
);

BUFx6f_ASAP7_75t_L g4060 ( 
.A(n_3543),
.Y(n_4060)
);

INVxp67_ASAP7_75t_L g4061 ( 
.A(n_3629),
.Y(n_4061)
);

INVx2_ASAP7_75t_SL g4062 ( 
.A(n_3689),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3676),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3677),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_SL g4065 ( 
.A1(n_3644),
.A2(n_2370),
.B1(n_2375),
.B2(n_2394),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3679),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3705),
.A2(n_2716),
.B1(n_2724),
.B2(n_2723),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3705),
.A2(n_2723),
.B1(n_2725),
.B2(n_2724),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3629),
.A2(n_2433),
.B1(n_2440),
.B2(n_2777),
.Y(n_4069)
);

BUFx5_ASAP7_75t_L g4070 ( 
.A(n_3602),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3648),
.B(n_3660),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3800),
.B(n_2725),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_L g4073 ( 
.A(n_3770),
.B(n_2433),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3680),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3777),
.B(n_3708),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3682),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_L g4077 ( 
.A(n_3777),
.B(n_2440),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3736),
.B(n_2897),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3800),
.B(n_3844),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3683),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3575),
.B(n_2727),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_SL g4082 ( 
.A(n_3771),
.B(n_2513),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3774),
.B(n_2513),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3575),
.B(n_2727),
.Y(n_4084)
);

INVxp67_ASAP7_75t_SL g4085 ( 
.A(n_3609),
.Y(n_4085)
);

O2A1O1Ixp33_ASAP7_75t_L g4086 ( 
.A1(n_3593),
.A2(n_3430),
.B(n_3118),
.C(n_2741),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_3609),
.A2(n_3046),
.B1(n_3267),
.B2(n_3381),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3685),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3675),
.B(n_2729),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3675),
.B(n_2729),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3702),
.B(n_2734),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_3457),
.B(n_3687),
.Y(n_4092)
);

INVxp67_ASAP7_75t_L g4093 ( 
.A(n_3852),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3702),
.B(n_2734),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3690),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_3687),
.B(n_2384),
.Y(n_4096)
);

OAI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3644),
.A2(n_2123),
.B1(n_2161),
.B2(n_2735),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3492),
.B(n_2513),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3694),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3695),
.Y(n_4100)
);

NOR3xp33_ASAP7_75t_L g4101 ( 
.A(n_3490),
.B(n_2351),
.C(n_2222),
.Y(n_4101)
);

INVx2_ASAP7_75t_SL g4102 ( 
.A(n_3741),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3697),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3692),
.B(n_2401),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3775),
.B(n_2735),
.Y(n_4105)
);

NAND2x1_ASAP7_75t_L g4106 ( 
.A(n_3602),
.B(n_3020),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3775),
.B(n_2737),
.Y(n_4107)
);

AOI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_3698),
.A2(n_3282),
.B1(n_2113),
.B2(n_2372),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3593),
.B(n_2737),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3492),
.B(n_2721),
.Y(n_4110)
);

CKINVDCx5p33_ASAP7_75t_R g4111 ( 
.A(n_3580),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3699),
.Y(n_4112)
);

NAND2xp33_ASAP7_75t_L g4113 ( 
.A(n_3602),
.B(n_3434),
.Y(n_4113)
);

NAND3xp33_ASAP7_75t_L g4114 ( 
.A(n_3563),
.B(n_2121),
.C(n_2129),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_3619),
.B(n_3497),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3462),
.B(n_2738),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3704),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3462),
.B(n_2738),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3507),
.B(n_2739),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3507),
.B(n_2129),
.Y(n_4120)
);

INVx3_ASAP7_75t_L g4121 ( 
.A(n_3468),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3840),
.B(n_2985),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3603),
.B(n_2739),
.Y(n_4123)
);

OR2x2_ASAP7_75t_L g4124 ( 
.A(n_3505),
.B(n_2503),
.Y(n_4124)
);

NOR2xp33_ASAP7_75t_L g4125 ( 
.A(n_3761),
.B(n_2255),
.Y(n_4125)
);

AOI221xp5_ASAP7_75t_L g4126 ( 
.A1(n_3822),
.A2(n_2490),
.B1(n_1194),
.B2(n_991),
.C(n_857),
.Y(n_4126)
);

AOI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_3754),
.A2(n_2241),
.B1(n_2910),
.B2(n_2124),
.Y(n_4127)
);

NOR2xp33_ASAP7_75t_L g4128 ( 
.A(n_3798),
.B(n_2255),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_3850),
.B(n_2503),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3710),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3603),
.B(n_2747),
.Y(n_4131)
);

OAI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_3849),
.A2(n_3415),
.B(n_2993),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_3711),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3743),
.B(n_2747),
.Y(n_4134)
);

INVx8_ASAP7_75t_L g4135 ( 
.A(n_3602),
.Y(n_4135)
);

NOR2xp33_ASAP7_75t_L g4136 ( 
.A(n_3636),
.B(n_2241),
.Y(n_4136)
);

BUFx6f_ASAP7_75t_L g4137 ( 
.A(n_3544),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3716),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_SL g4139 ( 
.A(n_3743),
.B(n_2985),
.Y(n_4139)
);

NOR2xp33_ASAP7_75t_L g4140 ( 
.A(n_3616),
.B(n_2824),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_L g4141 ( 
.A(n_3517),
.B(n_2183),
.C(n_2167),
.Y(n_4141)
);

CKINVDCx11_ASAP7_75t_R g4142 ( 
.A(n_3627),
.Y(n_4142)
);

NOR3xp33_ASAP7_75t_L g4143 ( 
.A(n_3809),
.B(n_2188),
.C(n_2585),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_3809),
.B(n_2985),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3813),
.B(n_2749),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3813),
.B(n_2749),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_SL g4147 ( 
.A(n_3652),
.B(n_2985),
.Y(n_4147)
);

INVx2_ASAP7_75t_SL g4148 ( 
.A(n_3686),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3718),
.B(n_2756),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3719),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_SL g4151 ( 
.A1(n_3825),
.A2(n_2900),
.B1(n_2490),
.B2(n_2444),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3720),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3721),
.Y(n_4153)
);

NOR2xp33_ASAP7_75t_L g4154 ( 
.A(n_3722),
.B(n_2874),
.Y(n_4154)
);

NOR3xp33_ASAP7_75t_L g4155 ( 
.A(n_3606),
.B(n_2444),
.C(n_2971),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3724),
.B(n_2756),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3728),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_3544),
.B(n_2910),
.Y(n_4158)
);

OAI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_3729),
.A2(n_3267),
.B1(n_3381),
.B2(n_3360),
.Y(n_4159)
);

OAI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_3731),
.A2(n_3381),
.B1(n_3064),
.B2(n_3272),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_3735),
.Y(n_4161)
);

NOR2xp67_ASAP7_75t_L g4162 ( 
.A(n_3696),
.B(n_2166),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3737),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3738),
.B(n_2757),
.Y(n_4164)
);

NOR2xp33_ASAP7_75t_SL g4165 ( 
.A(n_3502),
.B(n_2121),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3739),
.B(n_2757),
.Y(n_4166)
);

BUFx3_ASAP7_75t_L g4167 ( 
.A(n_3506),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_SL g4168 ( 
.A(n_3544),
.B(n_2760),
.Y(n_4168)
);

AND2x6_ASAP7_75t_SL g4169 ( 
.A(n_3525),
.B(n_2194),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3755),
.A2(n_3805),
.B1(n_3847),
.B2(n_3790),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3740),
.B(n_2758),
.Y(n_4171)
);

OR2x6_ASAP7_75t_L g4172 ( 
.A(n_3525),
.B(n_3381),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3744),
.B(n_2758),
.Y(n_4173)
);

NOR2xp33_ASAP7_75t_L g4174 ( 
.A(n_3747),
.B(n_2759),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3485),
.B(n_2759),
.Y(n_4175)
);

NOR3xp33_ASAP7_75t_L g4176 ( 
.A(n_3591),
.B(n_3324),
.C(n_3313),
.Y(n_4176)
);

BUFx6f_ASAP7_75t_L g4177 ( 
.A(n_3588),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_3527),
.A2(n_3048),
.B(n_2999),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_3527),
.A2(n_3048),
.B(n_2999),
.Y(n_4179)
);

AND2x4_ASAP7_75t_L g4180 ( 
.A(n_3588),
.B(n_3330),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3486),
.B(n_2769),
.Y(n_4181)
);

OR2x6_ASAP7_75t_L g4182 ( 
.A(n_3588),
.B(n_3044),
.Y(n_4182)
);

AND2x4_ASAP7_75t_L g4183 ( 
.A(n_3599),
.B(n_3330),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3493),
.B(n_2769),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3495),
.B(n_2772),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_L g4186 ( 
.A(n_3649),
.B(n_3540),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_3799),
.Y(n_4187)
);

AOI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_3849),
.A2(n_3048),
.B(n_2999),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_3599),
.B(n_3663),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_3599),
.B(n_2760),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3454),
.Y(n_4191)
);

NOR2xp33_ASAP7_75t_L g4192 ( 
.A(n_3830),
.B(n_2900),
.Y(n_4192)
);

INVx2_ASAP7_75t_L g4193 ( 
.A(n_3802),
.Y(n_4193)
);

INVx2_ASAP7_75t_SL g4194 ( 
.A(n_3663),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_3459),
.Y(n_4195)
);

AOI22xp5_ASAP7_75t_L g4196 ( 
.A1(n_3723),
.A2(n_3398),
.B1(n_3283),
.B2(n_3321),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3499),
.B(n_2772),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_3663),
.B(n_2760),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_3803),
.Y(n_4199)
);

BUFx6f_ASAP7_75t_L g4200 ( 
.A(n_3703),
.Y(n_4200)
);

NAND2xp33_ASAP7_75t_L g4201 ( 
.A(n_3655),
.B(n_3434),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3500),
.B(n_2775),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_3804),
.Y(n_4203)
);

INVxp67_ASAP7_75t_SL g4204 ( 
.A(n_3501),
.Y(n_4204)
);

NOR2xp33_ASAP7_75t_L g4205 ( 
.A(n_3703),
.B(n_2189),
.Y(n_4205)
);

NOR2xp33_ASAP7_75t_L g4206 ( 
.A(n_3703),
.B(n_2676),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3806),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3811),
.A2(n_3276),
.B1(n_3038),
.B2(n_2175),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_3714),
.B(n_2676),
.Y(n_4209)
);

BUFx6f_ASAP7_75t_SL g4210 ( 
.A(n_3714),
.Y(n_4210)
);

INVx2_ASAP7_75t_SL g4211 ( 
.A(n_3714),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_3810),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3841),
.B(n_3642),
.Y(n_4213)
);

INVx3_ASAP7_75t_L g4214 ( 
.A(n_3654),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3503),
.B(n_2775),
.Y(n_4215)
);

OAI22xp5_ASAP7_75t_L g4216 ( 
.A1(n_3504),
.A2(n_3265),
.B1(n_3007),
.B2(n_3342),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3812),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3508),
.B(n_2778),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3461),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3841),
.B(n_2764),
.Y(n_4220)
);

NAND3xp33_ASAP7_75t_L g4221 ( 
.A(n_3818),
.B(n_2121),
.C(n_2837),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_SL g4222 ( 
.A(n_3841),
.B(n_2764),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3768),
.B(n_2764),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_3509),
.B(n_2778),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_3838),
.B(n_2764),
.Y(n_4225)
);

AOI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_3769),
.A2(n_2175),
.B1(n_2121),
.B2(n_2837),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_3512),
.B(n_2780),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3514),
.B(n_2780),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_3819),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_3518),
.B(n_2789),
.Y(n_4230)
);

NOR2x2_ASAP7_75t_L g4231 ( 
.A(n_3871),
.B(n_2446),
.Y(n_4231)
);

INVx5_ASAP7_75t_L g4232 ( 
.A(n_4172),
.Y(n_4232)
);

BUFx3_ASAP7_75t_L g4233 ( 
.A(n_4111),
.Y(n_4233)
);

AND2x4_ASAP7_75t_SL g4234 ( 
.A(n_4056),
.B(n_3700),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3863),
.A2(n_3521),
.B1(n_3522),
.B2(n_3519),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_R g4236 ( 
.A(n_3934),
.B(n_3506),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3983),
.B(n_3523),
.Y(n_4237)
);

NOR2x1_ASAP7_75t_L g4238 ( 
.A(n_4017),
.B(n_2544),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3893),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_3863),
.B(n_4030),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4003),
.A2(n_3531),
.B1(n_3532),
.B2(n_3530),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4057),
.B(n_3533),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4071),
.B(n_3535),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_3886),
.A2(n_2852),
.B1(n_2872),
.B2(n_2558),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_3911),
.B(n_4056),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4042),
.Y(n_4246)
);

AND2x6_ASAP7_75t_SL g4247 ( 
.A(n_4192),
.B(n_2446),
.Y(n_4247)
);

INVx3_ASAP7_75t_L g4248 ( 
.A(n_3867),
.Y(n_4248)
);

AND2x6_ASAP7_75t_SL g4249 ( 
.A(n_4136),
.B(n_2852),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4063),
.Y(n_4250)
);

BUFx3_ASAP7_75t_L g4251 ( 
.A(n_3902),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_4059),
.B(n_2764),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4003),
.B(n_3537),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_3907),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4066),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_SL g4256 ( 
.A(n_3901),
.B(n_2787),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_4031),
.Y(n_4257)
);

NOR2xp33_ASAP7_75t_L g4258 ( 
.A(n_4043),
.B(n_2499),
.Y(n_4258)
);

HB1xp67_ASAP7_75t_L g4259 ( 
.A(n_4031),
.Y(n_4259)
);

NOR2x2_ASAP7_75t_L g4260 ( 
.A(n_3871),
.B(n_3407),
.Y(n_4260)
);

INVx5_ASAP7_75t_L g4261 ( 
.A(n_4172),
.Y(n_4261)
);

INVxp67_ASAP7_75t_SL g4262 ( 
.A(n_4019),
.Y(n_4262)
);

INVx2_ASAP7_75t_SL g4263 ( 
.A(n_4148),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3916),
.Y(n_4264)
);

BUFx2_ASAP7_75t_L g4265 ( 
.A(n_3897),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4019),
.B(n_3539),
.Y(n_4266)
);

BUFx3_ASAP7_75t_L g4267 ( 
.A(n_4102),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3901),
.B(n_2787),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3918),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4085),
.A2(n_3076),
.B(n_3065),
.Y(n_4270)
);

AND2x4_ASAP7_75t_L g4271 ( 
.A(n_3911),
.B(n_3310),
.Y(n_4271)
);

HB1xp67_ASAP7_75t_L g4272 ( 
.A(n_3976),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4076),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4085),
.B(n_3541),
.Y(n_4274)
);

AND2x4_ASAP7_75t_L g4275 ( 
.A(n_4058),
.B(n_3310),
.Y(n_4275)
);

AOI22xp33_ASAP7_75t_L g4276 ( 
.A1(n_3886),
.A2(n_2558),
.B1(n_2600),
.B2(n_2555),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_L g4277 ( 
.A(n_3868),
.B(n_3551),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_3898),
.B(n_3547),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3858),
.B(n_3549),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_3919),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4058),
.B(n_3310),
.Y(n_4281)
);

AND2x4_ASAP7_75t_L g4282 ( 
.A(n_4122),
.B(n_3349),
.Y(n_4282)
);

INVx4_ASAP7_75t_L g4283 ( 
.A(n_4210),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3873),
.B(n_3552),
.Y(n_4284)
);

INVx3_ASAP7_75t_L g4285 ( 
.A(n_3867),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_4073),
.B(n_4077),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4088),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_3924),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_3926),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_3874),
.B(n_3555),
.Y(n_4290)
);

AND2x4_ASAP7_75t_L g4291 ( 
.A(n_4172),
.B(n_4194),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_3867),
.Y(n_4292)
);

INVx3_ASAP7_75t_L g4293 ( 
.A(n_3892),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_3892),
.Y(n_4294)
);

BUFx6f_ASAP7_75t_L g4295 ( 
.A(n_3892),
.Y(n_4295)
);

AOI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_4006),
.A2(n_2771),
.B1(n_2600),
.B2(n_2622),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_R g4297 ( 
.A(n_3999),
.B(n_3551),
.Y(n_4297)
);

AOI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_4006),
.A2(n_2600),
.B1(n_2622),
.B2(n_2558),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_3903),
.B(n_3876),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_3869),
.A2(n_3415),
.B(n_3185),
.Y(n_4300)
);

NAND2x1p5_ASAP7_75t_L g4301 ( 
.A(n_4106),
.B(n_3349),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_4073),
.B(n_2787),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4095),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_3979),
.B(n_3556),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3927),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3933),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_3885),
.B(n_2789),
.Y(n_4307)
);

BUFx2_ASAP7_75t_L g4308 ( 
.A(n_3888),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3955),
.Y(n_4309)
);

NAND2xp33_ASAP7_75t_SL g4310 ( 
.A(n_3953),
.B(n_3123),
.Y(n_4310)
);

BUFx3_ASAP7_75t_L g4311 ( 
.A(n_4021),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4109),
.B(n_3559),
.Y(n_4312)
);

BUFx6f_ASAP7_75t_L g4313 ( 
.A(n_4021),
.Y(n_4313)
);

BUFx3_ASAP7_75t_L g4314 ( 
.A(n_4021),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_R g4315 ( 
.A(n_4165),
.B(n_2182),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3968),
.Y(n_4316)
);

INVx4_ASAP7_75t_L g4317 ( 
.A(n_4210),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_4099),
.Y(n_4318)
);

HB1xp67_ASAP7_75t_L g4319 ( 
.A(n_4044),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_3988),
.B(n_3561),
.Y(n_4320)
);

BUFx3_ASAP7_75t_L g4321 ( 
.A(n_4060),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_3865),
.Y(n_4322)
);

AND2x2_ASAP7_75t_SL g4323 ( 
.A(n_3965),
.B(n_2389),
.Y(n_4323)
);

AOI22x1_ASAP7_75t_L g4324 ( 
.A1(n_4204),
.A2(n_2790),
.B1(n_2893),
.B2(n_2792),
.Y(n_4324)
);

HB1xp67_ASAP7_75t_L g4325 ( 
.A(n_3865),
.Y(n_4325)
);

INVx5_ASAP7_75t_L g4326 ( 
.A(n_3871),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3973),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_3981),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_3862),
.B(n_3562),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4117),
.Y(n_4330)
);

INVx2_ASAP7_75t_SL g4331 ( 
.A(n_4062),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_3992),
.Y(n_4332)
);

INVxp67_ASAP7_75t_SL g4333 ( 
.A(n_4204),
.Y(n_4333)
);

INVx3_ASAP7_75t_L g4334 ( 
.A(n_4060),
.Y(n_4334)
);

AND2x4_ASAP7_75t_L g4335 ( 
.A(n_4211),
.B(n_4180),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4133),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3862),
.B(n_3564),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4138),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_SL g4339 ( 
.A(n_4077),
.B(n_2787),
.Y(n_4339)
);

BUFx3_ASAP7_75t_L g4340 ( 
.A(n_4060),
.Y(n_4340)
);

NOR2x1_ASAP7_75t_L g4341 ( 
.A(n_4046),
.B(n_4045),
.Y(n_4341)
);

BUFx3_ASAP7_75t_L g4342 ( 
.A(n_4137),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4150),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_SL g4344 ( 
.A(n_3885),
.B(n_2787),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_3895),
.B(n_3977),
.Y(n_4345)
);

NOR3xp33_ASAP7_75t_SL g4346 ( 
.A(n_4221),
.B(n_975),
.C(n_974),
.Y(n_4346)
);

INVxp67_ASAP7_75t_L g4347 ( 
.A(n_3980),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4180),
.B(n_4183),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_3997),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_SL g4350 ( 
.A(n_3895),
.B(n_2805),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_3998),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_SL g4352 ( 
.A1(n_3939),
.A2(n_1010),
.B1(n_1085),
.B2(n_1008),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4153),
.Y(n_4353)
);

OR2x2_ASAP7_75t_L g4354 ( 
.A(n_3923),
.B(n_3464),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_3969),
.B(n_3469),
.Y(n_4355)
);

AOI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4140),
.A2(n_2626),
.B1(n_2675),
.B2(n_2622),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4161),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4002),
.Y(n_4358)
);

A2O1A1Ixp33_ASAP7_75t_L g4359 ( 
.A1(n_4101),
.A2(n_3857),
.B(n_3987),
.C(n_4154),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_3914),
.B(n_3915),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_3956),
.B(n_2626),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_4142),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4004),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_3872),
.A2(n_4201),
.B(n_4113),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4013),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3856),
.B(n_3938),
.Y(n_4366)
);

BUFx6f_ASAP7_75t_L g4367 ( 
.A(n_4137),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4016),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4020),
.Y(n_4369)
);

AND2x4_ASAP7_75t_L g4370 ( 
.A(n_4183),
.B(n_3349),
.Y(n_4370)
);

BUFx6f_ASAP7_75t_L g4371 ( 
.A(n_4137),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4075),
.B(n_2626),
.Y(n_4372)
);

NOR2x1_ASAP7_75t_L g4373 ( 
.A(n_4054),
.B(n_3382),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_4187),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4024),
.Y(n_4375)
);

AO22x1_ASAP7_75t_L g4376 ( 
.A1(n_4049),
.A2(n_2360),
.B1(n_2182),
.B2(n_1085),
.Y(n_4376)
);

INVx2_ASAP7_75t_SL g4377 ( 
.A(n_4177),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4028),
.Y(n_4378)
);

AND2x4_ASAP7_75t_L g4379 ( 
.A(n_4139),
.B(n_3382),
.Y(n_4379)
);

AOI22xp33_ASAP7_75t_L g4380 ( 
.A1(n_4065),
.A2(n_2707),
.B1(n_2675),
.B2(n_3342),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4029),
.Y(n_4381)
);

NAND2x1p5_ASAP7_75t_L g4382 ( 
.A(n_3879),
.B(n_3382),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_3953),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_3984),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4038),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_3877),
.B(n_2675),
.Y(n_4386)
);

HB1xp67_ASAP7_75t_L g4387 ( 
.A(n_3984),
.Y(n_4387)
);

BUFx6f_ASAP7_75t_L g4388 ( 
.A(n_4177),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_3856),
.B(n_3940),
.Y(n_4389)
);

CKINVDCx20_ASAP7_75t_R g4390 ( 
.A(n_4170),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4064),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4035),
.B(n_3565),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_SL g4393 ( 
.A(n_4032),
.B(n_2805),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_L g4394 ( 
.A(n_3929),
.B(n_2790),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4193),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4074),
.Y(n_4396)
);

NAND2xp33_ASAP7_75t_L g4397 ( 
.A(n_4101),
.B(n_3434),
.Y(n_4397)
);

INVxp67_ASAP7_75t_L g4398 ( 
.A(n_3980),
.Y(n_4398)
);

AND2x4_ASAP7_75t_L g4399 ( 
.A(n_4144),
.B(n_3427),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4080),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_SL g4401 ( 
.A(n_3971),
.B(n_2805),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_3935),
.B(n_4012),
.Y(n_4402)
);

AND2x4_ASAP7_75t_L g4403 ( 
.A(n_3920),
.B(n_3427),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4100),
.Y(n_4404)
);

AND2x4_ASAP7_75t_L g4405 ( 
.A(n_3920),
.B(n_3427),
.Y(n_4405)
);

INVxp67_ASAP7_75t_L g4406 ( 
.A(n_3978),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4103),
.Y(n_4407)
);

INVx2_ASAP7_75t_SL g4408 ( 
.A(n_4177),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4112),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4130),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4152),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4140),
.A2(n_2707),
.B1(n_2893),
.B2(n_2792),
.Y(n_4412)
);

AND2x4_ASAP7_75t_L g4413 ( 
.A(n_3921),
.B(n_3442),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_4199),
.Y(n_4414)
);

OR2x2_ASAP7_75t_L g4415 ( 
.A(n_3957),
.B(n_3474),
.Y(n_4415)
);

INVx2_ASAP7_75t_SL g4416 ( 
.A(n_4200),
.Y(n_4416)
);

NOR2xp33_ASAP7_75t_L g4417 ( 
.A(n_3995),
.B(n_2895),
.Y(n_4417)
);

BUFx3_ASAP7_75t_L g4418 ( 
.A(n_4200),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4157),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4163),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_SL g4421 ( 
.A(n_3971),
.B(n_2805),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4050),
.B(n_3567),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4191),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_4200),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4195),
.Y(n_4425)
);

BUFx3_ASAP7_75t_L g4426 ( 
.A(n_4167),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4052),
.B(n_3568),
.Y(n_4427)
);

INVx4_ASAP7_75t_L g4428 ( 
.A(n_3921),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4053),
.B(n_3569),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_L g4430 ( 
.A(n_3958),
.B(n_2895),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_SL g4431 ( 
.A(n_4040),
.B(n_2805),
.Y(n_4431)
);

INVx4_ASAP7_75t_L g4432 ( 
.A(n_4011),
.Y(n_4432)
);

INVx3_ASAP7_75t_L g4433 ( 
.A(n_4135),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_4040),
.B(n_2854),
.Y(n_4434)
);

HB1xp67_ASAP7_75t_L g4435 ( 
.A(n_4093),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4219),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4203),
.Y(n_4437)
);

BUFx6f_ASAP7_75t_L g4438 ( 
.A(n_4011),
.Y(n_4438)
);

BUFx3_ASAP7_75t_L g4439 ( 
.A(n_4206),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_3908),
.B(n_3570),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_3962),
.B(n_2913),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_4169),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3894),
.B(n_3571),
.Y(n_4443)
);

NOR2xp33_ASAP7_75t_L g4444 ( 
.A(n_3910),
.B(n_2913),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4207),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4212),
.Y(n_4446)
);

AOI22xp5_ASAP7_75t_L g4447 ( 
.A1(n_4104),
.A2(n_2707),
.B1(n_2917),
.B2(n_2915),
.Y(n_4447)
);

CKINVDCx5p33_ASAP7_75t_R g4448 ( 
.A(n_3917),
.Y(n_4448)
);

AND2x4_ASAP7_75t_L g4449 ( 
.A(n_4047),
.B(n_3442),
.Y(n_4449)
);

INVx2_ASAP7_75t_SL g4450 ( 
.A(n_4092),
.Y(n_4450)
);

INVx1_ASAP7_75t_SL g4451 ( 
.A(n_3967),
.Y(n_4451)
);

OR2x6_ASAP7_75t_L g4452 ( 
.A(n_4135),
.B(n_3654),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_SL g4453 ( 
.A(n_3994),
.B(n_4069),
.Y(n_4453)
);

INVx2_ASAP7_75t_SL g4454 ( 
.A(n_4047),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4217),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4229),
.Y(n_4456)
);

AOI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_4108),
.A2(n_2917),
.B1(n_2918),
.B2(n_2915),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_3854),
.Y(n_4458)
);

OR2x2_ASAP7_75t_L g4459 ( 
.A(n_4225),
.B(n_3477),
.Y(n_4459)
);

AOI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4065),
.A2(n_3414),
.B1(n_3428),
.B2(n_3392),
.Y(n_4460)
);

BUFx6f_ASAP7_75t_L g4461 ( 
.A(n_4135),
.Y(n_4461)
);

INVx3_ASAP7_75t_L g4462 ( 
.A(n_4037),
.Y(n_4462)
);

INVxp67_ASAP7_75t_L g4463 ( 
.A(n_3978),
.Y(n_4463)
);

NOR3xp33_ASAP7_75t_SL g4464 ( 
.A(n_4114),
.B(n_979),
.C(n_977),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_SL g4465 ( 
.A(n_4007),
.B(n_2918),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_3872),
.A2(n_3076),
.B(n_3065),
.Y(n_4466)
);

BUFx6f_ASAP7_75t_L g4467 ( 
.A(n_4037),
.Y(n_4467)
);

AOI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4155),
.A2(n_2929),
.B1(n_2933),
.B2(n_2921),
.Y(n_4468)
);

NOR2xp33_ASAP7_75t_L g4469 ( 
.A(n_4051),
.B(n_2921),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_SL g4470 ( 
.A(n_4061),
.B(n_2929),
.Y(n_4470)
);

OR2x2_ASAP7_75t_L g4471 ( 
.A(n_4061),
.B(n_3481),
.Y(n_4471)
);

INVx6_ASAP7_75t_L g4472 ( 
.A(n_4182),
.Y(n_4472)
);

NOR2xp33_ASAP7_75t_L g4473 ( 
.A(n_4115),
.B(n_2933),
.Y(n_4473)
);

NAND2x1p5_ASAP7_75t_L g4474 ( 
.A(n_3879),
.B(n_3020),
.Y(n_4474)
);

INVx3_ASAP7_75t_L g4475 ( 
.A(n_4182),
.Y(n_4475)
);

OR2x2_ASAP7_75t_L g4476 ( 
.A(n_4093),
.B(n_3576),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_3899),
.B(n_3578),
.Y(n_4477)
);

BUFx12f_ASAP7_75t_L g4478 ( 
.A(n_4124),
.Y(n_4478)
);

AOI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4155),
.A2(n_4141),
.B1(n_4143),
.B2(n_4208),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4079),
.B(n_3581),
.Y(n_4480)
);

INVx2_ASAP7_75t_SL g4481 ( 
.A(n_4158),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_3864),
.Y(n_4482)
);

NOR2xp33_ASAP7_75t_R g4483 ( 
.A(n_4125),
.B(n_4128),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3875),
.B(n_3582),
.Y(n_4484)
);

AOI211xp5_ASAP7_75t_L g4485 ( 
.A1(n_4126),
.A2(n_1091),
.B(n_1108),
.C(n_1010),
.Y(n_4485)
);

BUFx3_ASAP7_75t_L g4486 ( 
.A(n_4209),
.Y(n_4486)
);

NOR2x1p5_ASAP7_75t_L g4487 ( 
.A(n_4014),
.B(n_2389),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_3890),
.Y(n_4488)
);

CKINVDCx20_ASAP7_75t_R g4489 ( 
.A(n_4120),
.Y(n_4489)
);

OAI22xp5_ASAP7_75t_SL g4490 ( 
.A1(n_3939),
.A2(n_1091),
.B1(n_1120),
.B2(n_1108),
.Y(n_4490)
);

AND2x4_ASAP7_75t_L g4491 ( 
.A(n_4182),
.B(n_4147),
.Y(n_4491)
);

NOR2xp33_ASAP7_75t_R g4492 ( 
.A(n_4129),
.B(n_2182),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4072),
.B(n_3583),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_3896),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_3949),
.B(n_3584),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_3909),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_3912),
.B(n_3585),
.Y(n_4497)
);

OAI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4055),
.A2(n_2936),
.B1(n_2939),
.B2(n_2935),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_3884),
.B(n_3586),
.Y(n_4499)
);

AND2x2_ASAP7_75t_SL g4500 ( 
.A(n_4126),
.B(n_2389),
.Y(n_4500)
);

CKINVDCx5p33_ASAP7_75t_R g4501 ( 
.A(n_3972),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_3881),
.B(n_4067),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_4067),
.B(n_3589),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4068),
.B(n_3590),
.Y(n_4504)
);

AOI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_4141),
.A2(n_2936),
.B1(n_2939),
.B2(n_2935),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_3922),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4068),
.B(n_3592),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4081),
.B(n_3594),
.Y(n_4508)
);

INVx4_ASAP7_75t_L g4509 ( 
.A(n_3880),
.Y(n_4509)
);

OR2x6_ASAP7_75t_L g4510 ( 
.A(n_4087),
.B(n_3712),
.Y(n_4510)
);

INVx4_ASAP7_75t_L g4511 ( 
.A(n_3880),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_3931),
.Y(n_4512)
);

AND2x4_ASAP7_75t_L g4513 ( 
.A(n_3904),
.B(n_3392),
.Y(n_4513)
);

AND2x6_ASAP7_75t_L g4514 ( 
.A(n_3904),
.B(n_3596),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_3937),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_L g4516 ( 
.A(n_3950),
.B(n_2940),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_3913),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_3944),
.Y(n_4518)
);

BUFx6f_ASAP7_75t_L g4519 ( 
.A(n_4189),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4084),
.B(n_3598),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4089),
.B(n_3600),
.Y(n_4521)
);

NOR2x2_ASAP7_75t_L g4522 ( 
.A(n_4151),
.B(n_3407),
.Y(n_4522)
);

AND2x2_ASAP7_75t_L g4523 ( 
.A(n_3970),
.B(n_3414),
.Y(n_4523)
);

AND2x4_ASAP7_75t_L g4524 ( 
.A(n_3913),
.B(n_3428),
.Y(n_4524)
);

AND2x4_ASAP7_75t_L g4525 ( 
.A(n_4110),
.B(n_3601),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3945),
.Y(n_4526)
);

INVx3_ASAP7_75t_L g4527 ( 
.A(n_3954),
.Y(n_4527)
);

OAI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_4097),
.A2(n_3612),
.B1(n_3614),
.B2(n_3607),
.Y(n_4528)
);

HB1xp67_ASAP7_75t_L g4529 ( 
.A(n_3970),
.Y(n_4529)
);

INVxp67_ASAP7_75t_SL g4530 ( 
.A(n_3928),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_3946),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_3951),
.Y(n_4532)
);

NOR3xp33_ASAP7_75t_SL g4533 ( 
.A(n_4097),
.B(n_983),
.C(n_981),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4090),
.B(n_3824),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_L g4535 ( 
.A(n_4091),
.B(n_3828),
.Y(n_4535)
);

BUFx8_ASAP7_75t_L g4536 ( 
.A(n_3959),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4094),
.B(n_3831),
.Y(n_4537)
);

NOR2xp67_ASAP7_75t_L g4538 ( 
.A(n_3906),
.B(n_3400),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4105),
.B(n_3833),
.Y(n_4539)
);

BUFx12f_ASAP7_75t_SL g4540 ( 
.A(n_4162),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4107),
.B(n_3834),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_3961),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_3960),
.B(n_2940),
.Y(n_4543)
);

INVx2_ASAP7_75t_SL g4544 ( 
.A(n_4078),
.Y(n_4544)
);

OR2x6_ASAP7_75t_SL g4545 ( 
.A(n_3964),
.B(n_984),
.Y(n_4545)
);

BUFx3_ASAP7_75t_L g4546 ( 
.A(n_4096),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_3982),
.Y(n_4547)
);

INVx2_ASAP7_75t_SL g4548 ( 
.A(n_4082),
.Y(n_4548)
);

AOI22xp33_ASAP7_75t_L g4549 ( 
.A1(n_3861),
.A2(n_4154),
.B1(n_3905),
.B2(n_4143),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_3993),
.Y(n_4550)
);

CKINVDCx5p33_ASAP7_75t_R g4551 ( 
.A(n_4186),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4086),
.B(n_3835),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_4086),
.B(n_3843),
.Y(n_4553)
);

INVxp67_ASAP7_75t_SL g4554 ( 
.A(n_4116),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_3996),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4008),
.Y(n_4556)
);

AOI22xp5_ASAP7_75t_L g4557 ( 
.A1(n_4196),
.A2(n_2943),
.B1(n_2945),
.B2(n_2942),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4010),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_3861),
.A2(n_2943),
.B1(n_2945),
.B2(n_2942),
.Y(n_4559)
);

NAND2x1p5_ASAP7_75t_L g4560 ( 
.A(n_3954),
.B(n_3020),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4009),
.B(n_3845),
.Y(n_4561)
);

AOI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_4226),
.A2(n_2949),
.B1(n_2952),
.B2(n_2947),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4015),
.Y(n_4563)
);

OAI22xp5_ASAP7_75t_L g4564 ( 
.A1(n_4009),
.A2(n_2949),
.B1(n_2952),
.B2(n_2947),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4034),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4174),
.Y(n_4566)
);

BUFx3_ASAP7_75t_L g4567 ( 
.A(n_4205),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_3990),
.B(n_3848),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_SL g4569 ( 
.A(n_3966),
.B(n_2953),
.Y(n_4569)
);

INVx2_ASAP7_75t_SL g4570 ( 
.A(n_4083),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4098),
.A2(n_2954),
.B1(n_2957),
.B2(n_2953),
.Y(n_4571)
);

INVx3_ASAP7_75t_L g4572 ( 
.A(n_4121),
.Y(n_4572)
);

HB1xp67_ASAP7_75t_L g4573 ( 
.A(n_4118),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4119),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_3990),
.B(n_3851),
.Y(n_4575)
);

INVx2_ASAP7_75t_SL g4576 ( 
.A(n_4121),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_3975),
.B(n_3853),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4123),
.Y(n_4578)
);

AOI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_3986),
.A2(n_2957),
.B1(n_2959),
.B2(n_2954),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4174),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4227),
.B(n_4005),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4227),
.Y(n_4582)
);

OR2x2_ASAP7_75t_SL g4583 ( 
.A(n_4131),
.B(n_820),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_4134),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_SL g4585 ( 
.A(n_4005),
.B(n_2959),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4025),
.B(n_3748),
.Y(n_4586)
);

INVxp67_ASAP7_75t_SL g4587 ( 
.A(n_3941),
.Y(n_4587)
);

CKINVDCx5p33_ASAP7_75t_R g4588 ( 
.A(n_4127),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4149),
.Y(n_4589)
);

AOI22xp33_ASAP7_75t_L g4590 ( 
.A1(n_3936),
.A2(n_2965),
.B1(n_2968),
.B2(n_2960),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4145),
.Y(n_4591)
);

OAI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_3869),
.A2(n_3448),
.B(n_3238),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_SL g4593 ( 
.A(n_3855),
.B(n_2960),
.Y(n_4593)
);

HB1xp67_ASAP7_75t_L g4594 ( 
.A(n_4146),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4027),
.B(n_3751),
.Y(n_4595)
);

AOI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_3878),
.A2(n_3076),
.B(n_3065),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_3952),
.B(n_2965),
.Y(n_4597)
);

NOR2xp33_ASAP7_75t_L g4598 ( 
.A(n_3866),
.B(n_2973),
.Y(n_4598)
);

INVx3_ASAP7_75t_L g4599 ( 
.A(n_4214),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4156),
.Y(n_4600)
);

AND2x6_ASAP7_75t_SL g4601 ( 
.A(n_3887),
.B(n_820),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4164),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4166),
.Y(n_4603)
);

NOR3xp33_ASAP7_75t_SL g4604 ( 
.A(n_3942),
.B(n_988),
.C(n_985),
.Y(n_4604)
);

BUFx3_ASAP7_75t_L g4605 ( 
.A(n_4214),
.Y(n_4605)
);

BUFx2_ASAP7_75t_L g4606 ( 
.A(n_3889),
.Y(n_4606)
);

CKINVDCx20_ASAP7_75t_R g4607 ( 
.A(n_4213),
.Y(n_4607)
);

INVx2_ASAP7_75t_SL g4608 ( 
.A(n_4168),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4018),
.B(n_3756),
.Y(n_4609)
);

NOR2xp33_ASAP7_75t_R g4610 ( 
.A(n_3882),
.B(n_2182),
.Y(n_4610)
);

INVx3_ASAP7_75t_L g4611 ( 
.A(n_3925),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4022),
.B(n_3758),
.Y(n_4612)
);

INVx5_ASAP7_75t_L g4613 ( 
.A(n_3925),
.Y(n_4613)
);

BUFx3_ASAP7_75t_L g4614 ( 
.A(n_3883),
.Y(n_4614)
);

A2O1A1Ixp33_ASAP7_75t_SL g4615 ( 
.A1(n_3987),
.A2(n_3405),
.B(n_3406),
.C(n_3400),
.Y(n_4615)
);

INVx3_ASAP7_75t_L g4616 ( 
.A(n_3925),
.Y(n_4616)
);

AOI21xp5_ASAP7_75t_L g4617 ( 
.A1(n_3974),
.A2(n_3085),
.B(n_3082),
.Y(n_4617)
);

AND3x1_ASAP7_75t_L g4618 ( 
.A(n_4176),
.B(n_825),
.C(n_750),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_SL g4619 ( 
.A(n_3943),
.B(n_3226),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4171),
.Y(n_4620)
);

BUFx8_ASAP7_75t_L g4621 ( 
.A(n_3925),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4173),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4175),
.Y(n_4623)
);

OR2x2_ASAP7_75t_L g4624 ( 
.A(n_3948),
.B(n_3759),
.Y(n_4624)
);

CKINVDCx5p33_ASAP7_75t_R g4625 ( 
.A(n_4023),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_SL g4626 ( 
.A(n_3963),
.B(n_3264),
.Y(n_4626)
);

INVx2_ASAP7_75t_L g4627 ( 
.A(n_4181),
.Y(n_4627)
);

AND2x6_ASAP7_75t_SL g4628 ( 
.A(n_4184),
.B(n_826),
.Y(n_4628)
);

AND2x6_ASAP7_75t_L g4629 ( 
.A(n_4185),
.B(n_3762),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4197),
.Y(n_4630)
);

AOI22xp33_ASAP7_75t_L g4631 ( 
.A1(n_3991),
.A2(n_2563),
.B1(n_2564),
.B2(n_2562),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4202),
.B(n_3763),
.Y(n_4632)
);

AO32x1_ASAP7_75t_L g4633 ( 
.A1(n_4235),
.A2(n_3900),
.A3(n_3932),
.B1(n_4026),
.B2(n_3870),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4308),
.B(n_4000),
.Y(n_4634)
);

OAI321xp33_ASAP7_75t_L g4635 ( 
.A1(n_4352),
.A2(n_1194),
.A3(n_1024),
.B1(n_4001),
.B2(n_1037),
.C(n_1075),
.Y(n_4635)
);

AOI22xp33_ASAP7_75t_L g4636 ( 
.A1(n_4286),
.A2(n_3859),
.B1(n_3860),
.B2(n_4176),
.Y(n_4636)
);

AOI21xp5_ASAP7_75t_L g4637 ( 
.A1(n_4434),
.A2(n_3930),
.B(n_3974),
.Y(n_4637)
);

O2A1O1Ixp33_ASAP7_75t_L g4638 ( 
.A1(n_4359),
.A2(n_3947),
.B(n_3891),
.C(n_4048),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4240),
.B(n_4215),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4240),
.B(n_4218),
.Y(n_4640)
);

AOI21xp5_ASAP7_75t_L g4641 ( 
.A1(n_4397),
.A2(n_4364),
.B(n_4323),
.Y(n_4641)
);

INVx3_ASAP7_75t_L g4642 ( 
.A(n_4461),
.Y(n_4642)
);

AOI33xp33_ASAP7_75t_L g4643 ( 
.A1(n_4485),
.A2(n_1188),
.A3(n_1121),
.B1(n_1148),
.B2(n_1120),
.B3(n_826),
.Y(n_4643)
);

AND2x4_ASAP7_75t_L g4644 ( 
.A(n_4291),
.B(n_4190),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4299),
.B(n_4224),
.Y(n_4645)
);

AOI21xp5_ASAP7_75t_L g4646 ( 
.A1(n_4364),
.A2(n_3930),
.B(n_3985),
.Y(n_4646)
);

OAI22xp5_ASAP7_75t_L g4647 ( 
.A1(n_4479),
.A2(n_4228),
.B1(n_4230),
.B2(n_4159),
.Y(n_4647)
);

O2A1O1Ixp33_ASAP7_75t_L g4648 ( 
.A1(n_4345),
.A2(n_4465),
.B(n_4533),
.C(n_4453),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4299),
.B(n_4178),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4366),
.B(n_4178),
.Y(n_4650)
);

OAI22xp33_ASAP7_75t_L g4651 ( 
.A1(n_4588),
.A2(n_3286),
.B1(n_3323),
.B2(n_3268),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4361),
.B(n_4033),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4451),
.B(n_4036),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4246),
.Y(n_4654)
);

NOR2xp67_ASAP7_75t_L g4655 ( 
.A(n_4406),
.B(n_4039),
.Y(n_4655)
);

NAND3xp33_ASAP7_75t_SL g4656 ( 
.A(n_4562),
.B(n_1148),
.C(n_1121),
.Y(n_4656)
);

AND2x2_ASAP7_75t_L g4657 ( 
.A(n_4451),
.B(n_4198),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_SL g4658 ( 
.A(n_4362),
.B(n_2360),
.Y(n_4658)
);

O2A1O1Ixp33_ASAP7_75t_L g4659 ( 
.A1(n_4307),
.A2(n_1188),
.B(n_825),
.C(n_1037),
.Y(n_4659)
);

BUFx6f_ASAP7_75t_SL g4660 ( 
.A(n_4233),
.Y(n_4660)
);

OAI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4406),
.A2(n_4463),
.B1(n_4473),
.B2(n_4490),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4366),
.B(n_4179),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4389),
.B(n_4179),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4552),
.A2(n_3985),
.B(n_4132),
.Y(n_4664)
);

NOR2xp33_ASAP7_75t_L g4665 ( 
.A(n_4567),
.B(n_2360),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4389),
.B(n_4188),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4360),
.B(n_4188),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4360),
.B(n_3764),
.Y(n_4668)
);

NOR2x1_ASAP7_75t_L g4669 ( 
.A(n_4341),
.B(n_4041),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_SL g4670 ( 
.A(n_4444),
.B(n_3989),
.Y(n_4670)
);

NAND3xp33_ASAP7_75t_L g4671 ( 
.A(n_4549),
.B(n_2360),
.C(n_995),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4554),
.B(n_3765),
.Y(n_4672)
);

INVx3_ASAP7_75t_L g4673 ( 
.A(n_4461),
.Y(n_4673)
);

NOR2xp33_ASAP7_75t_L g4674 ( 
.A(n_4402),
.B(n_992),
.Y(n_4674)
);

A2O1A1Ixp33_ASAP7_75t_L g4675 ( 
.A1(n_4500),
.A2(n_3989),
.B(n_4160),
.C(n_4216),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4574),
.B(n_3766),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4578),
.B(n_3773),
.Y(n_4677)
);

OAI22xp5_ASAP7_75t_L g4678 ( 
.A1(n_4463),
.A2(n_4546),
.B1(n_4244),
.B2(n_4398),
.Y(n_4678)
);

NOR3xp33_ASAP7_75t_L g4679 ( 
.A(n_4376),
.B(n_4223),
.C(n_976),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4552),
.A2(n_3068),
.B(n_3044),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4584),
.B(n_3778),
.Y(n_4681)
);

INVx2_ASAP7_75t_SL g4682 ( 
.A(n_4234),
.Y(n_4682)
);

CKINVDCx20_ASAP7_75t_R g4683 ( 
.A(n_4236),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4347),
.A2(n_3320),
.B1(n_3715),
.B2(n_3712),
.Y(n_4684)
);

NOR2xp67_ASAP7_75t_L g4685 ( 
.A(n_4263),
.B(n_4220),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4591),
.B(n_3779),
.Y(n_4686)
);

O2A1O1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4258),
.A2(n_825),
.B(n_1037),
.C(n_976),
.Y(n_4687)
);

NAND3xp33_ASAP7_75t_L g4688 ( 
.A(n_4604),
.B(n_1000),
.C(n_997),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_SL g4689 ( 
.A(n_4394),
.B(n_4430),
.Y(n_4689)
);

BUFx2_ASAP7_75t_L g4690 ( 
.A(n_4272),
.Y(n_4690)
);

AOI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4553),
.A2(n_3068),
.B(n_3044),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4239),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4553),
.A2(n_3068),
.B(n_3044),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4573),
.B(n_3780),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4594),
.B(n_3783),
.Y(n_4695)
);

NAND2x1p5_ASAP7_75t_L g4696 ( 
.A(n_4613),
.B(n_4326),
.Y(n_4696)
);

AOI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4401),
.A2(n_3068),
.B(n_3044),
.Y(n_4697)
);

OAI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4441),
.A2(n_2867),
.B(n_2889),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4606),
.B(n_3785),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4250),
.Y(n_4700)
);

AOI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4421),
.A2(n_3364),
.B(n_3068),
.Y(n_4701)
);

AO21x1_ASAP7_75t_L g4702 ( 
.A1(n_4235),
.A2(n_4222),
.B(n_835),
.Y(n_4702)
);

CKINVDCx8_ASAP7_75t_R g4703 ( 
.A(n_4249),
.Y(n_4703)
);

OAI21xp5_ASAP7_75t_L g4704 ( 
.A1(n_4238),
.A2(n_3362),
.B(n_3325),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4254),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4530),
.B(n_3786),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_SL g4707 ( 
.A(n_4610),
.B(n_3386),
.Y(n_4707)
);

AOI21xp5_ASAP7_75t_L g4708 ( 
.A1(n_4431),
.A2(n_3364),
.B(n_3085),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_SL g4709 ( 
.A(n_4457),
.B(n_3402),
.Y(n_4709)
);

NAND2x1p5_ASAP7_75t_L g4710 ( 
.A(n_4613),
.B(n_3082),
.Y(n_4710)
);

CKINVDCx10_ASAP7_75t_R g4711 ( 
.A(n_4231),
.Y(n_4711)
);

A2O1A1Ixp33_ASAP7_75t_L g4712 ( 
.A1(n_4468),
.A2(n_1075),
.B(n_1234),
.C(n_1079),
.Y(n_4712)
);

AND2x4_ASAP7_75t_L g4713 ( 
.A(n_4291),
.B(n_3789),
.Y(n_4713)
);

OAI21xp5_ASAP7_75t_L g4714 ( 
.A1(n_4593),
.A2(n_3424),
.B(n_3419),
.Y(n_4714)
);

AOI21xp5_ASAP7_75t_L g4715 ( 
.A1(n_4278),
.A2(n_4237),
.B(n_4262),
.Y(n_4715)
);

OAI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_4447),
.A2(n_3320),
.B1(n_3715),
.B2(n_3448),
.Y(n_4716)
);

AOI21x1_ASAP7_75t_L g4717 ( 
.A1(n_4617),
.A2(n_3631),
.B(n_4596),
.Y(n_4717)
);

BUFx2_ASAP7_75t_SL g4718 ( 
.A(n_4283),
.Y(n_4718)
);

INVx3_ASAP7_75t_L g4719 ( 
.A(n_4461),
.Y(n_4719)
);

INVxp67_ASAP7_75t_L g4720 ( 
.A(n_4319),
.Y(n_4720)
);

OR2x2_ASAP7_75t_L g4721 ( 
.A(n_4529),
.B(n_3791),
.Y(n_4721)
);

INVx3_ASAP7_75t_L g4722 ( 
.A(n_4467),
.Y(n_4722)
);

OAI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4607),
.A2(n_3437),
.B1(n_3431),
.B2(n_3792),
.Y(n_4723)
);

A2O1A1Ixp33_ASAP7_75t_L g4724 ( 
.A1(n_4581),
.A2(n_1075),
.B(n_1234),
.C(n_1079),
.Y(n_4724)
);

O2A1O1Ixp33_ASAP7_75t_L g4725 ( 
.A1(n_4393),
.A2(n_4498),
.B(n_4585),
.C(n_4615),
.Y(n_4725)
);

AOI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4278),
.A2(n_4237),
.B(n_4242),
.Y(n_4726)
);

OR2x6_ASAP7_75t_L g4727 ( 
.A(n_4510),
.B(n_3364),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4587),
.B(n_3793),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4589),
.B(n_3794),
.Y(n_4729)
);

O2A1O1Ixp33_ASAP7_75t_SL g4730 ( 
.A1(n_4329),
.A2(n_1079),
.B(n_1234),
.C(n_976),
.Y(n_4730)
);

AND2x4_ASAP7_75t_L g4731 ( 
.A(n_4475),
.B(n_3795),
.Y(n_4731)
);

AND2x4_ASAP7_75t_L g4732 ( 
.A(n_4475),
.B(n_4491),
.Y(n_4732)
);

NOR3xp33_ASAP7_75t_L g4733 ( 
.A(n_4481),
.B(n_835),
.C(n_829),
.Y(n_4733)
);

NAND2x1p5_ASAP7_75t_L g4734 ( 
.A(n_4613),
.B(n_3082),
.Y(n_4734)
);

NOR2xp33_ASAP7_75t_L g4735 ( 
.A(n_4448),
.B(n_1002),
.Y(n_4735)
);

INVx5_ASAP7_75t_L g4736 ( 
.A(n_4514),
.Y(n_4736)
);

OAI21xp5_ASAP7_75t_L g4737 ( 
.A1(n_4505),
.A2(n_2843),
.B(n_2894),
.Y(n_4737)
);

NAND3xp33_ASAP7_75t_L g4738 ( 
.A(n_4618),
.B(n_1005),
.C(n_1003),
.Y(n_4738)
);

OAI21xp5_ASAP7_75t_L g4739 ( 
.A1(n_4516),
.A2(n_2956),
.B(n_2896),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4600),
.B(n_3796),
.Y(n_4740)
);

NOR2xp33_ASAP7_75t_L g4741 ( 
.A(n_4551),
.B(n_1014),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4602),
.B(n_2181),
.Y(n_4742)
);

AOI21xp5_ASAP7_75t_L g4743 ( 
.A1(n_4242),
.A2(n_4243),
.B(n_4270),
.Y(n_4743)
);

A2O1A1Ixp33_ASAP7_75t_L g4744 ( 
.A1(n_4581),
.A2(n_3364),
.B(n_837),
.C(n_842),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4603),
.B(n_2181),
.Y(n_4745)
);

NAND2x1p5_ASAP7_75t_L g4746 ( 
.A(n_4613),
.B(n_3085),
.Y(n_4746)
);

AND2x2_ASAP7_75t_L g4747 ( 
.A(n_4523),
.B(n_1641),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4622),
.B(n_2181),
.Y(n_4748)
);

AOI22xp5_ASAP7_75t_L g4749 ( 
.A1(n_4489),
.A2(n_4277),
.B1(n_4390),
.B2(n_4450),
.Y(n_4749)
);

INVx4_ASAP7_75t_L g4750 ( 
.A(n_4438),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4623),
.B(n_4630),
.Y(n_4751)
);

NOR2xp33_ASAP7_75t_L g4752 ( 
.A(n_4545),
.B(n_1015),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_L g4753 ( 
.A(n_4620),
.B(n_2181),
.Y(n_4753)
);

HB1xp67_ASAP7_75t_L g4754 ( 
.A(n_4259),
.Y(n_4754)
);

NOR2xp33_ASAP7_75t_SL g4755 ( 
.A(n_4540),
.B(n_3072),
.Y(n_4755)
);

INVxp67_ASAP7_75t_L g4756 ( 
.A(n_4257),
.Y(n_4756)
);

OAI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4469),
.A2(n_2975),
.B(n_3350),
.Y(n_4757)
);

BUFx3_ASAP7_75t_L g4758 ( 
.A(n_4267),
.Y(n_4758)
);

AOI21xp5_ASAP7_75t_L g4759 ( 
.A1(n_4243),
.A2(n_3364),
.B(n_3202),
.Y(n_4759)
);

OAI22xp5_ASAP7_75t_L g4760 ( 
.A1(n_4412),
.A2(n_3094),
.B1(n_3063),
.B2(n_3353),
.Y(n_4760)
);

AOI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_4270),
.A2(n_3202),
.B(n_3142),
.Y(n_4761)
);

INVx3_ASAP7_75t_L g4762 ( 
.A(n_4467),
.Y(n_4762)
);

NOR2x1p5_ASAP7_75t_SL g4763 ( 
.A(n_4624),
.B(n_3925),
.Y(n_4763)
);

NAND3xp33_ASAP7_75t_L g4764 ( 
.A(n_4464),
.B(n_1019),
.C(n_1018),
.Y(n_4764)
);

BUFx6f_ASAP7_75t_L g4765 ( 
.A(n_4251),
.Y(n_4765)
);

OAI21xp5_ASAP7_75t_L g4766 ( 
.A1(n_4598),
.A2(n_3409),
.B(n_3367),
.Y(n_4766)
);

O2A1O1Ixp33_ASAP7_75t_L g4767 ( 
.A1(n_4470),
.A2(n_837),
.B(n_842),
.C(n_829),
.Y(n_4767)
);

A2O1A1Ixp33_ASAP7_75t_L g4768 ( 
.A1(n_4346),
.A2(n_847),
.B(n_849),
.C(n_844),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4264),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4592),
.A2(n_3202),
.B(n_3142),
.Y(n_4770)
);

NOR2xp33_ASAP7_75t_L g4771 ( 
.A(n_4439),
.B(n_1020),
.Y(n_4771)
);

AOI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4592),
.A2(n_3212),
.B(n_3142),
.Y(n_4772)
);

AND2x2_ASAP7_75t_L g4773 ( 
.A(n_4372),
.B(n_1641),
.Y(n_4773)
);

OAI21xp5_ASAP7_75t_L g4774 ( 
.A1(n_4296),
.A2(n_4557),
.B(n_4559),
.Y(n_4774)
);

AOI22xp33_ASAP7_75t_L g4775 ( 
.A1(n_4625),
.A2(n_1042),
.B1(n_2755),
.B2(n_2603),
.Y(n_4775)
);

CKINVDCx5p33_ASAP7_75t_R g4776 ( 
.A(n_4297),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4386),
.B(n_1646),
.Y(n_4777)
);

BUFx3_ASAP7_75t_L g4778 ( 
.A(n_4536),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_L g4779 ( 
.A(n_4614),
.B(n_3413),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4304),
.A2(n_3243),
.B(n_3212),
.Y(n_4780)
);

AOI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4304),
.A2(n_3243),
.B(n_3212),
.Y(n_4781)
);

INVx1_ASAP7_75t_SL g4782 ( 
.A(n_4265),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4486),
.B(n_4601),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4282),
.B(n_1646),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4255),
.Y(n_4785)
);

BUFx2_ASAP7_75t_L g4786 ( 
.A(n_4536),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4312),
.A2(n_3250),
.B(n_3243),
.Y(n_4787)
);

NAND2x1p5_ASAP7_75t_L g4788 ( 
.A(n_4326),
.B(n_3250),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4499),
.B(n_4329),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4499),
.B(n_3413),
.Y(n_4790)
);

BUFx2_ASAP7_75t_L g4791 ( 
.A(n_4384),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_SL g4792 ( 
.A(n_4337),
.B(n_3925),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4312),
.A2(n_3254),
.B(n_3250),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4337),
.B(n_3416),
.Y(n_4794)
);

NOR2xp33_ASAP7_75t_L g4795 ( 
.A(n_4245),
.B(n_1025),
.Y(n_4795)
);

NAND3xp33_ASAP7_75t_SL g4796 ( 
.A(n_4315),
.B(n_1038),
.C(n_1031),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4273),
.Y(n_4797)
);

OAI22xp5_ASAP7_75t_L g4798 ( 
.A1(n_4460),
.A2(n_3045),
.B1(n_3327),
.B2(n_3218),
.Y(n_4798)
);

NOR2xp33_ASAP7_75t_L g4799 ( 
.A(n_4245),
.B(n_1039),
.Y(n_4799)
);

CKINVDCx10_ASAP7_75t_R g4800 ( 
.A(n_4247),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_SL g4801 ( 
.A(n_4566),
.B(n_4070),
.Y(n_4801)
);

AO22x1_ASAP7_75t_L g4802 ( 
.A1(n_4501),
.A2(n_847),
.B1(n_849),
.B2(n_844),
.Y(n_4802)
);

NOR2xp33_ASAP7_75t_L g4803 ( 
.A(n_4628),
.B(n_1046),
.Y(n_4803)
);

NAND3xp33_ASAP7_75t_L g4804 ( 
.A(n_4417),
.B(n_1052),
.C(n_1049),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4287),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4627),
.B(n_2327),
.Y(n_4806)
);

INVx1_ASAP7_75t_SL g4807 ( 
.A(n_4331),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4253),
.B(n_4266),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4253),
.B(n_3416),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4269),
.Y(n_4810)
);

NOR2xp67_ASAP7_75t_L g4811 ( 
.A(n_4544),
.B(n_3400),
.Y(n_4811)
);

OR2x6_ASAP7_75t_SL g4812 ( 
.A(n_4442),
.B(n_1054),
.Y(n_4812)
);

NOR2xp33_ASAP7_75t_L g4813 ( 
.A(n_4478),
.B(n_1055),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4583),
.A2(n_3399),
.B1(n_3403),
.B2(n_3396),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4276),
.A2(n_3403),
.B1(n_3404),
.B2(n_3399),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4266),
.B(n_3425),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4274),
.B(n_3425),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4274),
.B(n_3429),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4348),
.B(n_1059),
.Y(n_4819)
);

AOI21xp5_ASAP7_75t_L g4820 ( 
.A1(n_4596),
.A2(n_3340),
.B(n_3254),
.Y(n_4820)
);

AOI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_4333),
.A2(n_3340),
.B(n_3254),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_SL g4822 ( 
.A(n_4580),
.B(n_4070),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4279),
.B(n_3429),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4303),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4279),
.B(n_3433),
.Y(n_4825)
);

A2O1A1Ixp33_ASAP7_75t_L g4826 ( 
.A1(n_4525),
.A2(n_855),
.B(n_858),
.C(n_851),
.Y(n_4826)
);

NOR3xp33_ASAP7_75t_L g4827 ( 
.A(n_4543),
.B(n_855),
.C(n_851),
.Y(n_4827)
);

NOR2xp33_ASAP7_75t_L g4828 ( 
.A(n_4348),
.B(n_1061),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4392),
.A2(n_3361),
.B(n_3340),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_SL g4830 ( 
.A(n_4582),
.B(n_4070),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4284),
.B(n_3433),
.Y(n_4831)
);

BUFx12f_ASAP7_75t_L g4832 ( 
.A(n_4383),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4284),
.B(n_3438),
.Y(n_4833)
);

INVx1_ASAP7_75t_SL g4834 ( 
.A(n_4483),
.Y(n_4834)
);

O2A1O1Ixp33_ASAP7_75t_L g4835 ( 
.A1(n_4548),
.A2(n_859),
.B(n_861),
.C(n_858),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4280),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4290),
.B(n_3438),
.Y(n_4837)
);

OAI21x1_ASAP7_75t_L g4838 ( 
.A1(n_4617),
.A2(n_3271),
.B(n_3204),
.Y(n_4838)
);

BUFx2_ASAP7_75t_L g4839 ( 
.A(n_4292),
.Y(n_4839)
);

OAI21xp5_ASAP7_75t_L g4840 ( 
.A1(n_4252),
.A2(n_4339),
.B(n_4302),
.Y(n_4840)
);

OAI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4619),
.A2(n_2810),
.B(n_2784),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4288),
.Y(n_4842)
);

NOR2xp33_ASAP7_75t_L g4843 ( 
.A(n_4570),
.B(n_1063),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_L g4844 ( 
.A(n_4387),
.B(n_1066),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4318),
.Y(n_4845)
);

CKINVDCx16_ASAP7_75t_R g4846 ( 
.A(n_4492),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_SL g4847 ( 
.A(n_4525),
.B(n_4477),
.Y(n_4847)
);

O2A1O1Ixp33_ASAP7_75t_L g4848 ( 
.A1(n_4344),
.A2(n_861),
.B(n_866),
.C(n_859),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4290),
.B(n_3441),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4443),
.B(n_3441),
.Y(n_4850)
);

OAI22xp5_ASAP7_75t_L g4851 ( 
.A1(n_4380),
.A2(n_3404),
.B1(n_3366),
.B2(n_3361),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4392),
.A2(n_3366),
.B(n_3361),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4422),
.A2(n_3366),
.B(n_3072),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4443),
.B(n_4497),
.Y(n_4854)
);

AOI22x1_ASAP7_75t_L g4855 ( 
.A1(n_4487),
.A2(n_1071),
.B1(n_1072),
.B2(n_1068),
.Y(n_4855)
);

OAI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4356),
.A2(n_3072),
.B1(n_3147),
.B2(n_3020),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4497),
.B(n_3443),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4289),
.Y(n_4858)
);

OAI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4626),
.A2(n_2755),
.B(n_2603),
.Y(n_4859)
);

OAI21xp33_ASAP7_75t_L g4860 ( 
.A1(n_4568),
.A2(n_1080),
.B(n_1078),
.Y(n_4860)
);

AOI21xp5_ASAP7_75t_L g4861 ( 
.A1(n_4422),
.A2(n_3147),
.B(n_3072),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4440),
.B(n_4480),
.Y(n_4862)
);

AOI21xp5_ASAP7_75t_L g4863 ( 
.A1(n_4427),
.A2(n_4429),
.B(n_4324),
.Y(n_4863)
);

BUFx6f_ASAP7_75t_L g4864 ( 
.A(n_4295),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_SL g4865 ( 
.A(n_4477),
.B(n_4373),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4629),
.A2(n_2755),
.B1(n_2970),
.B2(n_2603),
.Y(n_4866)
);

AND2x4_ASAP7_75t_L g4867 ( 
.A(n_4491),
.B(n_3443),
.Y(n_4867)
);

AND2x4_ASAP7_75t_SL g4868 ( 
.A(n_4283),
.B(n_3338),
.Y(n_4868)
);

AOI21xp5_ASAP7_75t_L g4869 ( 
.A1(n_4427),
.A2(n_4429),
.B(n_4466),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4330),
.Y(n_4870)
);

BUFx6f_ASAP7_75t_L g4871 ( 
.A(n_4295),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_SL g4872 ( 
.A(n_4495),
.B(n_4070),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4440),
.B(n_3445),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4415),
.B(n_2339),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4480),
.B(n_2339),
.Y(n_4875)
);

CKINVDCx14_ASAP7_75t_R g4876 ( 
.A(n_4426),
.Y(n_4876)
);

AOI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4466),
.A2(n_3177),
.B(n_3147),
.Y(n_4877)
);

AND2x4_ASAP7_75t_L g4878 ( 
.A(n_4232),
.B(n_3445),
.Y(n_4878)
);

AO21x1_ASAP7_75t_L g4879 ( 
.A1(n_4241),
.A2(n_868),
.B(n_866),
.Y(n_4879)
);

INVx3_ASAP7_75t_L g4880 ( 
.A(n_4467),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4495),
.B(n_2340),
.Y(n_4881)
);

NAND2xp33_ASAP7_75t_L g4882 ( 
.A(n_4514),
.B(n_3434),
.Y(n_4882)
);

AOI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4508),
.A2(n_3177),
.B(n_3147),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_4484),
.B(n_4070),
.Y(n_4884)
);

O2A1O1Ixp33_ASAP7_75t_L g4885 ( 
.A1(n_4350),
.A2(n_869),
.B(n_870),
.C(n_868),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4577),
.B(n_2340),
.Y(n_4886)
);

AOI21xp5_ASAP7_75t_L g4887 ( 
.A1(n_4508),
.A2(n_3196),
.B(n_3177),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4305),
.Y(n_4888)
);

AOI21xp5_ASAP7_75t_L g4889 ( 
.A1(n_4520),
.A2(n_3196),
.B(n_3177),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4336),
.Y(n_4890)
);

AOI21xp5_ASAP7_75t_L g4891 ( 
.A1(n_4520),
.A2(n_4521),
.B(n_4493),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_SL g4892 ( 
.A(n_4484),
.B(n_4070),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4521),
.A2(n_3255),
.B(n_3196),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4320),
.B(n_2364),
.Y(n_4894)
);

BUFx12f_ASAP7_75t_L g4895 ( 
.A(n_4317),
.Y(n_4895)
);

AOI22xp5_ASAP7_75t_L g4896 ( 
.A1(n_4629),
.A2(n_2369),
.B1(n_2374),
.B2(n_2364),
.Y(n_4896)
);

CKINVDCx20_ASAP7_75t_R g4897 ( 
.A(n_4311),
.Y(n_4897)
);

AOI21x1_ASAP7_75t_L g4898 ( 
.A1(n_4538),
.A2(n_3187),
.B(n_3183),
.Y(n_4898)
);

AOI22x1_ASAP7_75t_L g4899 ( 
.A1(n_4317),
.A2(n_1082),
.B1(n_1084),
.B2(n_1081),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4306),
.Y(n_4900)
);

INVx2_ASAP7_75t_SL g4901 ( 
.A(n_4314),
.Y(n_4901)
);

AND2x4_ASAP7_75t_L g4902 ( 
.A(n_4232),
.B(n_3405),
.Y(n_4902)
);

OAI22xp5_ASAP7_75t_L g4903 ( 
.A1(n_4459),
.A2(n_3255),
.B1(n_3279),
.B2(n_3196),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4338),
.Y(n_4904)
);

NAND2xp33_ASAP7_75t_L g4905 ( 
.A(n_4514),
.B(n_3434),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_4320),
.B(n_3380),
.Y(n_4906)
);

HB1xp67_ASAP7_75t_L g4907 ( 
.A(n_4435),
.Y(n_4907)
);

NAND2xp33_ASAP7_75t_L g4908 ( 
.A(n_4514),
.B(n_3434),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4493),
.B(n_2369),
.Y(n_4909)
);

O2A1O1Ixp33_ASAP7_75t_L g4910 ( 
.A1(n_4528),
.A2(n_870),
.B(n_871),
.C(n_869),
.Y(n_4910)
);

NOR2xp67_ASAP7_75t_L g4911 ( 
.A(n_4437),
.B(n_3405),
.Y(n_4911)
);

AOI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4300),
.A2(n_3279),
.B(n_3255),
.Y(n_4912)
);

O2A1O1Ixp5_ASAP7_75t_L g4913 ( 
.A1(n_4256),
.A2(n_3227),
.B(n_3302),
.C(n_3187),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4609),
.B(n_2374),
.Y(n_4914)
);

NOR2xp67_ASAP7_75t_L g4915 ( 
.A(n_4445),
.B(n_3406),
.Y(n_4915)
);

A2O1A1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_4579),
.A2(n_879),
.B(n_882),
.C(n_871),
.Y(n_4916)
);

BUFx6f_ASAP7_75t_L g4917 ( 
.A(n_4295),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4609),
.B(n_2304),
.Y(n_4918)
);

AOI21xp5_ASAP7_75t_L g4919 ( 
.A1(n_4300),
.A2(n_3279),
.B(n_3255),
.Y(n_4919)
);

NAND3xp33_ASAP7_75t_L g4920 ( 
.A(n_4568),
.B(n_1093),
.C(n_1089),
.Y(n_4920)
);

AOI22xp33_ASAP7_75t_L g4921 ( 
.A1(n_4629),
.A2(n_2755),
.B1(n_2970),
.B2(n_2603),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_4612),
.B(n_2304),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4612),
.B(n_2338),
.Y(n_4923)
);

NOR2xp67_ASAP7_75t_L g4924 ( 
.A(n_4446),
.B(n_3406),
.Y(n_4924)
);

OAI22xp5_ASAP7_75t_L g4925 ( 
.A1(n_4502),
.A2(n_4575),
.B1(n_4590),
.B2(n_4571),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4322),
.B(n_2338),
.Y(n_4926)
);

O2A1O1Ixp33_ASAP7_75t_L g4927 ( 
.A1(n_4528),
.A2(n_882),
.B(n_888),
.C(n_879),
.Y(n_4927)
);

NOR2xp33_ASAP7_75t_L g4928 ( 
.A(n_4282),
.B(n_1094),
.Y(n_4928)
);

A2O1A1Ixp33_ASAP7_75t_L g4929 ( 
.A1(n_4310),
.A2(n_898),
.B(n_900),
.C(n_888),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4513),
.B(n_3388),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4325),
.B(n_2338),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4502),
.B(n_4534),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4309),
.Y(n_4933)
);

BUFx8_ASAP7_75t_L g4934 ( 
.A(n_4313),
.Y(n_4934)
);

OAI22xp5_ASAP7_75t_L g4935 ( 
.A1(n_4575),
.A2(n_3288),
.B1(n_3370),
.B2(n_3279),
.Y(n_4935)
);

OAI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4569),
.A2(n_2970),
.B(n_2755),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_SL g4937 ( 
.A(n_4513),
.B(n_3388),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_SL g4938 ( 
.A(n_4524),
.B(n_3394),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4343),
.B(n_2338),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4353),
.B(n_2107),
.Y(n_4940)
);

OR2x6_ASAP7_75t_SL g4941 ( 
.A(n_4476),
.B(n_1099),
.Y(n_4941)
);

NOR2xp33_ASAP7_75t_SL g4942 ( 
.A(n_4428),
.B(n_3288),
.Y(n_4942)
);

OAI21xp33_ASAP7_75t_L g4943 ( 
.A1(n_4597),
.A2(n_1110),
.B(n_1105),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_SL g4944 ( 
.A(n_4524),
.B(n_3394),
.Y(n_4944)
);

AND2x2_ASAP7_75t_SL g4945 ( 
.A(n_4509),
.B(n_898),
.Y(n_4945)
);

OAI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4298),
.A2(n_2970),
.B(n_2755),
.Y(n_4946)
);

AOI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4564),
.A2(n_4535),
.B(n_4534),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4357),
.B(n_1648),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4564),
.A2(n_3370),
.B(n_3288),
.Y(n_4949)
);

NAND2x1_ASAP7_75t_L g4950 ( 
.A(n_4629),
.B(n_3655),
.Y(n_4950)
);

AOI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4535),
.A2(n_4539),
.B(n_4537),
.Y(n_4951)
);

AOI21xp5_ASAP7_75t_L g4952 ( 
.A1(n_4537),
.A2(n_3370),
.B(n_3288),
.Y(n_4952)
);

NOR2xp33_ASAP7_75t_L g4953 ( 
.A(n_4335),
.B(n_1112),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4374),
.B(n_2107),
.Y(n_4954)
);

AOI21x1_ASAP7_75t_L g4955 ( 
.A1(n_4268),
.A2(n_3302),
.B(n_3227),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4316),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4395),
.B(n_2107),
.Y(n_4957)
);

O2A1O1Ixp33_ASAP7_75t_L g4958 ( 
.A1(n_4586),
.A2(n_901),
.B(n_906),
.C(n_900),
.Y(n_4958)
);

NOR2x1p5_ASAP7_75t_L g4959 ( 
.A(n_4433),
.B(n_2562),
.Y(n_4959)
);

OR2x6_ASAP7_75t_SL g4960 ( 
.A(n_4471),
.B(n_1113),
.Y(n_4960)
);

BUFx12f_ASAP7_75t_L g4961 ( 
.A(n_4313),
.Y(n_4961)
);

AOI22x1_ASAP7_75t_L g4962 ( 
.A1(n_4509),
.A2(n_1115),
.B1(n_1116),
.B2(n_1114),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_SL g4963 ( 
.A(n_4519),
.B(n_3395),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4414),
.B(n_2107),
.Y(n_4964)
);

AO21x1_ASAP7_75t_L g4965 ( 
.A1(n_4241),
.A2(n_906),
.B(n_901),
.Y(n_4965)
);

OAI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4631),
.A2(n_3389),
.B1(n_3422),
.B2(n_3370),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4586),
.B(n_1122),
.Y(n_4967)
);

BUFx6f_ASAP7_75t_L g4968 ( 
.A(n_4313),
.Y(n_4968)
);

AOI21xp5_ASAP7_75t_L g4969 ( 
.A1(n_4539),
.A2(n_3389),
.B(n_3422),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4595),
.A2(n_2970),
.B(n_2755),
.Y(n_4970)
);

AOI21xp5_ASAP7_75t_L g4971 ( 
.A1(n_4541),
.A2(n_4632),
.B(n_4595),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4327),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_SL g4973 ( 
.A(n_4519),
.B(n_3395),
.Y(n_4973)
);

OAI21xp5_ASAP7_75t_L g4974 ( 
.A1(n_4541),
.A2(n_2970),
.B(n_3434),
.Y(n_4974)
);

AND2x2_ASAP7_75t_L g4975 ( 
.A(n_4354),
.B(n_4355),
.Y(n_4975)
);

NOR2xp67_ASAP7_75t_L g4976 ( 
.A(n_4455),
.B(n_3401),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4328),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_SL g4978 ( 
.A(n_4519),
.B(n_3401),
.Y(n_4978)
);

AOI22xp5_ASAP7_75t_L g4979 ( 
.A1(n_4271),
.A2(n_2970),
.B1(n_1128),
.B2(n_1131),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4632),
.A2(n_3422),
.B(n_3389),
.Y(n_4980)
);

AND2x4_ASAP7_75t_L g4981 ( 
.A(n_4232),
.B(n_4261),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_SL g4982 ( 
.A(n_4511),
.B(n_3389),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_SL g4983 ( 
.A(n_4511),
.B(n_3422),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4482),
.B(n_1124),
.Y(n_4984)
);

O2A1O1Ixp5_ASAP7_75t_L g4985 ( 
.A1(n_4503),
.A2(n_3420),
.B(n_2612),
.C(n_2605),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4458),
.Y(n_4986)
);

NOR2xp33_ASAP7_75t_L g4987 ( 
.A(n_4335),
.B(n_4271),
.Y(n_4987)
);

INVxp67_ASAP7_75t_L g4988 ( 
.A(n_4321),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4496),
.B(n_1133),
.Y(n_4989)
);

NOR2xp33_ASAP7_75t_L g4990 ( 
.A(n_4275),
.B(n_1134),
.Y(n_4990)
);

AND2x6_ASAP7_75t_SL g4991 ( 
.A(n_4452),
.B(n_907),
.Y(n_4991)
);

OAI22xp5_ASAP7_75t_L g4992 ( 
.A1(n_4510),
.A2(n_1137),
.B1(n_1139),
.B2(n_1136),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_SL g4993 ( 
.A(n_4232),
.B(n_3123),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4488),
.B(n_4563),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4506),
.B(n_1140),
.Y(n_4995)
);

INVxp67_ASAP7_75t_SL g4996 ( 
.A(n_4456),
.Y(n_4996)
);

INVx1_ASAP7_75t_SL g4997 ( 
.A(n_4522),
.Y(n_4997)
);

AOI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4503),
.A2(n_3148),
.B(n_2987),
.Y(n_4998)
);

NAND2xp5_ASAP7_75t_L g4999 ( 
.A(n_4512),
.B(n_1142),
.Y(n_4999)
);

OAI21xp33_ASAP7_75t_L g5000 ( 
.A1(n_4561),
.A2(n_1145),
.B(n_1144),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4515),
.B(n_1147),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4494),
.B(n_1648),
.Y(n_5002)
);

AO21x1_ASAP7_75t_L g5003 ( 
.A1(n_4561),
.A2(n_914),
.B(n_907),
.Y(n_5003)
);

NAND3xp33_ASAP7_75t_L g5004 ( 
.A(n_4326),
.B(n_1150),
.C(n_1149),
.Y(n_5004)
);

O2A1O1Ixp33_ASAP7_75t_L g5005 ( 
.A1(n_4504),
.A2(n_919),
.B(n_934),
.C(n_914),
.Y(n_5005)
);

CKINVDCx20_ASAP7_75t_R g5006 ( 
.A(n_4340),
.Y(n_5006)
);

AOI21xp5_ASAP7_75t_L g5007 ( 
.A1(n_4504),
.A2(n_3148),
.B(n_2987),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_SL g5008 ( 
.A(n_4261),
.B(n_3123),
.Y(n_5008)
);

INVx2_ASAP7_75t_L g5009 ( 
.A(n_4518),
.Y(n_5009)
);

OAI21x1_ASAP7_75t_L g5010 ( 
.A1(n_4611),
.A2(n_3271),
.B(n_3204),
.Y(n_5010)
);

A2O1A1Ixp33_ASAP7_75t_L g5011 ( 
.A1(n_4261),
.A2(n_934),
.B(n_938),
.C(n_919),
.Y(n_5011)
);

O2A1O1Ixp33_ASAP7_75t_L g5012 ( 
.A1(n_4507),
.A2(n_939),
.B(n_944),
.C(n_938),
.Y(n_5012)
);

AOI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4507),
.A2(n_3148),
.B(n_2987),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4326),
.A2(n_2987),
.B(n_2983),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_4261),
.B(n_3123),
.Y(n_5015)
);

NOR3xp33_ASAP7_75t_L g5016 ( 
.A(n_4462),
.B(n_944),
.C(n_939),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4452),
.A2(n_4510),
.B(n_4474),
.Y(n_5017)
);

NOR2xp33_ASAP7_75t_SL g5018 ( 
.A(n_4428),
.B(n_4432),
.Y(n_5018)
);

A2O1A1Ixp33_ASAP7_75t_L g5019 ( 
.A1(n_4332),
.A2(n_950),
.B(n_952),
.C(n_949),
.Y(n_5019)
);

OAI22xp5_ASAP7_75t_L g5020 ( 
.A1(n_4472),
.A2(n_1159),
.B1(n_1160),
.B2(n_1153),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4349),
.B(n_3300),
.Y(n_5021)
);

A2O1A1Ixp33_ASAP7_75t_L g5022 ( 
.A1(n_4351),
.A2(n_950),
.B(n_952),
.C(n_949),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4358),
.B(n_3300),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4363),
.B(n_3300),
.Y(n_5024)
);

OAI22xp5_ASAP7_75t_L g5025 ( 
.A1(n_4472),
.A2(n_1165),
.B1(n_1169),
.B2(n_1164),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4452),
.A2(n_3373),
.B(n_2987),
.Y(n_5026)
);

INVxp67_ASAP7_75t_L g5027 ( 
.A(n_4342),
.Y(n_5027)
);

AOI21xp5_ASAP7_75t_L g5028 ( 
.A1(n_4474),
.A2(n_3373),
.B(n_2987),
.Y(n_5028)
);

INVx4_ASAP7_75t_L g5029 ( 
.A(n_4438),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4365),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4368),
.B(n_4369),
.Y(n_5031)
);

AOI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4301),
.A2(n_3051),
.B(n_2983),
.Y(n_5032)
);

NOR2xp33_ASAP7_75t_L g5033 ( 
.A(n_4275),
.B(n_1173),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4605),
.B(n_3123),
.Y(n_5034)
);

A2O1A1Ixp33_ASAP7_75t_L g5035 ( 
.A1(n_4375),
.A2(n_961),
.B(n_965),
.C(n_960),
.Y(n_5035)
);

INVx2_ASAP7_75t_SL g5036 ( 
.A(n_4418),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4301),
.A2(n_3051),
.B(n_2983),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4378),
.Y(n_5038)
);

O2A1O1Ixp33_ASAP7_75t_L g5039 ( 
.A1(n_4381),
.A2(n_961),
.B(n_965),
.C(n_960),
.Y(n_5039)
);

AOI21x1_ASAP7_75t_L g5040 ( 
.A1(n_4385),
.A2(n_3420),
.B(n_2532),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4391),
.B(n_3375),
.Y(n_5041)
);

AOI21xp5_ASAP7_75t_L g5042 ( 
.A1(n_4611),
.A2(n_3051),
.B(n_2983),
.Y(n_5042)
);

OAI22xp5_ASAP7_75t_SL g5043 ( 
.A1(n_4472),
.A2(n_986),
.B1(n_993),
.B2(n_971),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4556),
.B(n_1649),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_4396),
.B(n_3375),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4616),
.A2(n_3051),
.B(n_2983),
.Y(n_5046)
);

AOI21xp5_ASAP7_75t_L g5047 ( 
.A1(n_4616),
.A2(n_3051),
.B(n_2983),
.Y(n_5047)
);

AOI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4382),
.A2(n_3097),
.B(n_3051),
.Y(n_5048)
);

CKINVDCx20_ASAP7_75t_R g5049 ( 
.A(n_4438),
.Y(n_5049)
);

INVx3_ASAP7_75t_L g5050 ( 
.A(n_4367),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4400),
.Y(n_5051)
);

O2A1O1Ixp33_ASAP7_75t_L g5052 ( 
.A1(n_4404),
.A2(n_986),
.B(n_993),
.C(n_971),
.Y(n_5052)
);

INVx3_ASAP7_75t_L g5053 ( 
.A(n_4732),
.Y(n_5053)
);

OAI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4689),
.A2(n_4608),
.B(n_4399),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_4832),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4862),
.B(n_4407),
.Y(n_5056)
);

BUFx12f_ASAP7_75t_L g5057 ( 
.A(n_4776),
.Y(n_5057)
);

OAI21x1_ASAP7_75t_L g5058 ( 
.A1(n_4717),
.A2(n_4410),
.B(n_4409),
.Y(n_5058)
);

NAND3xp33_ASAP7_75t_SL g5059 ( 
.A(n_4643),
.B(n_1176),
.C(n_1175),
.Y(n_5059)
);

INVx2_ASAP7_75t_L g5060 ( 
.A(n_4692),
.Y(n_5060)
);

CKINVDCx5p33_ASAP7_75t_R g5061 ( 
.A(n_4683),
.Y(n_5061)
);

A2O1A1Ixp33_ASAP7_75t_L g5062 ( 
.A1(n_4648),
.A2(n_1006),
.B(n_1011),
.C(n_1004),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4862),
.B(n_4789),
.Y(n_5063)
);

AOI21x1_ASAP7_75t_L g5064 ( 
.A1(n_4670),
.A2(n_4419),
.B(n_4411),
.Y(n_5064)
);

OAI21x1_ASAP7_75t_L g5065 ( 
.A1(n_4646),
.A2(n_4423),
.B(n_4420),
.Y(n_5065)
);

BUFx5_ASAP7_75t_L g5066 ( 
.A(n_4878),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_4789),
.B(n_4425),
.Y(n_5067)
);

OAI21x1_ASAP7_75t_L g5068 ( 
.A1(n_4838),
.A2(n_4436),
.B(n_4517),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4705),
.Y(n_5069)
);

AO21x1_ASAP7_75t_L g5070 ( 
.A1(n_4661),
.A2(n_1006),
.B(n_1004),
.Y(n_5070)
);

INVx2_ASAP7_75t_SL g5071 ( 
.A(n_4765),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4854),
.B(n_4526),
.Y(n_5072)
);

AND2x2_ASAP7_75t_L g5073 ( 
.A(n_4975),
.B(n_4634),
.Y(n_5073)
);

INVxp67_ASAP7_75t_L g5074 ( 
.A(n_4690),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_4715),
.B(n_4531),
.Y(n_5075)
);

AOI22xp33_ASAP7_75t_L g5076 ( 
.A1(n_4656),
.A2(n_4399),
.B1(n_4379),
.B2(n_1013),
.Y(n_5076)
);

OA22x2_ASAP7_75t_L g5077 ( 
.A1(n_4997),
.A2(n_4576),
.B1(n_4532),
.B2(n_4547),
.Y(n_5077)
);

AOI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_4664),
.A2(n_4382),
.B(n_4517),
.Y(n_5078)
);

BUFx2_ASAP7_75t_L g5079 ( 
.A(n_4791),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4769),
.Y(n_5080)
);

AO21x1_ASAP7_75t_L g5081 ( 
.A1(n_4910),
.A2(n_1013),
.B(n_1011),
.Y(n_5081)
);

AOI21xp5_ASAP7_75t_L g5082 ( 
.A1(n_4637),
.A2(n_4951),
.B(n_4638),
.Y(n_5082)
);

OAI21x1_ASAP7_75t_L g5083 ( 
.A1(n_4680),
.A2(n_4433),
.B(n_2612),
.Y(n_5083)
);

NAND2x1_ASAP7_75t_L g5084 ( 
.A(n_4669),
.B(n_4527),
.Y(n_5084)
);

AOI21xp5_ASAP7_75t_L g5085 ( 
.A1(n_4891),
.A2(n_4379),
.B(n_4560),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4810),
.Y(n_5086)
);

AOI21xp5_ASAP7_75t_L g5087 ( 
.A1(n_4882),
.A2(n_4560),
.B(n_4281),
.Y(n_5087)
);

OAI21x1_ASAP7_75t_L g5088 ( 
.A1(n_4691),
.A2(n_4572),
.B(n_4527),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4726),
.B(n_4542),
.Y(n_5089)
);

OAI21x1_ASAP7_75t_L g5090 ( 
.A1(n_4693),
.A2(n_4599),
.B(n_4572),
.Y(n_5090)
);

AOI21x1_ASAP7_75t_L g5091 ( 
.A1(n_4707),
.A2(n_4555),
.B(n_4550),
.Y(n_5091)
);

A2O1A1Ixp33_ASAP7_75t_L g5092 ( 
.A1(n_4671),
.A2(n_1017),
.B(n_1023),
.C(n_1016),
.Y(n_5092)
);

NAND2x1_ASAP7_75t_L g5093 ( 
.A(n_4981),
.B(n_4599),
.Y(n_5093)
);

OAI21x1_ASAP7_75t_L g5094 ( 
.A1(n_4998),
.A2(n_4462),
.B(n_2876),
.Y(n_5094)
);

INVx2_ASAP7_75t_SL g5095 ( 
.A(n_4765),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4836),
.Y(n_5096)
);

OAI21x1_ASAP7_75t_L g5097 ( 
.A1(n_5007),
.A2(n_2876),
.B(n_2860),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4842),
.Y(n_5098)
);

INVx5_ASAP7_75t_L g5099 ( 
.A(n_4736),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_4649),
.B(n_4558),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4905),
.A2(n_4281),
.B(n_4370),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_L g5102 ( 
.A(n_4649),
.B(n_4565),
.Y(n_5102)
);

A2O1A1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_4659),
.A2(n_1017),
.B(n_1023),
.C(n_1016),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4908),
.A2(n_4370),
.B(n_3299),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_4932),
.B(n_4621),
.Y(n_5105)
);

AOI21x1_ASAP7_75t_L g5106 ( 
.A1(n_5040),
.A2(n_1650),
.B(n_1649),
.Y(n_5106)
);

CKINVDCx5p33_ASAP7_75t_R g5107 ( 
.A(n_4876),
.Y(n_5107)
);

OAI21x1_ASAP7_75t_L g5108 ( 
.A1(n_5013),
.A2(n_2860),
.B(n_2981),
.Y(n_5108)
);

NAND2xp5_ASAP7_75t_L g5109 ( 
.A(n_4932),
.B(n_4621),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4858),
.Y(n_5110)
);

AOI21xp5_ASAP7_75t_L g5111 ( 
.A1(n_4971),
.A2(n_3299),
.B(n_3097),
.Y(n_5111)
);

AO21x1_ASAP7_75t_L g5112 ( 
.A1(n_4927),
.A2(n_1032),
.B(n_1030),
.Y(n_5112)
);

OAI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_4675),
.A2(n_4774),
.B(n_4920),
.Y(n_5113)
);

OAI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4725),
.A2(n_4405),
.B(n_4403),
.Y(n_5114)
);

BUFx12f_ASAP7_75t_L g5115 ( 
.A(n_4895),
.Y(n_5115)
);

OAI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4744),
.A2(n_4405),
.B(n_4403),
.Y(n_5116)
);

AOI21xp33_ASAP7_75t_L g5117 ( 
.A1(n_5005),
.A2(n_3418),
.B(n_3375),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4888),
.Y(n_5118)
);

OAI21xp5_ASAP7_75t_L g5119 ( 
.A1(n_4647),
.A2(n_4449),
.B(n_4413),
.Y(n_5119)
);

AO21x1_ASAP7_75t_L g5120 ( 
.A1(n_4865),
.A2(n_1032),
.B(n_1030),
.Y(n_5120)
);

OAI21x1_ASAP7_75t_L g5121 ( 
.A1(n_5010),
.A2(n_3001),
.B(n_2981),
.Y(n_5121)
);

BUFx3_ASAP7_75t_L g5122 ( 
.A(n_4897),
.Y(n_5122)
);

AO31x2_ASAP7_75t_L g5123 ( 
.A1(n_4702),
.A2(n_3447),
.A3(n_3451),
.B(n_3446),
.Y(n_5123)
);

OAI21x1_ASAP7_75t_L g5124 ( 
.A1(n_4759),
.A2(n_3003),
.B(n_3001),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_4854),
.B(n_4248),
.Y(n_5125)
);

AOI22xp5_ASAP7_75t_L g5126 ( 
.A1(n_4783),
.A2(n_1178),
.B1(n_1181),
.B2(n_1177),
.Y(n_5126)
);

AOI21xp5_ASAP7_75t_L g5127 ( 
.A1(n_4869),
.A2(n_3299),
.B(n_3097),
.Y(n_5127)
);

BUFx6f_ASAP7_75t_L g5128 ( 
.A(n_4765),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4900),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_SL g5130 ( 
.A(n_4651),
.B(n_4413),
.Y(n_5130)
);

OAI21x1_ASAP7_75t_L g5131 ( 
.A1(n_4697),
.A2(n_3004),
.B(n_3003),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4933),
.Y(n_5132)
);

A2O1A1Ixp33_ASAP7_75t_L g5133 ( 
.A1(n_4687),
.A2(n_1034),
.B(n_1035),
.C(n_1033),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_4907),
.B(n_4293),
.Y(n_5134)
);

NOR2xp67_ASAP7_75t_L g5135 ( 
.A(n_5004),
.B(n_4454),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_4847),
.B(n_4754),
.Y(n_5136)
);

INVx2_ASAP7_75t_SL g5137 ( 
.A(n_4758),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_4653),
.B(n_4248),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_SL g5139 ( 
.A(n_4723),
.B(n_4449),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_SL g5140 ( 
.A1(n_4698),
.A2(n_4432),
.B(n_2658),
.Y(n_5140)
);

NOR2xp33_ASAP7_75t_L g5141 ( 
.A(n_4834),
.B(n_4285),
.Y(n_5141)
);

NOR2xp33_ASAP7_75t_L g5142 ( 
.A(n_4741),
.B(n_4735),
.Y(n_5142)
);

BUFx2_ASAP7_75t_L g5143 ( 
.A(n_4934),
.Y(n_5143)
);

OAI21x1_ASAP7_75t_SL g5144 ( 
.A1(n_4879),
.A2(n_4408),
.B(n_4377),
.Y(n_5144)
);

INVx2_ASAP7_75t_SL g5145 ( 
.A(n_4934),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4956),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_4808),
.B(n_4294),
.Y(n_5147)
);

OAI21x1_ASAP7_75t_L g5148 ( 
.A1(n_4701),
.A2(n_3005),
.B(n_3004),
.Y(n_5148)
);

INVxp67_ASAP7_75t_L g5149 ( 
.A(n_4844),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4972),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_4808),
.B(n_4334),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4743),
.A2(n_3299),
.B(n_3097),
.Y(n_5152)
);

AOI21x1_ASAP7_75t_SL g5153 ( 
.A1(n_4773),
.A2(n_4260),
.B(n_2793),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_4732),
.B(n_4285),
.Y(n_5154)
);

BUFx12f_ASAP7_75t_L g5155 ( 
.A(n_4991),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_4977),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_5030),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5038),
.Y(n_5158)
);

AOI21x1_ASAP7_75t_L g5159 ( 
.A1(n_4863),
.A2(n_1651),
.B(n_1650),
.Y(n_5159)
);

BUFx2_ASAP7_75t_L g5160 ( 
.A(n_4756),
.Y(n_5160)
);

AOI21xp5_ASAP7_75t_SL g5161 ( 
.A1(n_4970),
.A2(n_2658),
.B(n_2653),
.Y(n_5161)
);

OAI21x1_ASAP7_75t_L g5162 ( 
.A1(n_4877),
.A2(n_3014),
.B(n_3005),
.Y(n_5162)
);

OAI22xp5_ASAP7_75t_L g5163 ( 
.A1(n_4945),
.A2(n_1034),
.B1(n_1035),
.B2(n_1033),
.Y(n_5163)
);

OAI21x1_ASAP7_75t_L g5164 ( 
.A1(n_4708),
.A2(n_3015),
.B(n_3014),
.Y(n_5164)
);

AO31x2_ASAP7_75t_L g5165 ( 
.A1(n_5003),
.A2(n_3447),
.A3(n_3451),
.B(n_3446),
.Y(n_5165)
);

OAI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4912),
.A2(n_3018),
.B(n_3015),
.Y(n_5166)
);

NOR2xp33_ASAP7_75t_L g5167 ( 
.A(n_4674),
.B(n_4293),
.Y(n_5167)
);

A2O1A1Ixp33_ASAP7_75t_L g5168 ( 
.A1(n_4635),
.A2(n_1043),
.B(n_1044),
.C(n_1041),
.Y(n_5168)
);

AO21x2_ASAP7_75t_L g5169 ( 
.A1(n_4641),
.A2(n_2532),
.B(n_2529),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_4947),
.A2(n_3299),
.B(n_3097),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4919),
.A2(n_3299),
.B(n_3097),
.Y(n_5171)
);

OAI21x1_ASAP7_75t_L g5172 ( 
.A1(n_4770),
.A2(n_3019),
.B(n_3018),
.Y(n_5172)
);

AOI21xp5_ASAP7_75t_L g5173 ( 
.A1(n_4739),
.A2(n_3372),
.B(n_3304),
.Y(n_5173)
);

AO21x1_ASAP7_75t_L g5174 ( 
.A1(n_5012),
.A2(n_1043),
.B(n_1041),
.Y(n_5174)
);

INVx2_ASAP7_75t_SL g5175 ( 
.A(n_4778),
.Y(n_5175)
);

OAI21x1_ASAP7_75t_L g5176 ( 
.A1(n_4772),
.A2(n_3022),
.B(n_3019),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5051),
.Y(n_5177)
);

NOR2xp33_ASAP7_75t_L g5178 ( 
.A(n_4960),
.B(n_4941),
.Y(n_5178)
);

OAI21xp5_ASAP7_75t_L g5179 ( 
.A1(n_4712),
.A2(n_3665),
.B(n_3655),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_4898),
.A2(n_3024),
.B(n_3022),
.Y(n_5180)
);

INVx2_ASAP7_75t_SL g5181 ( 
.A(n_4864),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4751),
.B(n_4645),
.Y(n_5182)
);

OAI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_4737),
.A2(n_3665),
.B(n_3655),
.Y(n_5183)
);

BUFx6f_ASAP7_75t_L g5184 ( 
.A(n_4864),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_4645),
.B(n_4294),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_4657),
.B(n_4334),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_4996),
.B(n_4416),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5031),
.Y(n_5188)
);

AOI21xp5_ASAP7_75t_L g5189 ( 
.A1(n_4667),
.A2(n_3372),
.B(n_3304),
.Y(n_5189)
);

OAI22x1_ASAP7_75t_L g5190 ( 
.A1(n_4749),
.A2(n_4424),
.B1(n_1047),
.B2(n_1048),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4639),
.B(n_4367),
.Y(n_5191)
);

OAI21x1_ASAP7_75t_L g5192 ( 
.A1(n_4761),
.A2(n_3028),
.B(n_3024),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5031),
.Y(n_5193)
);

INVx5_ASAP7_75t_L g5194 ( 
.A(n_4736),
.Y(n_5194)
);

AOI21xp5_ASAP7_75t_SL g5195 ( 
.A1(n_4709),
.A2(n_4859),
.B(n_4757),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_4667),
.A2(n_3372),
.B(n_3304),
.Y(n_5196)
);

AOI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_4633),
.A2(n_3372),
.B(n_3304),
.Y(n_5197)
);

AOI22xp5_ASAP7_75t_L g5198 ( 
.A1(n_4752),
.A2(n_1187),
.B1(n_1190),
.B2(n_1185),
.Y(n_5198)
);

OR2x6_ASAP7_75t_L g5199 ( 
.A(n_5017),
.B(n_4367),
.Y(n_5199)
);

OAI22x1_ASAP7_75t_L g5200 ( 
.A1(n_4782),
.A2(n_1047),
.B1(n_1048),
.B2(n_1044),
.Y(n_5200)
);

OAI22xp5_ASAP7_75t_L g5201 ( 
.A1(n_5043),
.A2(n_1056),
.B1(n_1064),
.B2(n_1051),
.Y(n_5201)
);

BUFx6f_ASAP7_75t_L g5202 ( 
.A(n_4864),
.Y(n_5202)
);

AOI21xp5_ASAP7_75t_L g5203 ( 
.A1(n_4633),
.A2(n_3372),
.B(n_3304),
.Y(n_5203)
);

OAI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_4925),
.A2(n_3665),
.B(n_3655),
.Y(n_5204)
);

OR2x2_ASAP7_75t_L g5205 ( 
.A(n_4650),
.B(n_1645),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_4639),
.B(n_4371),
.Y(n_5206)
);

AND2x4_ASAP7_75t_L g5207 ( 
.A(n_4981),
.B(n_4371),
.Y(n_5207)
);

AOI21xp33_ASAP7_75t_L g5208 ( 
.A1(n_4958),
.A2(n_3418),
.B(n_1056),
.Y(n_5208)
);

A2O1A1Ixp33_ASAP7_75t_L g5209 ( 
.A1(n_4679),
.A2(n_1064),
.B(n_1067),
.C(n_1051),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_4652),
.B(n_4371),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4633),
.A2(n_3304),
.B(n_3372),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5021),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_SL g5213 ( 
.A(n_4736),
.B(n_4388),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5021),
.Y(n_5214)
);

AOI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_4946),
.A2(n_3373),
.B(n_2812),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_SL g5216 ( 
.A(n_4736),
.B(n_4388),
.Y(n_5216)
);

AOI221x1_ASAP7_75t_L g5217 ( 
.A1(n_4678),
.A2(n_1070),
.B1(n_1074),
.B2(n_1069),
.C(n_1067),
.Y(n_5217)
);

AND2x2_ASAP7_75t_SL g5218 ( 
.A(n_4846),
.B(n_4388),
.Y(n_5218)
);

AO21x1_ASAP7_75t_L g5219 ( 
.A1(n_4992),
.A2(n_1070),
.B(n_1069),
.Y(n_5219)
);

NOR2xp33_ASAP7_75t_L g5220 ( 
.A(n_4771),
.B(n_1191),
.Y(n_5220)
);

AOI21xp5_ASAP7_75t_SL g5221 ( 
.A1(n_5011),
.A2(n_2667),
.B(n_2658),
.Y(n_5221)
);

BUFx3_ASAP7_75t_L g5222 ( 
.A(n_5006),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4853),
.A2(n_3028),
.B(n_2529),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4640),
.B(n_1193),
.Y(n_5224)
);

OAI21x1_ASAP7_75t_L g5225 ( 
.A1(n_4820),
.A2(n_2812),
.B(n_2808),
.Y(n_5225)
);

OAI21xp5_ASAP7_75t_SL g5226 ( 
.A1(n_4803),
.A2(n_4768),
.B(n_4733),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_4640),
.B(n_1196),
.Y(n_5227)
);

AOI21xp33_ASAP7_75t_L g5228 ( 
.A1(n_4965),
.A2(n_3418),
.B(n_1086),
.Y(n_5228)
);

NAND2xp5_ASAP7_75t_L g5229 ( 
.A(n_4650),
.B(n_1074),
.Y(n_5229)
);

OA22x2_ASAP7_75t_L g5230 ( 
.A1(n_4713),
.A2(n_1087),
.B1(n_1088),
.B2(n_1086),
.Y(n_5230)
);

BUFx6f_ASAP7_75t_L g5231 ( 
.A(n_4871),
.Y(n_5231)
);

OAI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_4826),
.A2(n_1088),
.B1(n_1090),
.B2(n_1087),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5023),
.Y(n_5233)
);

AO21x1_ASAP7_75t_L g5234 ( 
.A1(n_4706),
.A2(n_4728),
.B(n_4672),
.Y(n_5234)
);

AOI21xp5_ASAP7_75t_L g5235 ( 
.A1(n_5014),
.A2(n_3373),
.B(n_2814),
.Y(n_5235)
);

OAI21x1_ASAP7_75t_L g5236 ( 
.A1(n_4821),
.A2(n_2814),
.B(n_2808),
.Y(n_5236)
);

NAND2xp5_ASAP7_75t_L g5237 ( 
.A(n_4662),
.B(n_1090),
.Y(n_5237)
);

AOI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_5032),
.A2(n_3373),
.B(n_2825),
.Y(n_5238)
);

NAND2x1p5_ASAP7_75t_L g5239 ( 
.A(n_4950),
.B(n_3368),
.Y(n_5239)
);

INVx3_ASAP7_75t_L g5240 ( 
.A(n_4722),
.Y(n_5240)
);

AO31x2_ASAP7_75t_L g5241 ( 
.A1(n_5026),
.A2(n_2825),
.A3(n_2817),
.B(n_2616),
.Y(n_5241)
);

AOI21xp5_ASAP7_75t_L g5242 ( 
.A1(n_5037),
.A2(n_3373),
.B(n_2817),
.Y(n_5242)
);

AOI21xp33_ASAP7_75t_L g5243 ( 
.A1(n_4860),
.A2(n_1098),
.B(n_1095),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_4987),
.B(n_1095),
.Y(n_5244)
);

AO21x2_ASAP7_75t_L g5245 ( 
.A1(n_4840),
.A2(n_1101),
.B(n_1098),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_4974),
.A2(n_3239),
.B(n_3233),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_5023),
.Y(n_5247)
);

OAI21x1_ASAP7_75t_L g5248 ( 
.A1(n_4780),
.A2(n_2651),
.B(n_2633),
.Y(n_5248)
);

NAND2xp5_ASAP7_75t_L g5249 ( 
.A(n_4662),
.B(n_1101),
.Y(n_5249)
);

AO31x2_ASAP7_75t_L g5250 ( 
.A1(n_5042),
.A2(n_2616),
.A3(n_2610),
.B(n_1104),
.Y(n_5250)
);

OAI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_4724),
.A2(n_3665),
.B(n_3745),
.Y(n_5251)
);

OAI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_4766),
.A2(n_3665),
.B(n_3745),
.Y(n_5252)
);

OAI21x1_ASAP7_75t_L g5253 ( 
.A1(n_4781),
.A2(n_2651),
.B(n_2633),
.Y(n_5253)
);

AND2x4_ASAP7_75t_L g5254 ( 
.A(n_4727),
.B(n_1645),
.Y(n_5254)
);

OAI21x1_ASAP7_75t_L g5255 ( 
.A1(n_4787),
.A2(n_2651),
.B(n_2633),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_4747),
.B(n_1103),
.Y(n_5256)
);

OR2x6_ASAP7_75t_L g5257 ( 
.A(n_4727),
.B(n_3136),
.Y(n_5257)
);

NOR2xp33_ASAP7_75t_L g5258 ( 
.A(n_4682),
.B(n_1197),
.Y(n_5258)
);

OAI21xp5_ASAP7_75t_L g5259 ( 
.A1(n_4636),
.A2(n_3746),
.B(n_3745),
.Y(n_5259)
);

BUFx6f_ASAP7_75t_L g5260 ( 
.A(n_4871),
.Y(n_5260)
);

NAND2x1p5_ASAP7_75t_L g5261 ( 
.A(n_4993),
.B(n_3351),
.Y(n_5261)
);

OAI21x1_ASAP7_75t_L g5262 ( 
.A1(n_4793),
.A2(n_4852),
.B(n_4829),
.Y(n_5262)
);

INVx2_ASAP7_75t_L g5263 ( 
.A(n_4654),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4663),
.B(n_1103),
.Y(n_5264)
);

INVx6_ASAP7_75t_L g5265 ( 
.A(n_4961),
.Y(n_5265)
);

OAI21x1_ASAP7_75t_L g5266 ( 
.A1(n_4955),
.A2(n_2690),
.B(n_2666),
.Y(n_5266)
);

O2A1O1Ixp33_ASAP7_75t_L g5267 ( 
.A1(n_4916),
.A2(n_4943),
.B(n_4730),
.C(n_4929),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_4663),
.B(n_1104),
.Y(n_5268)
);

OAI21x1_ASAP7_75t_L g5269 ( 
.A1(n_5046),
.A2(n_2690),
.B(n_2666),
.Y(n_5269)
);

OAI21x1_ASAP7_75t_L g5270 ( 
.A1(n_5047),
.A2(n_2690),
.B(n_2666),
.Y(n_5270)
);

A2O1A1Ixp33_ASAP7_75t_L g5271 ( 
.A1(n_5000),
.A2(n_1109),
.B(n_1111),
.C(n_1107),
.Y(n_5271)
);

OAI22xp5_ASAP7_75t_L g5272 ( 
.A1(n_4874),
.A2(n_1109),
.B1(n_1111),
.B2(n_1107),
.Y(n_5272)
);

OAI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_4714),
.A2(n_3746),
.B(n_3745),
.Y(n_5273)
);

INVx4_ASAP7_75t_L g5274 ( 
.A(n_4871),
.Y(n_5274)
);

BUFx3_ASAP7_75t_L g5275 ( 
.A(n_5049),
.Y(n_5275)
);

OAI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4985),
.A2(n_2712),
.B(n_2704),
.Y(n_5276)
);

INVxp67_ASAP7_75t_SL g5277 ( 
.A(n_5024),
.Y(n_5277)
);

INVx2_ASAP7_75t_SL g5278 ( 
.A(n_4917),
.Y(n_5278)
);

OAI21x1_ASAP7_75t_L g5279 ( 
.A1(n_4949),
.A2(n_2712),
.B(n_2704),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_4666),
.B(n_1117),
.Y(n_5280)
);

NAND2xp5_ASAP7_75t_L g5281 ( 
.A(n_4666),
.B(n_1117),
.Y(n_5281)
);

AO31x2_ASAP7_75t_L g5282 ( 
.A1(n_5024),
.A2(n_1123),
.A3(n_1127),
.B(n_1118),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_L g5283 ( 
.A1(n_4883),
.A2(n_3239),
.B(n_3233),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4696),
.A2(n_2712),
.B(n_2704),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_5041),
.B(n_1118),
.Y(n_5285)
);

AOI21xp5_ASAP7_75t_L g5286 ( 
.A1(n_4887),
.A2(n_3242),
.B(n_3240),
.Y(n_5286)
);

AO31x2_ASAP7_75t_L g5287 ( 
.A1(n_5041),
.A2(n_1127),
.A3(n_1129),
.B(n_1123),
.Y(n_5287)
);

O2A1O1Ixp5_ASAP7_75t_L g5288 ( 
.A1(n_4802),
.A2(n_1132),
.B(n_1135),
.C(n_1129),
.Y(n_5288)
);

AO21x1_ASAP7_75t_L g5289 ( 
.A1(n_4848),
.A2(n_1135),
.B(n_1132),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_4889),
.A2(n_4952),
.B(n_4893),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5045),
.B(n_1138),
.Y(n_5291)
);

OAI21x1_ASAP7_75t_L g5292 ( 
.A1(n_4696),
.A2(n_4913),
.B(n_4969),
.Y(n_5292)
);

OAI21xp5_ASAP7_75t_L g5293 ( 
.A1(n_4704),
.A2(n_3746),
.B(n_3745),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_5045),
.B(n_1138),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_SL g5295 ( 
.A(n_4755),
.B(n_1667),
.Y(n_5295)
);

OAI21x1_ASAP7_75t_L g5296 ( 
.A1(n_4861),
.A2(n_2815),
.B(n_2776),
.Y(n_5296)
);

AOI21xp5_ASAP7_75t_L g5297 ( 
.A1(n_5028),
.A2(n_3242),
.B(n_3240),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4936),
.A2(n_3261),
.B(n_3256),
.Y(n_5298)
);

BUFx2_ASAP7_75t_L g5299 ( 
.A(n_4839),
.Y(n_5299)
);

A2O1A1Ixp33_ASAP7_75t_L g5300 ( 
.A1(n_5016),
.A2(n_1143),
.B(n_1151),
.C(n_1141),
.Y(n_5300)
);

AOI22xp5_ASAP7_75t_L g5301 ( 
.A1(n_4796),
.A2(n_1206),
.B1(n_1209),
.B2(n_1202),
.Y(n_5301)
);

OAI21xp5_ASAP7_75t_L g5302 ( 
.A1(n_4804),
.A2(n_3746),
.B(n_1143),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_4784),
.B(n_4994),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4700),
.Y(n_5304)
);

AO31x2_ASAP7_75t_L g5305 ( 
.A1(n_4716),
.A2(n_1151),
.A3(n_1152),
.B(n_1141),
.Y(n_5305)
);

AOI21xp33_ASAP7_75t_L g5306 ( 
.A1(n_5039),
.A2(n_1154),
.B(n_1152),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_L g5307 ( 
.A1(n_4980),
.A2(n_5048),
.B(n_5015),
.Y(n_5307)
);

AOI22xp5_ASAP7_75t_L g5308 ( 
.A1(n_4813),
.A2(n_1214),
.B1(n_1218),
.B2(n_1216),
.Y(n_5308)
);

BUFx3_ASAP7_75t_L g5309 ( 
.A(n_4786),
.Y(n_5309)
);

AOI21xp5_ASAP7_75t_L g5310 ( 
.A1(n_5008),
.A2(n_4942),
.B(n_4668),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_4785),
.Y(n_5311)
);

INVx2_ASAP7_75t_SL g5312 ( 
.A(n_4917),
.Y(n_5312)
);

OAI21x1_ASAP7_75t_L g5313 ( 
.A1(n_4841),
.A2(n_2815),
.B(n_2776),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_4809),
.B(n_1154),
.Y(n_5314)
);

INVx4_ASAP7_75t_L g5315 ( 
.A(n_4917),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_4809),
.B(n_1156),
.Y(n_5316)
);

A2O1A1Ixp33_ASAP7_75t_L g5317 ( 
.A1(n_5052),
.A2(n_1157),
.B(n_1158),
.C(n_1156),
.Y(n_5317)
);

AOI21xp5_ASAP7_75t_L g5318 ( 
.A1(n_4668),
.A2(n_3261),
.B(n_3256),
.Y(n_5318)
);

AOI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_4727),
.A2(n_3269),
.B(n_3266),
.Y(n_5319)
);

BUFx6f_ASAP7_75t_SL g5320 ( 
.A(n_4750),
.Y(n_5320)
);

AND2x6_ASAP7_75t_SL g5321 ( 
.A(n_4665),
.B(n_1157),
.Y(n_5321)
);

AOI21x1_ASAP7_75t_L g5322 ( 
.A1(n_4976),
.A2(n_1652),
.B(n_1651),
.Y(n_5322)
);

OAI21xp5_ASAP7_75t_L g5323 ( 
.A1(n_4896),
.A2(n_3746),
.B(n_1162),
.Y(n_5323)
);

A2O1A1Ixp33_ASAP7_75t_L g5324 ( 
.A1(n_4835),
.A2(n_4843),
.B(n_4979),
.C(n_4738),
.Y(n_5324)
);

OAI22xp5_ASAP7_75t_L g5325 ( 
.A1(n_4886),
.A2(n_1162),
.B1(n_1163),
.B2(n_1158),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_4699),
.B(n_1213),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_4710),
.A2(n_2815),
.B(n_2776),
.Y(n_5327)
);

BUFx2_ASAP7_75t_L g5328 ( 
.A(n_4722),
.Y(n_5328)
);

OAI21x1_ASAP7_75t_L g5329 ( 
.A1(n_4710),
.A2(n_2820),
.B(n_2816),
.Y(n_5329)
);

OAI22xp5_ASAP7_75t_L g5330 ( 
.A1(n_4875),
.A2(n_1167),
.B1(n_1171),
.B2(n_1163),
.Y(n_5330)
);

INVx2_ASAP7_75t_L g5331 ( 
.A(n_4797),
.Y(n_5331)
);

OAI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_4814),
.A2(n_1171),
.B(n_1167),
.Y(n_5332)
);

INVxp67_ASAP7_75t_L g5333 ( 
.A(n_4807),
.Y(n_5333)
);

AOI22xp33_ASAP7_75t_L g5334 ( 
.A1(n_4855),
.A2(n_1179),
.B1(n_1180),
.B2(n_1172),
.Y(n_5334)
);

OAI21x1_ASAP7_75t_L g5335 ( 
.A1(n_4734),
.A2(n_2820),
.B(n_2816),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4694),
.B(n_1219),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_4982),
.A2(n_3269),
.B(n_3266),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_4805),
.Y(n_5338)
);

OAI21x1_ASAP7_75t_L g5339 ( 
.A1(n_4734),
.A2(n_2820),
.B(n_2816),
.Y(n_5339)
);

INVx3_ASAP7_75t_L g5340 ( 
.A(n_4762),
.Y(n_5340)
);

OAI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_4815),
.A2(n_1179),
.B(n_1172),
.Y(n_5341)
);

INVxp67_ASAP7_75t_SL g5342 ( 
.A(n_4816),
.Y(n_5342)
);

OAI22xp5_ASAP7_75t_L g5343 ( 
.A1(n_4881),
.A2(n_1182),
.B1(n_1183),
.B2(n_1180),
.Y(n_5343)
);

OAI21x1_ASAP7_75t_L g5344 ( 
.A1(n_4746),
.A2(n_2857),
.B(n_2830),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_4824),
.Y(n_5345)
);

INVx2_ASAP7_75t_L g5346 ( 
.A(n_4845),
.Y(n_5346)
);

OAI21x1_ASAP7_75t_SL g5347 ( 
.A1(n_4794),
.A2(n_1183),
.B(n_1182),
.Y(n_5347)
);

BUFx3_ASAP7_75t_L g5348 ( 
.A(n_4901),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_L g5349 ( 
.A(n_4695),
.B(n_1223),
.Y(n_5349)
);

AOI21x1_ASAP7_75t_L g5350 ( 
.A1(n_4655),
.A2(n_1657),
.B(n_1652),
.Y(n_5350)
);

AO31x2_ASAP7_75t_L g5351 ( 
.A1(n_4935),
.A2(n_1186),
.A3(n_1198),
.B(n_1184),
.Y(n_5351)
);

AND3x4_ASAP7_75t_L g5352 ( 
.A(n_4711),
.B(n_1670),
.C(n_1667),
.Y(n_5352)
);

AND2x4_ASAP7_75t_L g5353 ( 
.A(n_4763),
.B(n_1670),
.Y(n_5353)
);

OAI21x1_ASAP7_75t_L g5354 ( 
.A1(n_4746),
.A2(n_2857),
.B(n_2830),
.Y(n_5354)
);

NAND2xp5_ASAP7_75t_L g5355 ( 
.A(n_4870),
.B(n_1224),
.Y(n_5355)
);

OAI21x1_ASAP7_75t_L g5356 ( 
.A1(n_4801),
.A2(n_2857),
.B(n_2830),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_4644),
.B(n_1184),
.Y(n_5357)
);

A2O1A1Ixp33_ASAP7_75t_L g5358 ( 
.A1(n_4885),
.A2(n_1198),
.B(n_1199),
.C(n_1186),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_4644),
.B(n_4928),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_4890),
.B(n_1226),
.Y(n_5360)
);

AO31x2_ASAP7_75t_L g5361 ( 
.A1(n_4903),
.A2(n_1200),
.A3(n_1205),
.B(n_1199),
.Y(n_5361)
);

AND2x4_ASAP7_75t_L g5362 ( 
.A(n_4762),
.B(n_1680),
.Y(n_5362)
);

AND2x4_ASAP7_75t_L g5363 ( 
.A(n_4880),
.B(n_1680),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_4983),
.A2(n_3280),
.B(n_3270),
.Y(n_5364)
);

OAI21x1_ASAP7_75t_L g5365 ( 
.A1(n_4822),
.A2(n_2866),
.B(n_2863),
.Y(n_5365)
);

NAND2xp5_ASAP7_75t_L g5366 ( 
.A(n_4904),
.B(n_1230),
.Y(n_5366)
);

AOI21xp5_ASAP7_75t_L g5367 ( 
.A1(n_4906),
.A2(n_3280),
.B(n_3270),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_4986),
.B(n_1232),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_5009),
.B(n_4720),
.Y(n_5369)
);

NAND2xp5_ASAP7_75t_SL g5370 ( 
.A(n_5018),
.B(n_1685),
.Y(n_5370)
);

AND2x6_ASAP7_75t_SL g5371 ( 
.A(n_4800),
.B(n_1200),
.Y(n_5371)
);

NOR2xp33_ASAP7_75t_L g5372 ( 
.A(n_4812),
.B(n_1235),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_4713),
.B(n_1205),
.Y(n_5373)
);

OAI21x1_ASAP7_75t_L g5374 ( 
.A1(n_4830),
.A2(n_2866),
.B(n_2863),
.Y(n_5374)
);

BUFx12f_ASAP7_75t_L g5375 ( 
.A(n_5036),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_4721),
.B(n_1236),
.Y(n_5376)
);

CKINVDCx20_ASAP7_75t_R g5377 ( 
.A(n_4703),
.Y(n_5377)
);

BUFx12f_ASAP7_75t_L g5378 ( 
.A(n_4750),
.Y(n_5378)
);

AND2x2_ASAP7_75t_L g5379 ( 
.A(n_4867),
.B(n_1208),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_4816),
.B(n_1208),
.Y(n_5380)
);

AOI21xp5_ASAP7_75t_L g5381 ( 
.A1(n_4872),
.A2(n_3294),
.B(n_3292),
.Y(n_5381)
);

AND2x2_ASAP7_75t_L g5382 ( 
.A(n_4867),
.B(n_1210),
.Y(n_5382)
);

NAND2xp5_ASAP7_75t_L g5383 ( 
.A(n_4817),
.B(n_1210),
.Y(n_5383)
);

AOI21x1_ASAP7_75t_L g5384 ( 
.A1(n_4911),
.A2(n_1658),
.B(n_1657),
.Y(n_5384)
);

AOI21xp33_ASAP7_75t_L g5385 ( 
.A1(n_4779),
.A2(n_4894),
.B(n_4909),
.Y(n_5385)
);

OA21x2_ASAP7_75t_L g5386 ( 
.A1(n_4884),
.A2(n_1659),
.B(n_1658),
.Y(n_5386)
);

AOI21xp5_ASAP7_75t_L g5387 ( 
.A1(n_4892),
.A2(n_3294),
.B(n_3292),
.Y(n_5387)
);

A2O1A1Ixp33_ASAP7_75t_L g5388 ( 
.A1(n_4767),
.A2(n_1217),
.B(n_1222),
.C(n_1215),
.Y(n_5388)
);

OR2x2_ASAP7_75t_L g5389 ( 
.A(n_4792),
.B(n_1685),
.Y(n_5389)
);

BUFx6f_ASAP7_75t_L g5390 ( 
.A(n_4968),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_4817),
.B(n_1215),
.Y(n_5391)
);

OAI21xp5_ASAP7_75t_L g5392 ( 
.A1(n_4827),
.A2(n_4967),
.B(n_4760),
.Y(n_5392)
);

BUFx2_ASAP7_75t_SL g5393 ( 
.A(n_4660),
.Y(n_5393)
);

OAI21x1_ASAP7_75t_L g5394 ( 
.A1(n_4788),
.A2(n_2866),
.B(n_2863),
.Y(n_5394)
);

INVx1_ASAP7_75t_SL g5395 ( 
.A(n_4779),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_4818),
.B(n_1217),
.Y(n_5396)
);

AOI21x1_ASAP7_75t_L g5397 ( 
.A1(n_4915),
.A2(n_1660),
.B(n_1659),
.Y(n_5397)
);

OAI21xp5_ASAP7_75t_L g5398 ( 
.A1(n_4851),
.A2(n_1229),
.B(n_1222),
.Y(n_5398)
);

AOI221x1_ASAP7_75t_L g5399 ( 
.A1(n_5019),
.A2(n_1240),
.B1(n_1233),
.B2(n_1229),
.C(n_1660),
.Y(n_5399)
);

OAI21x1_ASAP7_75t_L g5400 ( 
.A1(n_4788),
.A2(n_2891),
.B(n_2875),
.Y(n_5400)
);

NAND2xp5_ASAP7_75t_L g5401 ( 
.A(n_4818),
.B(n_1233),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4948),
.Y(n_5402)
);

AOI21xp33_ASAP7_75t_L g5403 ( 
.A1(n_4918),
.A2(n_4923),
.B(n_4922),
.Y(n_5403)
);

AOI21xp5_ASAP7_75t_L g5404 ( 
.A1(n_4914),
.A2(n_3312),
.B(n_3307),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_4857),
.A2(n_3312),
.B(n_3307),
.Y(n_5405)
);

CKINVDCx5p33_ASAP7_75t_R g5406 ( 
.A(n_4660),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_4777),
.B(n_1238),
.Y(n_5407)
);

BUFx2_ASAP7_75t_L g5408 ( 
.A(n_4880),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_4794),
.B(n_1242),
.Y(n_5409)
);

AOI21xp33_ASAP7_75t_L g5410 ( 
.A1(n_4857),
.A2(n_4873),
.B(n_4790),
.Y(n_5410)
);

NAND2xp5_ASAP7_75t_L g5411 ( 
.A(n_4823),
.B(n_1243),
.Y(n_5411)
);

AOI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_4873),
.A2(n_3318),
.B(n_3314),
.Y(n_5412)
);

NOR2x1_ASAP7_75t_SL g5413 ( 
.A(n_4718),
.B(n_4790),
.Y(n_5413)
);

OAI22xp5_ASAP7_75t_L g5414 ( 
.A1(n_4806),
.A2(n_4740),
.B1(n_4729),
.B2(n_5035),
.Y(n_5414)
);

INVxp67_ASAP7_75t_SL g5415 ( 
.A(n_4850),
.Y(n_5415)
);

OAI21x1_ASAP7_75t_L g5416 ( 
.A1(n_4850),
.A2(n_2891),
.B(n_2875),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_L g5417 ( 
.A(n_4823),
.B(n_1247),
.Y(n_5417)
);

AO21x1_ASAP7_75t_L g5418 ( 
.A1(n_4963),
.A2(n_1240),
.B(n_1662),
.Y(n_5418)
);

OAI21x1_ASAP7_75t_L g5419 ( 
.A1(n_4825),
.A2(n_2891),
.B(n_2875),
.Y(n_5419)
);

BUFx3_ASAP7_75t_L g5420 ( 
.A(n_4968),
.Y(n_5420)
);

BUFx6f_ASAP7_75t_L g5421 ( 
.A(n_4968),
.Y(n_5421)
);

OAI21x1_ASAP7_75t_SL g5422 ( 
.A1(n_4825),
.A2(n_1699),
.B(n_1690),
.Y(n_5422)
);

AOI21xp5_ASAP7_75t_L g5423 ( 
.A1(n_4866),
.A2(n_3318),
.B(n_3314),
.Y(n_5423)
);

AOI21x1_ASAP7_75t_L g5424 ( 
.A1(n_4924),
.A2(n_5034),
.B(n_4978),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_4831),
.B(n_1249),
.Y(n_5425)
);

OAI21x1_ASAP7_75t_L g5426 ( 
.A1(n_4831),
.A2(n_2914),
.B(n_2892),
.Y(n_5426)
);

OAI21x1_ASAP7_75t_L g5427 ( 
.A1(n_4833),
.A2(n_2914),
.B(n_2892),
.Y(n_5427)
);

OAI21xp5_ASAP7_75t_L g5428 ( 
.A1(n_4798),
.A2(n_3291),
.B(n_2564),
.Y(n_5428)
);

NAND2xp5_ASAP7_75t_L g5429 ( 
.A(n_4833),
.B(n_1251),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_4731),
.Y(n_5430)
);

OAI21xp5_ASAP7_75t_L g5431 ( 
.A1(n_4684),
.A2(n_3291),
.B(n_2563),
.Y(n_5431)
);

OAI21x1_ASAP7_75t_L g5432 ( 
.A1(n_4837),
.A2(n_2914),
.B(n_2892),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_4837),
.B(n_1690),
.Y(n_5433)
);

NOR2x1_ASAP7_75t_SL g5434 ( 
.A(n_4849),
.B(n_3136),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_4731),
.Y(n_5435)
);

OAI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_5022),
.A2(n_3291),
.B(n_1669),
.Y(n_5436)
);

AOI21xp5_ASAP7_75t_L g5437 ( 
.A1(n_4921),
.A2(n_3331),
.B(n_3328),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5050),
.Y(n_5438)
);

BUFx6f_ASAP7_75t_L g5439 ( 
.A(n_5050),
.Y(n_5439)
);

AOI21x1_ASAP7_75t_L g5440 ( 
.A1(n_4973),
.A2(n_1669),
.B(n_1662),
.Y(n_5440)
);

AOI21xp5_ASAP7_75t_L g5441 ( 
.A1(n_4849),
.A2(n_3331),
.B(n_3328),
.Y(n_5441)
);

AOI21xp5_ASAP7_75t_L g5442 ( 
.A1(n_4676),
.A2(n_3341),
.B(n_3334),
.Y(n_5442)
);

OAI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_4775),
.A2(n_4688),
.B(n_4742),
.Y(n_5443)
);

OAI21xp5_ASAP7_75t_L g5444 ( 
.A1(n_4745),
.A2(n_3291),
.B(n_1679),
.Y(n_5444)
);

OAI21x1_ASAP7_75t_L g5445 ( 
.A1(n_4856),
.A2(n_2941),
.B(n_3035),
.Y(n_5445)
);

AOI21xp5_ASAP7_75t_L g5446 ( 
.A1(n_4677),
.A2(n_3341),
.B(n_3334),
.Y(n_5446)
);

AOI21xp5_ASAP7_75t_L g5447 ( 
.A1(n_4681),
.A2(n_3358),
.B(n_3348),
.Y(n_5447)
);

O2A1O1Ixp5_ASAP7_75t_L g5448 ( 
.A1(n_4930),
.A2(n_1679),
.B(n_1687),
.C(n_1673),
.Y(n_5448)
);

CKINVDCx16_ASAP7_75t_R g5449 ( 
.A(n_4658),
.Y(n_5449)
);

AOI21xp5_ASAP7_75t_L g5450 ( 
.A1(n_4686),
.A2(n_3358),
.B(n_3348),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_5002),
.B(n_1699),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_5044),
.B(n_1708),
.Y(n_5452)
);

INVx4_ASAP7_75t_L g5453 ( 
.A(n_5029),
.Y(n_5453)
);

AOI21xp5_ASAP7_75t_L g5454 ( 
.A1(n_4966),
.A2(n_3359),
.B(n_2355),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4926),
.Y(n_5455)
);

OAI21x1_ASAP7_75t_L g5456 ( 
.A1(n_4748),
.A2(n_2941),
.B(n_3035),
.Y(n_5456)
);

OAI21x1_ASAP7_75t_L g5457 ( 
.A1(n_4939),
.A2(n_2941),
.B(n_3052),
.Y(n_5457)
);

AOI21xp5_ASAP7_75t_L g5458 ( 
.A1(n_4937),
.A2(n_4944),
.B(n_4938),
.Y(n_5458)
);

OAI21xp5_ASAP7_75t_L g5459 ( 
.A1(n_5113),
.A2(n_4764),
.B(n_4685),
.Y(n_5459)
);

AO31x2_ASAP7_75t_L g5460 ( 
.A1(n_5290),
.A2(n_5029),
.A3(n_4931),
.B(n_4954),
.Y(n_5460)
);

AO22x1_ASAP7_75t_L g5461 ( 
.A1(n_5113),
.A2(n_4953),
.B1(n_5033),
.B2(n_4990),
.Y(n_5461)
);

NOR2xp33_ASAP7_75t_L g5462 ( 
.A(n_5149),
.B(n_4988),
.Y(n_5462)
);

OAI21x1_ASAP7_75t_L g5463 ( 
.A1(n_5127),
.A2(n_4957),
.B(n_4940),
.Y(n_5463)
);

OAI21x1_ASAP7_75t_L g5464 ( 
.A1(n_5152),
.A2(n_4964),
.B(n_4753),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5069),
.Y(n_5465)
);

AND2x4_ASAP7_75t_L g5466 ( 
.A(n_5053),
.B(n_4642),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_5063),
.B(n_4989),
.Y(n_5467)
);

AOI221x1_ASAP7_75t_L g5468 ( 
.A1(n_5200),
.A2(n_4819),
.B1(n_4828),
.B2(n_5025),
.C(n_5020),
.Y(n_5468)
);

AOI21xp5_ASAP7_75t_L g5469 ( 
.A1(n_5082),
.A2(n_4878),
.B(n_4902),
.Y(n_5469)
);

NAND2xp5_ASAP7_75t_L g5470 ( 
.A(n_5395),
.B(n_4984),
.Y(n_5470)
);

OAI21xp5_ASAP7_75t_L g5471 ( 
.A1(n_5392),
.A2(n_4799),
.B(n_4795),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_5395),
.B(n_4995),
.Y(n_5472)
);

OAI21x1_ASAP7_75t_L g5473 ( 
.A1(n_5159),
.A2(n_5170),
.B(n_5171),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_5195),
.A2(n_4902),
.B(n_4868),
.Y(n_5474)
);

NOR4xp25_ASAP7_75t_L g5475 ( 
.A(n_5392),
.B(n_5001),
.C(n_4999),
.D(n_5027),
.Y(n_5475)
);

A2O1A1Ixp33_ASAP7_75t_L g5476 ( 
.A1(n_5226),
.A2(n_4811),
.B(n_4959),
.C(n_4673),
.Y(n_5476)
);

OAI21x1_ASAP7_75t_L g5477 ( 
.A1(n_5292),
.A2(n_4673),
.B(n_4642),
.Y(n_5477)
);

AOI21x1_ASAP7_75t_SL g5478 ( 
.A1(n_5229),
.A2(n_4899),
.B(n_4),
.Y(n_5478)
);

AND2x6_ASAP7_75t_L g5479 ( 
.A(n_5254),
.B(n_4719),
.Y(n_5479)
);

OAI21x1_ASAP7_75t_L g5480 ( 
.A1(n_5111),
.A2(n_4719),
.B(n_4962),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5080),
.Y(n_5481)
);

INVx1_ASAP7_75t_SL g5482 ( 
.A(n_5328),
.Y(n_5482)
);

OAI21xp5_ASAP7_75t_L g5483 ( 
.A1(n_5324),
.A2(n_1687),
.B(n_1673),
.Y(n_5483)
);

AO31x2_ASAP7_75t_L g5484 ( 
.A1(n_5234),
.A2(n_1694),
.A3(n_1696),
.B(n_1689),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5086),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5060),
.Y(n_5486)
);

OAI21xp5_ASAP7_75t_L g5487 ( 
.A1(n_5226),
.A2(n_1694),
.B(n_1689),
.Y(n_5487)
);

AOI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_5140),
.A2(n_5173),
.B(n_5161),
.Y(n_5488)
);

OAI21xp33_ASAP7_75t_L g5489 ( 
.A1(n_5062),
.A2(n_1700),
.B(n_1696),
.Y(n_5489)
);

INVx2_ASAP7_75t_L g5490 ( 
.A(n_5098),
.Y(n_5490)
);

OAI22xp5_ASAP7_75t_L g5491 ( 
.A1(n_5076),
.A2(n_1702),
.B1(n_1706),
.B2(n_1700),
.Y(n_5491)
);

OAI21x1_ASAP7_75t_L g5492 ( 
.A1(n_5262),
.A2(n_2944),
.B(n_2932),
.Y(n_5492)
);

AOI21xp5_ASAP7_75t_L g5493 ( 
.A1(n_5104),
.A2(n_2355),
.B(n_2321),
.Y(n_5493)
);

AOI21xp5_ASAP7_75t_L g5494 ( 
.A1(n_5085),
.A2(n_2355),
.B(n_2321),
.Y(n_5494)
);

AOI22xp5_ASAP7_75t_L g5495 ( 
.A1(n_5070),
.A2(n_758),
.B1(n_867),
.B2(n_748),
.Y(n_5495)
);

OAI22xp5_ASAP7_75t_L g5496 ( 
.A1(n_5449),
.A2(n_1706),
.B1(n_1709),
.B2(n_1702),
.Y(n_5496)
);

NOR2xp33_ASAP7_75t_L g5497 ( 
.A(n_5142),
.B(n_1708),
.Y(n_5497)
);

OAI21x1_ASAP7_75t_SL g5498 ( 
.A1(n_5091),
.A2(n_5413),
.B(n_5064),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_5182),
.B(n_1478),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_5342),
.B(n_1478),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5096),
.Y(n_5501)
);

NOR2xp33_ASAP7_75t_L g5502 ( 
.A(n_5167),
.B(n_1457),
.Y(n_5502)
);

OR2x2_ASAP7_75t_L g5503 ( 
.A(n_5277),
.B(n_1459),
.Y(n_5503)
);

NOR4xp25_ASAP7_75t_L g5504 ( 
.A(n_5059),
.B(n_5163),
.C(n_5209),
.D(n_5133),
.Y(n_5504)
);

BUFx3_ASAP7_75t_L g5505 ( 
.A(n_5122),
.Y(n_5505)
);

OAI21x1_ASAP7_75t_L g5506 ( 
.A1(n_5189),
.A2(n_2944),
.B(n_1710),
.Y(n_5506)
);

INVx2_ASAP7_75t_L g5507 ( 
.A(n_5156),
.Y(n_5507)
);

BUFx6f_ASAP7_75t_L g5508 ( 
.A(n_5128),
.Y(n_5508)
);

OAI21x1_ASAP7_75t_L g5509 ( 
.A1(n_5196),
.A2(n_2944),
.B(n_1710),
.Y(n_5509)
);

OR2x2_ASAP7_75t_L g5510 ( 
.A(n_5136),
.B(n_1459),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_5415),
.B(n_1540),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_L g5512 ( 
.A(n_5193),
.B(n_1540),
.Y(n_5512)
);

OAI21x1_ASAP7_75t_L g5513 ( 
.A1(n_5106),
.A2(n_2944),
.B(n_1709),
.Y(n_5513)
);

INVx3_ASAP7_75t_L g5514 ( 
.A(n_5093),
.Y(n_5514)
);

AOI21xp5_ASAP7_75t_L g5515 ( 
.A1(n_5215),
.A2(n_2355),
.B(n_2321),
.Y(n_5515)
);

OAI21x1_ASAP7_75t_L g5516 ( 
.A1(n_5083),
.A2(n_3054),
.B(n_3052),
.Y(n_5516)
);

AOI21xp5_ASAP7_75t_L g5517 ( 
.A1(n_5221),
.A2(n_2355),
.B(n_2321),
.Y(n_5517)
);

AOI22xp33_ASAP7_75t_L g5518 ( 
.A1(n_5219),
.A2(n_867),
.B1(n_957),
.B2(n_758),
.Y(n_5518)
);

AOI21xp5_ASAP7_75t_L g5519 ( 
.A1(n_5183),
.A2(n_2355),
.B(n_2321),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5157),
.Y(n_5520)
);

AND2x4_ASAP7_75t_L g5521 ( 
.A(n_5053),
.B(n_1613),
.Y(n_5521)
);

OAI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5217),
.A2(n_1464),
.B(n_1463),
.Y(n_5522)
);

AOI21xp5_ASAP7_75t_L g5523 ( 
.A1(n_5183),
.A2(n_2321),
.B(n_3359),
.Y(n_5523)
);

OAI21x1_ASAP7_75t_L g5524 ( 
.A1(n_5307),
.A2(n_3057),
.B(n_3054),
.Y(n_5524)
);

AO31x2_ASAP7_75t_L g5525 ( 
.A1(n_5434),
.A2(n_1625),
.A3(n_1630),
.B(n_1618),
.Y(n_5525)
);

OAI22x1_ASAP7_75t_L g5526 ( 
.A1(n_5079),
.A2(n_1625),
.B1(n_1630),
.B2(n_1618),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_L g5527 ( 
.A(n_5188),
.B(n_1463),
.Y(n_5527)
);

INVx2_ASAP7_75t_SL g5528 ( 
.A(n_5128),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5073),
.B(n_5100),
.Y(n_5529)
);

OAI21x1_ASAP7_75t_L g5530 ( 
.A1(n_5238),
.A2(n_3059),
.B(n_3057),
.Y(n_5530)
);

OAI21x1_ASAP7_75t_L g5531 ( 
.A1(n_5242),
.A2(n_3075),
.B(n_3059),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_5100),
.B(n_1464),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5299),
.B(n_1465),
.Y(n_5533)
);

OAI21xp5_ASAP7_75t_L g5534 ( 
.A1(n_5103),
.A2(n_1470),
.B(n_1465),
.Y(n_5534)
);

OAI21x1_ASAP7_75t_L g5535 ( 
.A1(n_5235),
.A2(n_3077),
.B(n_3075),
.Y(n_5535)
);

AO31x2_ASAP7_75t_L g5536 ( 
.A1(n_5075),
.A2(n_1636),
.A3(n_1638),
.B(n_1632),
.Y(n_5536)
);

NAND2xp5_ASAP7_75t_L g5537 ( 
.A(n_5074),
.B(n_5102),
.Y(n_5537)
);

NOR2xp33_ASAP7_75t_L g5538 ( 
.A(n_5105),
.B(n_1470),
.Y(n_5538)
);

AND2x4_ASAP7_75t_L g5539 ( 
.A(n_5430),
.B(n_1632),
.Y(n_5539)
);

AND2x2_ASAP7_75t_L g5540 ( 
.A(n_5160),
.B(n_1471),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_L g5541 ( 
.A(n_5102),
.B(n_5455),
.Y(n_5541)
);

AOI21xp5_ASAP7_75t_L g5542 ( 
.A1(n_5089),
.A2(n_2794),
.B(n_2946),
.Y(n_5542)
);

AOI21xp5_ASAP7_75t_L g5543 ( 
.A1(n_5089),
.A2(n_2955),
.B(n_2946),
.Y(n_5543)
);

OAI21xp5_ASAP7_75t_L g5544 ( 
.A1(n_5288),
.A2(n_1482),
.B(n_1471),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_5147),
.B(n_1482),
.Y(n_5545)
);

AOI22xp5_ASAP7_75t_L g5546 ( 
.A1(n_5081),
.A2(n_867),
.B1(n_957),
.B2(n_758),
.Y(n_5546)
);

O2A1O1Ixp33_ASAP7_75t_L g5547 ( 
.A1(n_5163),
.A2(n_1638),
.B(n_1639),
.C(n_1636),
.Y(n_5547)
);

BUFx2_ASAP7_75t_L g5548 ( 
.A(n_5408),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5110),
.Y(n_5549)
);

CKINVDCx5p33_ASAP7_75t_R g5550 ( 
.A(n_5061),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5151),
.B(n_1487),
.Y(n_5551)
);

AO21x2_ASAP7_75t_L g5552 ( 
.A1(n_5075),
.A2(n_1640),
.B(n_1639),
.Y(n_5552)
);

INVx6_ASAP7_75t_SL g5553 ( 
.A(n_5207),
.Y(n_5553)
);

OAI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5220),
.A2(n_1489),
.B(n_1487),
.Y(n_5554)
);

AO31x2_ASAP7_75t_L g5555 ( 
.A1(n_5454),
.A2(n_5174),
.A3(n_5078),
.B(n_5418),
.Y(n_5555)
);

INVx5_ASAP7_75t_L g5556 ( 
.A(n_5353),
.Y(n_5556)
);

OAI21x1_ASAP7_75t_SL g5557 ( 
.A1(n_5120),
.A2(n_1640),
.B(n_1491),
.Y(n_5557)
);

INVx5_ASAP7_75t_L g5558 ( 
.A(n_5353),
.Y(n_5558)
);

AOI22xp5_ASAP7_75t_L g5559 ( 
.A1(n_5112),
.A2(n_867),
.B1(n_957),
.B2(n_758),
.Y(n_5559)
);

AO21x1_ASAP7_75t_L g5560 ( 
.A1(n_5285),
.A2(n_1491),
.B(n_1489),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5118),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_5105),
.B(n_1495),
.Y(n_5562)
);

OAI21x1_ASAP7_75t_L g5563 ( 
.A1(n_5266),
.A2(n_3078),
.B(n_3077),
.Y(n_5563)
);

AOI211x1_ASAP7_75t_L g5564 ( 
.A1(n_5201),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_5564)
);

OAI21xp5_ASAP7_75t_L g5565 ( 
.A1(n_5267),
.A2(n_1496),
.B(n_1495),
.Y(n_5565)
);

OAI21x1_ASAP7_75t_L g5566 ( 
.A1(n_5279),
.A2(n_3083),
.B(n_3078),
.Y(n_5566)
);

NAND2xp5_ASAP7_75t_L g5567 ( 
.A(n_5056),
.B(n_1496),
.Y(n_5567)
);

AOI21xp5_ASAP7_75t_L g5568 ( 
.A1(n_5204),
.A2(n_2955),
.B(n_2906),
.Y(n_5568)
);

OAI21x1_ASAP7_75t_L g5569 ( 
.A1(n_5416),
.A2(n_3089),
.B(n_3083),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_5129),
.Y(n_5570)
);

AOI21xp5_ASAP7_75t_L g5571 ( 
.A1(n_5204),
.A2(n_2906),
.B(n_2904),
.Y(n_5571)
);

NAND3xp33_ASAP7_75t_L g5572 ( 
.A(n_5092),
.B(n_5243),
.C(n_5306),
.Y(n_5572)
);

AND2x4_ASAP7_75t_L g5573 ( 
.A(n_5435),
.B(n_1499),
.Y(n_5573)
);

OA21x2_ASAP7_75t_L g5574 ( 
.A1(n_5058),
.A2(n_1500),
.B(n_1499),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_5067),
.B(n_1500),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_SL g5576 ( 
.A(n_5218),
.B(n_1503),
.Y(n_5576)
);

AOI21xp5_ASAP7_75t_L g5577 ( 
.A1(n_5252),
.A2(n_2911),
.B(n_2904),
.Y(n_5577)
);

AOI221x1_ASAP7_75t_L g5578 ( 
.A1(n_5190),
.A2(n_1514),
.B1(n_1516),
.B2(n_1513),
.C(n_1503),
.Y(n_5578)
);

OAI22xp5_ASAP7_75t_L g5579 ( 
.A1(n_5109),
.A2(n_3101),
.B1(n_3111),
.B2(n_3089),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5385),
.B(n_1513),
.Y(n_5580)
);

INVx3_ASAP7_75t_L g5581 ( 
.A(n_5240),
.Y(n_5581)
);

AOI21xp5_ASAP7_75t_L g5582 ( 
.A1(n_5252),
.A2(n_2912),
.B(n_2911),
.Y(n_5582)
);

OAI22xp5_ASAP7_75t_L g5583 ( 
.A1(n_5109),
.A2(n_3111),
.B1(n_3114),
.B2(n_3101),
.Y(n_5583)
);

O2A1O1Ixp5_ASAP7_75t_L g5584 ( 
.A1(n_5139),
.A2(n_1516),
.B(n_1518),
.C(n_1514),
.Y(n_5584)
);

OAI22x1_ASAP7_75t_L g5585 ( 
.A1(n_5178),
.A2(n_5333),
.B1(n_5107),
.B2(n_5146),
.Y(n_5585)
);

OA21x2_ASAP7_75t_L g5586 ( 
.A1(n_5065),
.A2(n_1519),
.B(n_1518),
.Y(n_5586)
);

OAI22x1_ASAP7_75t_L g5587 ( 
.A1(n_5132),
.A2(n_1524),
.B1(n_1526),
.B2(n_1519),
.Y(n_5587)
);

A2O1A1Ixp33_ASAP7_75t_L g5588 ( 
.A1(n_5243),
.A2(n_1526),
.B(n_1528),
.C(n_1524),
.Y(n_5588)
);

OAI22xp5_ASAP7_75t_L g5589 ( 
.A1(n_5259),
.A2(n_3124),
.B1(n_3129),
.B2(n_3114),
.Y(n_5589)
);

OAI21x1_ASAP7_75t_L g5590 ( 
.A1(n_5419),
.A2(n_3129),
.B(n_3124),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5150),
.Y(n_5591)
);

INVx3_ASAP7_75t_L g5592 ( 
.A(n_5240),
.Y(n_5592)
);

BUFx3_ASAP7_75t_L g5593 ( 
.A(n_5222),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_5158),
.Y(n_5594)
);

AO21x1_ASAP7_75t_L g5595 ( 
.A1(n_5285),
.A2(n_1530),
.B(n_1528),
.Y(n_5595)
);

AND2x4_ASAP7_75t_L g5596 ( 
.A(n_5199),
.B(n_1530),
.Y(n_5596)
);

NOR2xp33_ASAP7_75t_L g5597 ( 
.A(n_5321),
.B(n_5359),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5177),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5304),
.Y(n_5599)
);

NAND3xp33_ASAP7_75t_L g5600 ( 
.A(n_5306),
.B(n_1532),
.C(n_1531),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5345),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_5263),
.Y(n_5602)
);

NAND3xp33_ASAP7_75t_L g5603 ( 
.A(n_5330),
.B(n_1532),
.C(n_1531),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5311),
.Y(n_5604)
);

OAI21x1_ASAP7_75t_L g5605 ( 
.A1(n_5426),
.A2(n_3134),
.B(n_3132),
.Y(n_5605)
);

AND2x2_ASAP7_75t_SL g5606 ( 
.A(n_5143),
.B(n_1541),
.Y(n_5606)
);

OAI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_5259),
.A2(n_3134),
.B1(n_3143),
.B2(n_3132),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_L g5608 ( 
.A(n_5385),
.B(n_1541),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_5125),
.B(n_1544),
.Y(n_5609)
);

BUFx2_ASAP7_75t_L g5610 ( 
.A(n_5199),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5331),
.Y(n_5611)
);

OAI22xp5_ASAP7_75t_L g5612 ( 
.A1(n_5135),
.A2(n_3153),
.B1(n_3154),
.B2(n_3143),
.Y(n_5612)
);

OAI21x1_ASAP7_75t_L g5613 ( 
.A1(n_5427),
.A2(n_5432),
.B(n_5296),
.Y(n_5613)
);

BUFx10_ASAP7_75t_L g5614 ( 
.A(n_5406),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5338),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_SL g5616 ( 
.A(n_5414),
.B(n_5054),
.Y(n_5616)
);

AOI21xp5_ASAP7_75t_L g5617 ( 
.A1(n_5101),
.A2(n_2922),
.B(n_2912),
.Y(n_5617)
);

OAI21x1_ASAP7_75t_L g5618 ( 
.A1(n_5313),
.A2(n_3154),
.B(n_3153),
.Y(n_5618)
);

INVx1_ASAP7_75t_SL g5619 ( 
.A(n_5077),
.Y(n_5619)
);

NAND3xp33_ASAP7_75t_L g5620 ( 
.A(n_5330),
.B(n_1546),
.C(n_1544),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_5302),
.A2(n_2923),
.B(n_2922),
.Y(n_5621)
);

A2O1A1Ixp33_ASAP7_75t_L g5622 ( 
.A1(n_5443),
.A2(n_1549),
.B(n_1550),
.C(n_1546),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5346),
.Y(n_5623)
);

AOI221x1_ASAP7_75t_L g5624 ( 
.A1(n_5402),
.A2(n_1552),
.B1(n_1555),
.B2(n_1550),
.C(n_1549),
.Y(n_5624)
);

OA21x2_ASAP7_75t_L g5625 ( 
.A1(n_5068),
.A2(n_1555),
.B(n_1552),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5134),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5212),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5214),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5233),
.Y(n_5629)
);

AND2x2_ASAP7_75t_L g5630 ( 
.A(n_5210),
.B(n_1557),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5247),
.Y(n_5631)
);

NAND3xp33_ASAP7_75t_L g5632 ( 
.A(n_5343),
.B(n_1560),
.C(n_1557),
.Y(n_5632)
);

BUFx3_ASAP7_75t_L g5633 ( 
.A(n_5375),
.Y(n_5633)
);

NAND2xp5_ASAP7_75t_L g5634 ( 
.A(n_5185),
.B(n_1560),
.Y(n_5634)
);

NAND2xp5_ASAP7_75t_L g5635 ( 
.A(n_5229),
.B(n_1562),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5369),
.Y(n_5636)
);

BUFx10_ASAP7_75t_L g5637 ( 
.A(n_5258),
.Y(n_5637)
);

OAI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5230),
.A2(n_3163),
.B1(n_3164),
.B2(n_3161),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_5237),
.B(n_1562),
.Y(n_5639)
);

AO21x1_ASAP7_75t_L g5640 ( 
.A1(n_5291),
.A2(n_1575),
.B(n_1570),
.Y(n_5640)
);

INVxp67_ASAP7_75t_SL g5641 ( 
.A(n_5187),
.Y(n_5641)
);

NOR2xp33_ASAP7_75t_L g5642 ( 
.A(n_5224),
.B(n_1570),
.Y(n_5642)
);

OAI21x1_ASAP7_75t_L g5643 ( 
.A1(n_5445),
.A2(n_3163),
.B(n_3161),
.Y(n_5643)
);

OAI21x1_ASAP7_75t_L g5644 ( 
.A1(n_5456),
.A2(n_3167),
.B(n_3164),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_5237),
.B(n_1575),
.Y(n_5645)
);

AOI21xp5_ASAP7_75t_L g5646 ( 
.A1(n_5302),
.A2(n_2926),
.B(n_2923),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5077),
.Y(n_5647)
);

BUFx10_ASAP7_75t_L g5648 ( 
.A(n_5055),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5249),
.B(n_1576),
.Y(n_5649)
);

INVx2_ASAP7_75t_L g5650 ( 
.A(n_5438),
.Y(n_5650)
);

OAI21x1_ASAP7_75t_L g5651 ( 
.A1(n_5457),
.A2(n_3167),
.B(n_1578),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5138),
.Y(n_5652)
);

AO31x2_ASAP7_75t_L g5653 ( 
.A1(n_5197),
.A2(n_1578),
.A3(n_1576),
.B(n_2593),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_5340),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5340),
.Y(n_5655)
);

AOI21xp33_ASAP7_75t_L g5656 ( 
.A1(n_5205),
.A2(n_2359),
.B(n_2357),
.Y(n_5656)
);

OAI21x1_ASAP7_75t_L g5657 ( 
.A1(n_5269),
.A2(n_2527),
.B(n_2597),
.Y(n_5657)
);

OAI21x1_ASAP7_75t_SL g5658 ( 
.A1(n_5310),
.A2(n_3),
.B(n_4),
.Y(n_5658)
);

OAI21x1_ASAP7_75t_L g5659 ( 
.A1(n_5270),
.A2(n_2527),
.B(n_2597),
.Y(n_5659)
);

NOR2xp33_ASAP7_75t_L g5660 ( 
.A(n_5227),
.B(n_57),
.Y(n_5660)
);

OAI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_5343),
.A2(n_2363),
.B(n_2362),
.Y(n_5661)
);

NAND2xp33_ASAP7_75t_L g5662 ( 
.A(n_5414),
.B(n_3291),
.Y(n_5662)
);

NAND2xp5_ASAP7_75t_L g5663 ( 
.A(n_5249),
.B(n_57),
.Y(n_5663)
);

OAI21x1_ASAP7_75t_L g5664 ( 
.A1(n_5121),
.A2(n_2527),
.B(n_2551),
.Y(n_5664)
);

AND2x4_ASAP7_75t_L g5665 ( 
.A(n_5199),
.B(n_58),
.Y(n_5665)
);

OAI21x1_ASAP7_75t_L g5666 ( 
.A1(n_5248),
.A2(n_2551),
.B(n_2926),
.Y(n_5666)
);

AOI21xp5_ASAP7_75t_L g5667 ( 
.A1(n_5099),
.A2(n_2950),
.B(n_2938),
.Y(n_5667)
);

AOI221x1_ASAP7_75t_L g5668 ( 
.A1(n_5291),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_5668)
);

NAND2x1p5_ASAP7_75t_L g5669 ( 
.A(n_5099),
.B(n_3136),
.Y(n_5669)
);

INVxp67_ASAP7_75t_L g5670 ( 
.A(n_5373),
.Y(n_5670)
);

AND2x4_ASAP7_75t_L g5671 ( 
.A(n_5099),
.B(n_58),
.Y(n_5671)
);

AND2x2_ASAP7_75t_L g5672 ( 
.A(n_5303),
.B(n_957),
.Y(n_5672)
);

OAI21xp5_ASAP7_75t_L g5673 ( 
.A1(n_5198),
.A2(n_2363),
.B(n_2362),
.Y(n_5673)
);

BUFx2_ASAP7_75t_R g5674 ( 
.A(n_5393),
.Y(n_5674)
);

AOI21xp5_ASAP7_75t_L g5675 ( 
.A1(n_5099),
.A2(n_2950),
.B(n_2938),
.Y(n_5675)
);

BUFx6f_ASAP7_75t_L g5676 ( 
.A(n_5128),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5282),
.Y(n_5677)
);

AOI21xp5_ASAP7_75t_L g5678 ( 
.A1(n_5194),
.A2(n_2961),
.B(n_2951),
.Y(n_5678)
);

AOI21xp5_ASAP7_75t_L g5679 ( 
.A1(n_5194),
.A2(n_5087),
.B(n_5293),
.Y(n_5679)
);

AOI22xp5_ASAP7_75t_L g5680 ( 
.A1(n_5323),
.A2(n_1221),
.B1(n_1239),
.B2(n_990),
.Y(n_5680)
);

AOI21xp5_ASAP7_75t_SL g5681 ( 
.A1(n_5295),
.A2(n_3166),
.B(n_3136),
.Y(n_5681)
);

AOI21x1_ASAP7_75t_L g5682 ( 
.A1(n_5084),
.A2(n_2407),
.B(n_2406),
.Y(n_5682)
);

O2A1O1Ixp33_ASAP7_75t_SL g5683 ( 
.A1(n_5145),
.A2(n_60),
.B(n_62),
.C(n_59),
.Y(n_5683)
);

NAND2xp5_ASAP7_75t_L g5684 ( 
.A(n_5264),
.B(n_59),
.Y(n_5684)
);

OAI21x1_ASAP7_75t_L g5685 ( 
.A1(n_5253),
.A2(n_2551),
.B(n_2951),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_5264),
.B(n_60),
.Y(n_5686)
);

AO31x2_ASAP7_75t_L g5687 ( 
.A1(n_5203),
.A2(n_5211),
.A3(n_5399),
.B(n_5294),
.Y(n_5687)
);

NAND2xp5_ASAP7_75t_L g5688 ( 
.A(n_5268),
.B(n_62),
.Y(n_5688)
);

AOI21xp5_ASAP7_75t_L g5689 ( 
.A1(n_5194),
.A2(n_2963),
.B(n_2961),
.Y(n_5689)
);

AOI21x1_ASAP7_75t_L g5690 ( 
.A1(n_5268),
.A2(n_2407),
.B(n_2406),
.Y(n_5690)
);

OAI21x1_ASAP7_75t_L g5691 ( 
.A1(n_5255),
.A2(n_2964),
.B(n_2963),
.Y(n_5691)
);

AOI21xp5_ASAP7_75t_L g5692 ( 
.A1(n_5194),
.A2(n_2967),
.B(n_2964),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5282),
.Y(n_5693)
);

OAI21x1_ASAP7_75t_L g5694 ( 
.A1(n_5094),
.A2(n_2972),
.B(n_2967),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5280),
.B(n_63),
.Y(n_5695)
);

O2A1O1Ixp33_ASAP7_75t_L g5696 ( 
.A1(n_5168),
.A2(n_5317),
.B(n_5300),
.C(n_5232),
.Y(n_5696)
);

INVx3_ASAP7_75t_L g5697 ( 
.A(n_5439),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_5280),
.B(n_63),
.Y(n_5698)
);

BUFx2_ASAP7_75t_L g5699 ( 
.A(n_5066),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5154),
.B(n_990),
.Y(n_5700)
);

AOI22xp5_ASAP7_75t_L g5701 ( 
.A1(n_5323),
.A2(n_1221),
.B1(n_1239),
.B2(n_990),
.Y(n_5701)
);

CKINVDCx5p33_ASAP7_75t_R g5702 ( 
.A(n_5057),
.Y(n_5702)
);

O2A1O1Ixp5_ASAP7_75t_L g5703 ( 
.A1(n_5213),
.A2(n_1221),
.B(n_1239),
.C(n_990),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5282),
.Y(n_5704)
);

BUFx4_ASAP7_75t_SL g5705 ( 
.A(n_5377),
.Y(n_5705)
);

AOI21xp5_ASAP7_75t_L g5706 ( 
.A1(n_5293),
.A2(n_5273),
.B(n_5208),
.Y(n_5706)
);

OR2x2_ASAP7_75t_L g5707 ( 
.A(n_5186),
.B(n_64),
.Y(n_5707)
);

NOR2xp67_ASAP7_75t_L g5708 ( 
.A(n_5294),
.B(n_5),
.Y(n_5708)
);

OAI21x1_ASAP7_75t_L g5709 ( 
.A1(n_5153),
.A2(n_5422),
.B(n_5365),
.Y(n_5709)
);

NAND2xp5_ASAP7_75t_L g5710 ( 
.A(n_5281),
.B(n_65),
.Y(n_5710)
);

AOI21xp5_ASAP7_75t_L g5711 ( 
.A1(n_5273),
.A2(n_2976),
.B(n_2974),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5287),
.Y(n_5712)
);

OAI21x1_ASAP7_75t_L g5713 ( 
.A1(n_5356),
.A2(n_5374),
.B(n_5090),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5287),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5281),
.B(n_65),
.Y(n_5715)
);

AO31x2_ASAP7_75t_L g5716 ( 
.A1(n_5289),
.A2(n_2402),
.A3(n_2377),
.B(n_2379),
.Y(n_5716)
);

OAI21xp33_ASAP7_75t_L g5717 ( 
.A1(n_5230),
.A2(n_1239),
.B(n_1221),
.Y(n_5717)
);

NAND3xp33_ASAP7_75t_L g5718 ( 
.A(n_5341),
.B(n_2978),
.C(n_2977),
.Y(n_5718)
);

O2A1O1Ixp5_ASAP7_75t_SL g5719 ( 
.A1(n_5410),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_5719)
);

BUFx6f_ASAP7_75t_L g5720 ( 
.A(n_5378),
.Y(n_5720)
);

AOI22xp5_ASAP7_75t_L g5721 ( 
.A1(n_5130),
.A2(n_3291),
.B1(n_2978),
.B2(n_2977),
.Y(n_5721)
);

CKINVDCx5p33_ASAP7_75t_R g5722 ( 
.A(n_5115),
.Y(n_5722)
);

OAI21x1_ASAP7_75t_L g5723 ( 
.A1(n_5088),
.A2(n_2577),
.B(n_2703),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_5155),
.Y(n_5724)
);

O2A1O1Ixp33_ASAP7_75t_L g5725 ( 
.A1(n_5232),
.A2(n_9),
.B(n_6),
.C(n_8),
.Y(n_5725)
);

XOR2xp5_ASAP7_75t_L g5726 ( 
.A(n_5275),
.B(n_5126),
.Y(n_5726)
);

OAI21x1_ASAP7_75t_L g5727 ( 
.A1(n_5276),
.A2(n_2577),
.B(n_2703),
.Y(n_5727)
);

AOI21xp5_ASAP7_75t_L g5728 ( 
.A1(n_5208),
.A2(n_5298),
.B(n_5403),
.Y(n_5728)
);

NOR2xp67_ASAP7_75t_L g5729 ( 
.A(n_5314),
.B(n_10),
.Y(n_5729)
);

AOI21xp5_ASAP7_75t_L g5730 ( 
.A1(n_5403),
.A2(n_2717),
.B(n_2706),
.Y(n_5730)
);

AO22x1_ASAP7_75t_L g5731 ( 
.A1(n_5309),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_5731)
);

AOI21xp5_ASAP7_75t_L g5732 ( 
.A1(n_5246),
.A2(n_2717),
.B(n_2706),
.Y(n_5732)
);

AOI21xp33_ASAP7_75t_L g5733 ( 
.A1(n_5443),
.A2(n_12),
.B(n_11),
.Y(n_5733)
);

OAI21xp5_ASAP7_75t_L g5734 ( 
.A1(n_5271),
.A2(n_3291),
.B(n_2402),
.Y(n_5734)
);

A2O1A1Ixp33_ASAP7_75t_L g5735 ( 
.A1(n_5341),
.A2(n_68),
.B(n_70),
.C(n_66),
.Y(n_5735)
);

INVx2_ASAP7_75t_L g5736 ( 
.A(n_5066),
.Y(n_5736)
);

BUFx2_ASAP7_75t_L g5737 ( 
.A(n_5066),
.Y(n_5737)
);

A2O1A1Ixp33_ASAP7_75t_L g5738 ( 
.A1(n_5388),
.A2(n_68),
.B(n_70),
.C(n_66),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5287),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5066),
.Y(n_5740)
);

AO21x2_ASAP7_75t_L g5741 ( 
.A1(n_5347),
.A2(n_2377),
.B(n_2373),
.Y(n_5741)
);

AOI21xp5_ASAP7_75t_L g5742 ( 
.A1(n_5216),
.A2(n_2722),
.B(n_2667),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5072),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_5191),
.B(n_71),
.Y(n_5744)
);

OAI21xp33_ASAP7_75t_L g5745 ( 
.A1(n_5201),
.A2(n_10),
.B(n_11),
.Y(n_5745)
);

BUFx3_ASAP7_75t_L g5746 ( 
.A(n_5348),
.Y(n_5746)
);

NAND2xp5_ASAP7_75t_L g5747 ( 
.A(n_5206),
.B(n_71),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5066),
.Y(n_5748)
);

BUFx3_ASAP7_75t_L g5749 ( 
.A(n_5137),
.Y(n_5749)
);

NOR2xp67_ASAP7_75t_L g5750 ( 
.A(n_5314),
.B(n_13),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5357),
.Y(n_5751)
);

AOI211x1_ASAP7_75t_L g5752 ( 
.A1(n_5054),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_5752)
);

OAI21xp5_ASAP7_75t_L g5753 ( 
.A1(n_5272),
.A2(n_2379),
.B(n_2373),
.Y(n_5753)
);

NAND2xp5_ASAP7_75t_L g5754 ( 
.A(n_5410),
.B(n_72),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5389),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5379),
.Y(n_5756)
);

AOI221xp5_ASAP7_75t_SL g5757 ( 
.A1(n_5272),
.A2(n_30),
.B1(n_39),
.B2(n_21),
.C(n_13),
.Y(n_5757)
);

OAI21xp5_ASAP7_75t_L g5758 ( 
.A1(n_5325),
.A2(n_2387),
.B(n_2382),
.Y(n_5758)
);

O2A1O1Ixp5_ASAP7_75t_SL g5759 ( 
.A1(n_5332),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_5759)
);

OAI21x1_ASAP7_75t_L g5760 ( 
.A1(n_5223),
.A2(n_2577),
.B(n_2722),
.Y(n_5760)
);

OA21x2_ASAP7_75t_L g5761 ( 
.A1(n_5114),
.A2(n_2387),
.B(n_2382),
.Y(n_5761)
);

AOI221x1_ASAP7_75t_L g5762 ( 
.A1(n_5144),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.C(n_19),
.Y(n_5762)
);

OAI21x1_ASAP7_75t_L g5763 ( 
.A1(n_5108),
.A2(n_2395),
.B(n_2388),
.Y(n_5763)
);

NAND3x1_ASAP7_75t_L g5764 ( 
.A(n_5372),
.B(n_16),
.C(n_17),
.Y(n_5764)
);

OAI21x1_ASAP7_75t_L g5765 ( 
.A1(n_5124),
.A2(n_2395),
.B(n_2388),
.Y(n_5765)
);

AOI21xp5_ASAP7_75t_L g5766 ( 
.A1(n_5228),
.A2(n_2667),
.B(n_2658),
.Y(n_5766)
);

AOI21xp33_ASAP7_75t_L g5767 ( 
.A1(n_5409),
.A2(n_5417),
.B(n_5411),
.Y(n_5767)
);

AOI21x1_ASAP7_75t_L g5768 ( 
.A1(n_5350),
.A2(n_17),
.B(n_18),
.Y(n_5768)
);

NOR2xp67_ASAP7_75t_L g5769 ( 
.A(n_5316),
.B(n_19),
.Y(n_5769)
);

AOI21xp5_ASAP7_75t_L g5770 ( 
.A1(n_5228),
.A2(n_2667),
.B(n_2658),
.Y(n_5770)
);

NAND2xp5_ASAP7_75t_SL g5771 ( 
.A(n_5114),
.B(n_2286),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5316),
.B(n_72),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5382),
.Y(n_5773)
);

AOI21xp5_ASAP7_75t_L g5774 ( 
.A1(n_5428),
.A2(n_2667),
.B(n_3136),
.Y(n_5774)
);

OAI21x1_ASAP7_75t_L g5775 ( 
.A1(n_5180),
.A2(n_2405),
.B(n_2378),
.Y(n_5775)
);

AO31x2_ASAP7_75t_L g5776 ( 
.A1(n_5380),
.A2(n_22),
.A3(n_20),
.B(n_21),
.Y(n_5776)
);

AOI21x1_ASAP7_75t_L g5777 ( 
.A1(n_5380),
.A2(n_20),
.B(n_23),
.Y(n_5777)
);

OAI21xp5_ASAP7_75t_L g5778 ( 
.A1(n_5325),
.A2(n_2343),
.B(n_2329),
.Y(n_5778)
);

NAND3xp33_ASAP7_75t_SL g5779 ( 
.A(n_5352),
.B(n_5301),
.C(n_5256),
.Y(n_5779)
);

AO31x2_ASAP7_75t_L g5780 ( 
.A1(n_5383),
.A2(n_26),
.A3(n_23),
.B(n_24),
.Y(n_5780)
);

OAI21x1_ASAP7_75t_L g5781 ( 
.A1(n_5166),
.A2(n_2405),
.B(n_2378),
.Y(n_5781)
);

OAI21xp5_ASAP7_75t_L g5782 ( 
.A1(n_5358),
.A2(n_2343),
.B(n_2329),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5305),
.Y(n_5783)
);

AOI31xp67_ASAP7_75t_L g5784 ( 
.A1(n_5370),
.A2(n_27),
.A3(n_23),
.B(n_26),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5305),
.Y(n_5785)
);

NAND2xp5_ASAP7_75t_L g5786 ( 
.A(n_5383),
.B(n_73),
.Y(n_5786)
);

OAI21x1_ASAP7_75t_L g5787 ( 
.A1(n_5284),
.A2(n_2405),
.B(n_2378),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5071),
.B(n_75),
.Y(n_5788)
);

OAI21xp5_ASAP7_75t_L g5789 ( 
.A1(n_5308),
.A2(n_2343),
.B(n_2329),
.Y(n_5789)
);

AO32x2_ASAP7_75t_L g5790 ( 
.A1(n_5181),
.A2(n_28),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_5790)
);

NOR2xp33_ASAP7_75t_L g5791 ( 
.A(n_5141),
.B(n_76),
.Y(n_5791)
);

INVx3_ASAP7_75t_L g5792 ( 
.A(n_5439),
.Y(n_5792)
);

A2O1A1Ixp33_ASAP7_75t_L g5793 ( 
.A1(n_5398),
.A2(n_77),
.B(n_79),
.C(n_76),
.Y(n_5793)
);

OAI21x1_ASAP7_75t_SL g5794 ( 
.A1(n_5119),
.A2(n_28),
.B(n_29),
.Y(n_5794)
);

NAND2xp5_ASAP7_75t_L g5795 ( 
.A(n_5391),
.B(n_77),
.Y(n_5795)
);

AOI221x1_ASAP7_75t_L g5796 ( 
.A1(n_5376),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.C(n_32),
.Y(n_5796)
);

AOI221x1_ASAP7_75t_L g5797 ( 
.A1(n_5391),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.C(n_35),
.Y(n_5797)
);

NAND2xp5_ASAP7_75t_SL g5798 ( 
.A(n_5119),
.B(n_5458),
.Y(n_5798)
);

OAI21x1_ASAP7_75t_L g5799 ( 
.A1(n_5172),
.A2(n_5176),
.B(n_5162),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5439),
.Y(n_5800)
);

AND2x4_ASAP7_75t_L g5801 ( 
.A(n_5207),
.B(n_80),
.Y(n_5801)
);

NAND2xp5_ASAP7_75t_L g5802 ( 
.A(n_5396),
.B(n_81),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5305),
.Y(n_5803)
);

OAI21x1_ASAP7_75t_L g5804 ( 
.A1(n_5131),
.A2(n_2405),
.B(n_2378),
.Y(n_5804)
);

NAND2xp5_ASAP7_75t_L g5805 ( 
.A(n_5396),
.B(n_81),
.Y(n_5805)
);

OAI21x1_ASAP7_75t_L g5806 ( 
.A1(n_5148),
.A2(n_2200),
.B(n_2195),
.Y(n_5806)
);

AO21x2_ASAP7_75t_L g5807 ( 
.A1(n_5498),
.A2(n_5401),
.B(n_5169),
.Y(n_5807)
);

OAI22x1_ASAP7_75t_L g5808 ( 
.A1(n_5619),
.A2(n_5095),
.B1(n_5175),
.B2(n_5371),
.Y(n_5808)
);

AO21x2_ASAP7_75t_L g5809 ( 
.A1(n_5475),
.A2(n_5401),
.B(n_5169),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5548),
.Y(n_5810)
);

INVx5_ASAP7_75t_L g5811 ( 
.A(n_5720),
.Y(n_5811)
);

BUFx2_ASAP7_75t_R g5812 ( 
.A(n_5724),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5594),
.Y(n_5813)
);

OR2x6_ASAP7_75t_L g5814 ( 
.A(n_5679),
.B(n_5257),
.Y(n_5814)
);

BUFx2_ASAP7_75t_L g5815 ( 
.A(n_5553),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5465),
.Y(n_5816)
);

OAI21x1_ASAP7_75t_L g5817 ( 
.A1(n_5488),
.A2(n_5424),
.B(n_5164),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5481),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_5705),
.Y(n_5819)
);

BUFx2_ASAP7_75t_L g5820 ( 
.A(n_5553),
.Y(n_5820)
);

OAI21x1_ASAP7_75t_L g5821 ( 
.A1(n_5713),
.A2(n_5239),
.B(n_5327),
.Y(n_5821)
);

INVx4_ASAP7_75t_L g5822 ( 
.A(n_5720),
.Y(n_5822)
);

INVx3_ASAP7_75t_L g5823 ( 
.A(n_5514),
.Y(n_5823)
);

INVx8_ASAP7_75t_L g5824 ( 
.A(n_5720),
.Y(n_5824)
);

OAI21xp5_ASAP7_75t_L g5825 ( 
.A1(n_5475),
.A2(n_5468),
.B(n_5616),
.Y(n_5825)
);

INVxp67_ASAP7_75t_SL g5826 ( 
.A(n_5503),
.Y(n_5826)
);

BUFx2_ASAP7_75t_L g5827 ( 
.A(n_5610),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5485),
.Y(n_5828)
);

OAI21x1_ASAP7_75t_L g5829 ( 
.A1(n_5477),
.A2(n_5239),
.B(n_5329),
.Y(n_5829)
);

BUFx2_ASAP7_75t_L g5830 ( 
.A(n_5466),
.Y(n_5830)
);

AND2x4_ASAP7_75t_L g5831 ( 
.A(n_5514),
.B(n_5420),
.Y(n_5831)
);

BUFx3_ASAP7_75t_L g5832 ( 
.A(n_5746),
.Y(n_5832)
);

OAI21x1_ASAP7_75t_SL g5833 ( 
.A1(n_5794),
.A2(n_5433),
.B(n_5332),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5501),
.Y(n_5834)
);

AOI22xp33_ASAP7_75t_L g5835 ( 
.A1(n_5572),
.A2(n_5245),
.B1(n_5334),
.B2(n_5398),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5549),
.Y(n_5836)
);

AO21x2_ASAP7_75t_L g5837 ( 
.A1(n_5677),
.A2(n_5429),
.B(n_5425),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5561),
.Y(n_5838)
);

OAI21x1_ASAP7_75t_L g5839 ( 
.A1(n_5494),
.A2(n_5339),
.B(n_5335),
.Y(n_5839)
);

INVx1_ASAP7_75t_L g5840 ( 
.A(n_5570),
.Y(n_5840)
);

INVxp67_ASAP7_75t_L g5841 ( 
.A(n_5533),
.Y(n_5841)
);

AND2x4_ASAP7_75t_L g5842 ( 
.A(n_5647),
.B(n_5278),
.Y(n_5842)
);

AOI22x1_ASAP7_75t_L g5843 ( 
.A1(n_5471),
.A2(n_5453),
.B1(n_5244),
.B2(n_5254),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5591),
.Y(n_5844)
);

OAI21x1_ASAP7_75t_L g5845 ( 
.A1(n_5723),
.A2(n_5354),
.B(n_5344),
.Y(n_5845)
);

BUFx3_ASAP7_75t_L g5846 ( 
.A(n_5633),
.Y(n_5846)
);

NAND2xp5_ASAP7_75t_L g5847 ( 
.A(n_5743),
.B(n_5351),
.Y(n_5847)
);

AOI21xp5_ASAP7_75t_L g5848 ( 
.A1(n_5519),
.A2(n_5428),
.B(n_5431),
.Y(n_5848)
);

NAND2x1p5_ASAP7_75t_L g5849 ( 
.A(n_5556),
.B(n_5386),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5598),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5601),
.Y(n_5851)
);

OA21x2_ASAP7_75t_L g5852 ( 
.A1(n_5798),
.A2(n_5400),
.B(n_5394),
.Y(n_5852)
);

HB1xp67_ASAP7_75t_L g5853 ( 
.A(n_5627),
.Y(n_5853)
);

INVxp67_ASAP7_75t_SL g5854 ( 
.A(n_5783),
.Y(n_5854)
);

AND2x4_ASAP7_75t_L g5855 ( 
.A(n_5619),
.B(n_5736),
.Y(n_5855)
);

OAI21xp5_ASAP7_75t_L g5856 ( 
.A1(n_5680),
.A2(n_5431),
.B(n_5251),
.Y(n_5856)
);

AND2x2_ASAP7_75t_L g5857 ( 
.A(n_5641),
.B(n_5482),
.Y(n_5857)
);

AND2x4_ASAP7_75t_L g5858 ( 
.A(n_5740),
.B(n_5312),
.Y(n_5858)
);

OAI21xp5_ASAP7_75t_L g5859 ( 
.A1(n_5680),
.A2(n_5251),
.B(n_5336),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5628),
.Y(n_5860)
);

BUFx3_ASAP7_75t_L g5861 ( 
.A(n_5505),
.Y(n_5861)
);

OR2x6_ASAP7_75t_L g5862 ( 
.A(n_5469),
.B(n_5257),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5629),
.Y(n_5863)
);

BUFx8_ASAP7_75t_L g5864 ( 
.A(n_5630),
.Y(n_5864)
);

OA21x2_ASAP7_75t_L g5865 ( 
.A1(n_5748),
.A2(n_5097),
.B(n_5349),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5599),
.Y(n_5866)
);

AO31x2_ASAP7_75t_L g5867 ( 
.A1(n_5693),
.A2(n_5453),
.A3(n_5315),
.B(n_5274),
.Y(n_5867)
);

HB1xp67_ASAP7_75t_L g5868 ( 
.A(n_5631),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5486),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5490),
.Y(n_5870)
);

INVx2_ASAP7_75t_SL g5871 ( 
.A(n_5749),
.Y(n_5871)
);

AND2x4_ASAP7_75t_L g5872 ( 
.A(n_5482),
.B(n_5274),
.Y(n_5872)
);

INVx3_ASAP7_75t_L g5873 ( 
.A(n_5581),
.Y(n_5873)
);

NAND2xp5_ASAP7_75t_L g5874 ( 
.A(n_5636),
.B(n_5351),
.Y(n_5874)
);

OAI21x1_ASAP7_75t_L g5875 ( 
.A1(n_5709),
.A2(n_5192),
.B(n_5261),
.Y(n_5875)
);

OAI21x1_ASAP7_75t_L g5876 ( 
.A1(n_5799),
.A2(n_5261),
.B(n_5386),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5652),
.B(n_5265),
.Y(n_5877)
);

OR2x2_ASAP7_75t_L g5878 ( 
.A(n_5529),
.B(n_5351),
.Y(n_5878)
);

OA21x2_ASAP7_75t_L g5879 ( 
.A1(n_5704),
.A2(n_5326),
.B(n_5117),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5626),
.B(n_5537),
.Y(n_5880)
);

OAI21x1_ASAP7_75t_L g5881 ( 
.A1(n_5613),
.A2(n_5322),
.B(n_5384),
.Y(n_5881)
);

OAI21x1_ASAP7_75t_L g5882 ( 
.A1(n_5694),
.A2(n_5397),
.B(n_5225),
.Y(n_5882)
);

OAI21x1_ASAP7_75t_L g5883 ( 
.A1(n_5682),
.A2(n_5236),
.B(n_5283),
.Y(n_5883)
);

OAI21x1_ASAP7_75t_SL g5884 ( 
.A1(n_5754),
.A2(n_5451),
.B(n_5116),
.Y(n_5884)
);

NOR2xp67_ASAP7_75t_SL g5885 ( 
.A(n_5459),
.B(n_5265),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5541),
.B(n_5361),
.Y(n_5886)
);

INVx6_ASAP7_75t_L g5887 ( 
.A(n_5614),
.Y(n_5887)
);

OAI21xp5_ASAP7_75t_L g5888 ( 
.A1(n_5701),
.A2(n_5451),
.B(n_5179),
.Y(n_5888)
);

OAI21x1_ASAP7_75t_L g5889 ( 
.A1(n_5543),
.A2(n_5286),
.B(n_5440),
.Y(n_5889)
);

OAI21x1_ASAP7_75t_L g5890 ( 
.A1(n_5473),
.A2(n_5318),
.B(n_5319),
.Y(n_5890)
);

OAI21x1_ASAP7_75t_L g5891 ( 
.A1(n_5785),
.A2(n_5116),
.B(n_5405),
.Y(n_5891)
);

OAI21x1_ASAP7_75t_L g5892 ( 
.A1(n_5803),
.A2(n_5441),
.B(n_5412),
.Y(n_5892)
);

INVx1_ASAP7_75t_SL g5893 ( 
.A(n_5699),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5650),
.Y(n_5894)
);

OAI21x1_ASAP7_75t_L g5895 ( 
.A1(n_5712),
.A2(n_5404),
.B(n_5297),
.Y(n_5895)
);

OAI21x1_ASAP7_75t_SL g5896 ( 
.A1(n_5658),
.A2(n_5315),
.B(n_5355),
.Y(n_5896)
);

OAI21x1_ASAP7_75t_L g5897 ( 
.A1(n_5714),
.A2(n_5446),
.B(n_5442),
.Y(n_5897)
);

INVx2_ASAP7_75t_L g5898 ( 
.A(n_5654),
.Y(n_5898)
);

INVx2_ASAP7_75t_SL g5899 ( 
.A(n_5593),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5602),
.B(n_5361),
.Y(n_5900)
);

OAI21xp5_ASAP7_75t_L g5901 ( 
.A1(n_5701),
.A2(n_5179),
.B(n_5452),
.Y(n_5901)
);

NOR2xp67_ASAP7_75t_L g5902 ( 
.A(n_5585),
.B(n_5360),
.Y(n_5902)
);

OAI21x1_ASAP7_75t_L g5903 ( 
.A1(n_5739),
.A2(n_5450),
.B(n_5447),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5507),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5737),
.B(n_5361),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5520),
.Y(n_5906)
);

OAI21x1_ASAP7_75t_L g5907 ( 
.A1(n_5763),
.A2(n_5387),
.B(n_5381),
.Y(n_5907)
);

OAI21x1_ASAP7_75t_SL g5908 ( 
.A1(n_5459),
.A2(n_5368),
.B(n_5366),
.Y(n_5908)
);

INVx3_ASAP7_75t_L g5909 ( 
.A(n_5581),
.Y(n_5909)
);

AOI21xp5_ASAP7_75t_L g5910 ( 
.A1(n_5774),
.A2(n_5245),
.B(n_5117),
.Y(n_5910)
);

OAI21x1_ASAP7_75t_L g5911 ( 
.A1(n_5506),
.A2(n_5448),
.B(n_5444),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_5655),
.Y(n_5912)
);

INVx6_ASAP7_75t_L g5913 ( 
.A(n_5614),
.Y(n_5913)
);

BUFx3_ASAP7_75t_L g5914 ( 
.A(n_5648),
.Y(n_5914)
);

CKINVDCx5p33_ASAP7_75t_R g5915 ( 
.A(n_5550),
.Y(n_5915)
);

AO21x1_ASAP7_75t_L g5916 ( 
.A1(n_5665),
.A2(n_5407),
.B(n_5363),
.Y(n_5916)
);

OAI21x1_ASAP7_75t_L g5917 ( 
.A1(n_5509),
.A2(n_5444),
.B(n_5364),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5604),
.Y(n_5918)
);

AO21x2_ASAP7_75t_L g5919 ( 
.A1(n_5542),
.A2(n_5363),
.B(n_5362),
.Y(n_5919)
);

OAI21x1_ASAP7_75t_L g5920 ( 
.A1(n_5493),
.A2(n_5523),
.B(n_5728),
.Y(n_5920)
);

OAI21x1_ASAP7_75t_L g5921 ( 
.A1(n_5515),
.A2(n_5337),
.B(n_5367),
.Y(n_5921)
);

OAI21x1_ASAP7_75t_L g5922 ( 
.A1(n_5480),
.A2(n_5437),
.B(n_5423),
.Y(n_5922)
);

AOI22x1_ASAP7_75t_L g5923 ( 
.A1(n_5526),
.A2(n_5665),
.B1(n_5474),
.B2(n_5483),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5611),
.Y(n_5924)
);

AOI21xp33_ASAP7_75t_L g5925 ( 
.A1(n_5757),
.A2(n_5362),
.B(n_5436),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5615),
.Y(n_5926)
);

OAI21x1_ASAP7_75t_L g5927 ( 
.A1(n_5464),
.A2(n_5436),
.B(n_5250),
.Y(n_5927)
);

CKINVDCx20_ASAP7_75t_R g5928 ( 
.A(n_5702),
.Y(n_5928)
);

OAI21x1_ASAP7_75t_L g5929 ( 
.A1(n_5463),
.A2(n_5250),
.B(n_5165),
.Y(n_5929)
);

AOI21x1_ASAP7_75t_L g5930 ( 
.A1(n_5461),
.A2(n_5257),
.B(n_5320),
.Y(n_5930)
);

BUFx12f_ASAP7_75t_L g5931 ( 
.A(n_5722),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5623),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5592),
.Y(n_5933)
);

AO21x2_ASAP7_75t_L g5934 ( 
.A1(n_5500),
.A2(n_5250),
.B(n_5320),
.Y(n_5934)
);

OAI21x1_ASAP7_75t_SL g5935 ( 
.A1(n_5777),
.A2(n_31),
.B(n_33),
.Y(n_5935)
);

INVx5_ASAP7_75t_L g5936 ( 
.A(n_5671),
.Y(n_5936)
);

NAND2x1p5_ASAP7_75t_L g5937 ( 
.A(n_5556),
.B(n_5184),
.Y(n_5937)
);

OAI22xp5_ASAP7_75t_L g5938 ( 
.A1(n_5752),
.A2(n_5184),
.B1(n_5231),
.B2(n_5202),
.Y(n_5938)
);

OAI21x1_ASAP7_75t_L g5939 ( 
.A1(n_5727),
.A2(n_5165),
.B(n_5241),
.Y(n_5939)
);

OAI21x1_ASAP7_75t_L g5940 ( 
.A1(n_5806),
.A2(n_5165),
.B(n_5241),
.Y(n_5940)
);

BUFx2_ASAP7_75t_L g5941 ( 
.A(n_5466),
.Y(n_5941)
);

OAI21xp5_ASAP7_75t_L g5942 ( 
.A1(n_5733),
.A2(n_5123),
.B(n_83),
.Y(n_5942)
);

BUFx12f_ASAP7_75t_L g5943 ( 
.A(n_5648),
.Y(n_5943)
);

AND2x4_ASAP7_75t_L g5944 ( 
.A(n_5592),
.B(n_5800),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5755),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5510),
.Y(n_5946)
);

OAI21x1_ASAP7_75t_L g5947 ( 
.A1(n_5666),
.A2(n_5241),
.B(n_5123),
.Y(n_5947)
);

OAI21x1_ASAP7_75t_L g5948 ( 
.A1(n_5685),
.A2(n_5123),
.B(n_5184),
.Y(n_5948)
);

AOI21xp5_ASAP7_75t_L g5949 ( 
.A1(n_5517),
.A2(n_5231),
.B(n_5202),
.Y(n_5949)
);

OAI21x1_ASAP7_75t_SL g5950 ( 
.A1(n_5470),
.A2(n_35),
.B(n_36),
.Y(n_5950)
);

AOI21x1_ASAP7_75t_L g5951 ( 
.A1(n_5580),
.A2(n_5231),
.B(n_5202),
.Y(n_5951)
);

OAI21x1_ASAP7_75t_L g5952 ( 
.A1(n_5804),
.A2(n_5390),
.B(n_5260),
.Y(n_5952)
);

NOR2xp33_ASAP7_75t_L g5953 ( 
.A(n_5767),
.B(n_5260),
.Y(n_5953)
);

BUFx6f_ASAP7_75t_L g5954 ( 
.A(n_5508),
.Y(n_5954)
);

OAI21x1_ASAP7_75t_L g5955 ( 
.A1(n_5706),
.A2(n_5390),
.B(n_5260),
.Y(n_5955)
);

AO21x2_ASAP7_75t_L g5956 ( 
.A1(n_5511),
.A2(n_5421),
.B(n_5390),
.Y(n_5956)
);

OAI21x1_ASAP7_75t_L g5957 ( 
.A1(n_5569),
.A2(n_5421),
.B(n_2200),
.Y(n_5957)
);

INVxp67_ASAP7_75t_SL g5958 ( 
.A(n_5472),
.Y(n_5958)
);

INVx3_ASAP7_75t_L g5959 ( 
.A(n_5697),
.Y(n_5959)
);

OA21x2_ASAP7_75t_L g5960 ( 
.A1(n_5762),
.A2(n_5421),
.B(n_35),
.Y(n_5960)
);

A2O1A1Ixp33_ASAP7_75t_L g5961 ( 
.A1(n_5717),
.A2(n_83),
.B(n_84),
.C(n_82),
.Y(n_5961)
);

CKINVDCx11_ASAP7_75t_R g5962 ( 
.A(n_5637),
.Y(n_5962)
);

OAI21x1_ASAP7_75t_L g5963 ( 
.A1(n_5590),
.A2(n_2200),
.B(n_2195),
.Y(n_5963)
);

INVx3_ASAP7_75t_L g5964 ( 
.A(n_5697),
.Y(n_5964)
);

INVx2_ASAP7_75t_L g5965 ( 
.A(n_5792),
.Y(n_5965)
);

INVx2_ASAP7_75t_SL g5966 ( 
.A(n_5540),
.Y(n_5966)
);

CKINVDCx14_ASAP7_75t_R g5967 ( 
.A(n_5779),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5536),
.Y(n_5968)
);

HB1xp67_ASAP7_75t_L g5969 ( 
.A(n_5536),
.Y(n_5969)
);

OA21x2_ASAP7_75t_L g5970 ( 
.A1(n_5608),
.A2(n_36),
.B(n_38),
.Y(n_5970)
);

O2A1O1Ixp33_ASAP7_75t_L g5971 ( 
.A1(n_5735),
.A2(n_86),
.B(n_87),
.C(n_85),
.Y(n_5971)
);

INVx1_ASAP7_75t_SL g5972 ( 
.A(n_5792),
.Y(n_5972)
);

INVx5_ASAP7_75t_L g5973 ( 
.A(n_5671),
.Y(n_5973)
);

OAI21x1_ASAP7_75t_L g5974 ( 
.A1(n_5605),
.A2(n_2200),
.B(n_2195),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5536),
.Y(n_5975)
);

OAI21x1_ASAP7_75t_L g5976 ( 
.A1(n_5781),
.A2(n_2210),
.B(n_2195),
.Y(n_5976)
);

OAI21x1_ASAP7_75t_SL g5977 ( 
.A1(n_5512),
.A2(n_38),
.B(n_39),
.Y(n_5977)
);

NAND2x1p5_ASAP7_75t_L g5978 ( 
.A(n_5556),
.B(n_3166),
.Y(n_5978)
);

NAND3xp33_ASAP7_75t_L g5979 ( 
.A(n_5796),
.B(n_86),
.C(n_85),
.Y(n_5979)
);

BUFx2_ASAP7_75t_R g5980 ( 
.A(n_5674),
.Y(n_5980)
);

OAI21x1_ASAP7_75t_L g5981 ( 
.A1(n_5775),
.A2(n_2224),
.B(n_2210),
.Y(n_5981)
);

NAND2xp5_ASAP7_75t_SL g5982 ( 
.A(n_5558),
.B(n_5596),
.Y(n_5982)
);

OAI21x1_ASAP7_75t_L g5983 ( 
.A1(n_5760),
.A2(n_2224),
.B(n_2210),
.Y(n_5983)
);

OR2x6_ASAP7_75t_L g5984 ( 
.A(n_5771),
.B(n_3166),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5527),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5751),
.Y(n_5986)
);

OA21x2_ASAP7_75t_L g5987 ( 
.A1(n_5757),
.A2(n_39),
.B(n_40),
.Y(n_5987)
);

OAI21x1_ASAP7_75t_L g5988 ( 
.A1(n_5524),
.A2(n_2224),
.B(n_2210),
.Y(n_5988)
);

OAI21x1_ASAP7_75t_L g5989 ( 
.A1(n_5625),
.A2(n_2229),
.B(n_2224),
.Y(n_5989)
);

AND2x2_ASAP7_75t_L g5990 ( 
.A(n_5670),
.B(n_40),
.Y(n_5990)
);

OAI21x1_ASAP7_75t_L g5991 ( 
.A1(n_5625),
.A2(n_2232),
.B(n_2229),
.Y(n_5991)
);

NAND3xp33_ASAP7_75t_L g5992 ( 
.A(n_5668),
.B(n_89),
.C(n_88),
.Y(n_5992)
);

OR2x2_ASAP7_75t_L g5993 ( 
.A(n_5756),
.B(n_5773),
.Y(n_5993)
);

INVx4_ASAP7_75t_L g5994 ( 
.A(n_5521),
.Y(n_5994)
);

BUFx2_ASAP7_75t_SL g5995 ( 
.A(n_5637),
.Y(n_5995)
);

AO21x2_ASAP7_75t_L g5996 ( 
.A1(n_5552),
.A2(n_40),
.B(n_41),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5460),
.Y(n_5997)
);

OAI21x1_ASAP7_75t_SL g5998 ( 
.A1(n_5532),
.A2(n_5575),
.B(n_5567),
.Y(n_5998)
);

BUFx12f_ASAP7_75t_L g5999 ( 
.A(n_5606),
.Y(n_5999)
);

BUFx2_ASAP7_75t_L g6000 ( 
.A(n_5528),
.Y(n_6000)
);

OR3x4_ASAP7_75t_SL g6001 ( 
.A(n_5764),
.B(n_5731),
.C(n_5726),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5460),
.B(n_42),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5460),
.Y(n_6003)
);

OAI21x1_ASAP7_75t_L g6004 ( 
.A1(n_5690),
.A2(n_5659),
.B(n_5657),
.Y(n_6004)
);

AOI22xp5_ASAP7_75t_L g6005 ( 
.A1(n_5745),
.A2(n_90),
.B1(n_91),
.B2(n_88),
.Y(n_6005)
);

AO21x2_ASAP7_75t_L g6006 ( 
.A1(n_5552),
.A2(n_42),
.B(n_43),
.Y(n_6006)
);

OA21x2_ASAP7_75t_L g6007 ( 
.A1(n_5476),
.A2(n_43),
.B(n_44),
.Y(n_6007)
);

OA21x2_ASAP7_75t_L g6008 ( 
.A1(n_5499),
.A2(n_5551),
.B(n_5545),
.Y(n_6008)
);

OAI21x1_ASAP7_75t_L g6009 ( 
.A1(n_5644),
.A2(n_2232),
.B(n_2229),
.Y(n_6009)
);

BUFx2_ASAP7_75t_R g6010 ( 
.A(n_5467),
.Y(n_6010)
);

AOI21xp5_ASAP7_75t_L g6011 ( 
.A1(n_5662),
.A2(n_3232),
.B(n_3166),
.Y(n_6011)
);

INVx2_ASAP7_75t_SL g6012 ( 
.A(n_5508),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5609),
.Y(n_6013)
);

OA21x2_ASAP7_75t_L g6014 ( 
.A1(n_5634),
.A2(n_44),
.B(n_45),
.Y(n_6014)
);

AO21x2_ASAP7_75t_L g6015 ( 
.A1(n_5708),
.A2(n_44),
.B(n_45),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5484),
.Y(n_6016)
);

AND2x4_ASAP7_75t_L g6017 ( 
.A(n_5558),
.B(n_46),
.Y(n_6017)
);

INVx2_ASAP7_75t_SL g6018 ( 
.A(n_5508),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5484),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5676),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5484),
.Y(n_6021)
);

BUFx2_ASAP7_75t_L g6022 ( 
.A(n_5676),
.Y(n_6022)
);

BUFx2_ASAP7_75t_SL g6023 ( 
.A(n_5700),
.Y(n_6023)
);

OAI21x1_ASAP7_75t_L g6024 ( 
.A1(n_5618),
.A2(n_2232),
.B(n_2229),
.Y(n_6024)
);

OAI21x1_ASAP7_75t_SL g6025 ( 
.A1(n_5663),
.A2(n_46),
.B(n_47),
.Y(n_6025)
);

OAI21xp5_ASAP7_75t_L g6026 ( 
.A1(n_5495),
.A2(n_92),
.B(n_90),
.Y(n_6026)
);

BUFx3_ASAP7_75t_L g6027 ( 
.A(n_5676),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5776),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5521),
.Y(n_6029)
);

OR2x2_ASAP7_75t_L g6030 ( 
.A(n_5707),
.B(n_47),
.Y(n_6030)
);

OA21x2_ASAP7_75t_L g6031 ( 
.A1(n_5797),
.A2(n_47),
.B(n_48),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5596),
.Y(n_6032)
);

AO21x1_ASAP7_75t_L g6033 ( 
.A1(n_5597),
.A2(n_48),
.B(n_49),
.Y(n_6033)
);

AO21x2_ASAP7_75t_L g6034 ( 
.A1(n_5708),
.A2(n_48),
.B(n_50),
.Y(n_6034)
);

HB1xp67_ASAP7_75t_L g6035 ( 
.A(n_5653),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5776),
.Y(n_6036)
);

OAI21x1_ASAP7_75t_L g6037 ( 
.A1(n_5765),
.A2(n_2234),
.B(n_2232),
.Y(n_6037)
);

AOI21xp5_ASAP7_75t_L g6038 ( 
.A1(n_5681),
.A2(n_3232),
.B(n_3166),
.Y(n_6038)
);

OAI21xp5_ASAP7_75t_L g6039 ( 
.A1(n_5495),
.A2(n_5504),
.B(n_5572),
.Y(n_6039)
);

OAI21x1_ASAP7_75t_L g6040 ( 
.A1(n_5787),
.A2(n_2234),
.B(n_2110),
.Y(n_6040)
);

BUFx3_ASAP7_75t_L g6041 ( 
.A(n_5462),
.Y(n_6041)
);

INVx5_ASAP7_75t_L g6042 ( 
.A(n_5479),
.Y(n_6042)
);

OAI22xp5_ASAP7_75t_L g6043 ( 
.A1(n_5752),
.A2(n_95),
.B1(n_114),
.B2(n_104),
.Y(n_6043)
);

HB1xp67_ASAP7_75t_L g6044 ( 
.A(n_5653),
.Y(n_6044)
);

BUFx3_ASAP7_75t_L g6045 ( 
.A(n_5801),
.Y(n_6045)
);

OR2x2_ASAP7_75t_L g6046 ( 
.A(n_5744),
.B(n_50),
.Y(n_6046)
);

NOR2x1_ASAP7_75t_R g6047 ( 
.A(n_5801),
.B(n_50),
.Y(n_6047)
);

NAND2x1p5_ASAP7_75t_L g6048 ( 
.A(n_5558),
.B(n_3232),
.Y(n_6048)
);

AND2x4_ASAP7_75t_L g6049 ( 
.A(n_5539),
.B(n_51),
.Y(n_6049)
);

OAI21x1_ASAP7_75t_L g6050 ( 
.A1(n_5742),
.A2(n_2234),
.B(n_2110),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5776),
.Y(n_6051)
);

AO21x2_ASAP7_75t_L g6052 ( 
.A1(n_5729),
.A2(n_51),
.B(n_52),
.Y(n_6052)
);

OAI21x1_ASAP7_75t_L g6053 ( 
.A1(n_5574),
.A2(n_2234),
.B(n_2110),
.Y(n_6053)
);

AOI22xp5_ASAP7_75t_L g6054 ( 
.A1(n_5745),
.A2(n_93),
.B1(n_97),
.B2(n_96),
.Y(n_6054)
);

OAI21x1_ASAP7_75t_L g6055 ( 
.A1(n_5574),
.A2(n_2110),
.B(n_2098),
.Y(n_6055)
);

OAI21x1_ASAP7_75t_L g6056 ( 
.A1(n_5664),
.A2(n_2146),
.B(n_2098),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5780),
.Y(n_6057)
);

INVx8_ASAP7_75t_L g6058 ( 
.A(n_5539),
.Y(n_6058)
);

OA21x2_ASAP7_75t_L g6059 ( 
.A1(n_5747),
.A2(n_52),
.B(n_53),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5780),
.Y(n_6060)
);

BUFx10_ASAP7_75t_L g6061 ( 
.A(n_5497),
.Y(n_6061)
);

BUFx3_ASAP7_75t_L g6062 ( 
.A(n_5788),
.Y(n_6062)
);

OA21x2_ASAP7_75t_L g6063 ( 
.A1(n_5538),
.A2(n_52),
.B(n_53),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_5687),
.B(n_53),
.Y(n_6064)
);

INVx3_ASAP7_75t_L g6065 ( 
.A(n_5479),
.Y(n_6065)
);

CKINVDCx5p33_ASAP7_75t_R g6066 ( 
.A(n_5672),
.Y(n_6066)
);

INVx2_ASAP7_75t_SL g6067 ( 
.A(n_5573),
.Y(n_6067)
);

NAND3xp33_ASAP7_75t_L g6068 ( 
.A(n_5793),
.B(n_96),
.C(n_93),
.Y(n_6068)
);

OR2x6_ASAP7_75t_L g6069 ( 
.A(n_5761),
.B(n_3232),
.Y(n_6069)
);

OAI21xp5_ASAP7_75t_L g6070 ( 
.A1(n_5504),
.A2(n_100),
.B(n_99),
.Y(n_6070)
);

OAI221xp5_ASAP7_75t_L g6071 ( 
.A1(n_5717),
.A2(n_54),
.B1(n_56),
.B2(n_55),
.C(n_99),
.Y(n_6071)
);

OAI21x1_ASAP7_75t_L g6072 ( 
.A1(n_5691),
.A2(n_2146),
.B(n_2098),
.Y(n_6072)
);

CKINVDCx20_ASAP7_75t_R g6073 ( 
.A(n_5791),
.Y(n_6073)
);

OAI21x1_ASAP7_75t_SL g6074 ( 
.A1(n_5684),
.A2(n_54),
.B(n_100),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_5687),
.B(n_54),
.Y(n_6075)
);

OAI21x1_ASAP7_75t_L g6076 ( 
.A1(n_5516),
.A2(n_2146),
.B(n_2098),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5780),
.Y(n_6077)
);

INVx1_ASAP7_75t_SL g6078 ( 
.A(n_5761),
.Y(n_6078)
);

OAI21x1_ASAP7_75t_SL g6079 ( 
.A1(n_5686),
.A2(n_101),
.B(n_102),
.Y(n_6079)
);

BUFx3_ASAP7_75t_L g6080 ( 
.A(n_5479),
.Y(n_6080)
);

INVx2_ASAP7_75t_L g6081 ( 
.A(n_5573),
.Y(n_6081)
);

BUFx2_ASAP7_75t_R g6082 ( 
.A(n_5576),
.Y(n_6082)
);

NOR2xp33_ASAP7_75t_L g6083 ( 
.A(n_5562),
.B(n_5688),
.Y(n_6083)
);

CKINVDCx5p33_ASAP7_75t_R g6084 ( 
.A(n_5502),
.Y(n_6084)
);

OAI21xp5_ASAP7_75t_L g6085 ( 
.A1(n_5703),
.A2(n_101),
.B(n_102),
.Y(n_6085)
);

BUFx3_ASAP7_75t_L g6086 ( 
.A(n_5479),
.Y(n_6086)
);

NAND2x1p5_ASAP7_75t_L g6087 ( 
.A(n_5586),
.B(n_3232),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5790),
.Y(n_6088)
);

AO21x2_ASAP7_75t_L g6089 ( 
.A1(n_5729),
.A2(n_113),
.B(n_103),
.Y(n_6089)
);

AO21x2_ASAP7_75t_L g6090 ( 
.A1(n_5750),
.A2(n_116),
.B(n_104),
.Y(n_6090)
);

NOR2xp67_ASAP7_75t_L g6091 ( 
.A(n_5772),
.B(n_106),
.Y(n_6091)
);

BUFx10_ASAP7_75t_L g6092 ( 
.A(n_5642),
.Y(n_6092)
);

OAI21x1_ASAP7_75t_L g6093 ( 
.A1(n_5930),
.A2(n_5586),
.B(n_5643),
.Y(n_6093)
);

AO31x2_ASAP7_75t_L g6094 ( 
.A1(n_6028),
.A2(n_5560),
.A3(n_5640),
.B(n_5595),
.Y(n_6094)
);

AND2x4_ASAP7_75t_L g6095 ( 
.A(n_6065),
.B(n_5750),
.Y(n_6095)
);

OAI21x1_ASAP7_75t_L g6096 ( 
.A1(n_5955),
.A2(n_5651),
.B(n_5768),
.Y(n_6096)
);

OAI21x1_ASAP7_75t_L g6097 ( 
.A1(n_5829),
.A2(n_5566),
.B(n_5492),
.Y(n_6097)
);

NAND2xp5_ASAP7_75t_L g6098 ( 
.A(n_5958),
.B(n_5769),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5855),
.Y(n_6099)
);

OA21x2_ASAP7_75t_L g6100 ( 
.A1(n_5825),
.A2(n_5698),
.B(n_5695),
.Y(n_6100)
);

OR2x2_ASAP7_75t_L g6101 ( 
.A(n_5958),
.B(n_5878),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5853),
.Y(n_6102)
);

AO21x2_ASAP7_75t_L g6103 ( 
.A1(n_5825),
.A2(n_5769),
.B(n_5487),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5853),
.Y(n_6104)
);

INVx1_ASAP7_75t_L g6105 ( 
.A(n_5868),
.Y(n_6105)
);

NAND2x1p5_ASAP7_75t_L g6106 ( 
.A(n_6042),
.B(n_5982),
.Y(n_6106)
);

INVx2_ASAP7_75t_L g6107 ( 
.A(n_5855),
.Y(n_6107)
);

OAI21x1_ASAP7_75t_L g6108 ( 
.A1(n_5817),
.A2(n_5770),
.B(n_5766),
.Y(n_6108)
);

AOI21xp5_ASAP7_75t_L g6109 ( 
.A1(n_6039),
.A2(n_5725),
.B(n_5696),
.Y(n_6109)
);

OAI21x1_ASAP7_75t_L g6110 ( 
.A1(n_6002),
.A2(n_5478),
.B(n_5563),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_5946),
.B(n_5660),
.Y(n_6111)
);

OA21x2_ASAP7_75t_L g6112 ( 
.A1(n_6039),
.A2(n_5854),
.B(n_6036),
.Y(n_6112)
);

OAI21x1_ASAP7_75t_L g6113 ( 
.A1(n_6002),
.A2(n_5669),
.B(n_5719),
.Y(n_6113)
);

NAND2x1p5_ASAP7_75t_L g6114 ( 
.A(n_6042),
.B(n_5721),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5868),
.Y(n_6115)
);

OAI21x1_ASAP7_75t_L g6116 ( 
.A1(n_5900),
.A2(n_5531),
.B(n_5530),
.Y(n_6116)
);

A2O1A1Ixp33_ASAP7_75t_L g6117 ( 
.A1(n_6070),
.A2(n_5546),
.B(n_5559),
.C(n_5738),
.Y(n_6117)
);

AND2x4_ASAP7_75t_L g6118 ( 
.A(n_6065),
.B(n_5525),
.Y(n_6118)
);

AO21x2_ASAP7_75t_L g6119 ( 
.A1(n_6064),
.A2(n_5559),
.B(n_5546),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_5827),
.Y(n_6120)
);

INVx3_ASAP7_75t_L g6121 ( 
.A(n_5823),
.Y(n_6121)
);

BUFx12f_ASAP7_75t_L g6122 ( 
.A(n_5962),
.Y(n_6122)
);

AOI21xp5_ASAP7_75t_L g6123 ( 
.A1(n_6070),
.A2(n_5715),
.B(n_5710),
.Y(n_6123)
);

OA21x2_ASAP7_75t_L g6124 ( 
.A1(n_5854),
.A2(n_5795),
.B(n_5786),
.Y(n_6124)
);

AOI21x1_ASAP7_75t_L g6125 ( 
.A1(n_5885),
.A2(n_5805),
.B(n_5802),
.Y(n_6125)
);

AO21x2_ASAP7_75t_L g6126 ( 
.A1(n_6064),
.A2(n_5683),
.B(n_5557),
.Y(n_6126)
);

BUFx2_ASAP7_75t_L g6127 ( 
.A(n_5864),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5842),
.Y(n_6128)
);

BUFx3_ASAP7_75t_L g6129 ( 
.A(n_5931),
.Y(n_6129)
);

OAI21x1_ASAP7_75t_L g6130 ( 
.A1(n_5900),
.A2(n_5535),
.B(n_5568),
.Y(n_6130)
);

OAI21x1_ASAP7_75t_L g6131 ( 
.A1(n_5847),
.A2(n_5675),
.B(n_5667),
.Y(n_6131)
);

OA21x2_ASAP7_75t_L g6132 ( 
.A1(n_6051),
.A2(n_5639),
.B(n_5635),
.Y(n_6132)
);

AO31x2_ASAP7_75t_L g6133 ( 
.A1(n_6057),
.A2(n_5587),
.A3(n_5624),
.B(n_5579),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_5816),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_5842),
.Y(n_6135)
);

OR2x2_ASAP7_75t_L g6136 ( 
.A(n_5993),
.B(n_5687),
.Y(n_6136)
);

INVx3_ASAP7_75t_L g6137 ( 
.A(n_5823),
.Y(n_6137)
);

NOR2xp33_ASAP7_75t_L g6138 ( 
.A(n_5812),
.B(n_5496),
.Y(n_6138)
);

CKINVDCx20_ASAP7_75t_R g6139 ( 
.A(n_5928),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5873),
.Y(n_6140)
);

AOI21x1_ASAP7_75t_L g6141 ( 
.A1(n_5808),
.A2(n_5649),
.B(n_5645),
.Y(n_6141)
);

OAI21xp5_ASAP7_75t_L g6142 ( 
.A1(n_5967),
.A2(n_5759),
.B(n_5518),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5818),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5828),
.Y(n_6144)
);

BUFx2_ASAP7_75t_L g6145 ( 
.A(n_5864),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5834),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_5873),
.Y(n_6147)
);

OA21x2_ASAP7_75t_L g6148 ( 
.A1(n_6060),
.A2(n_5689),
.B(n_5678),
.Y(n_6148)
);

OAI21x1_ASAP7_75t_L g6149 ( 
.A1(n_5847),
.A2(n_5692),
.B(n_5583),
.Y(n_6149)
);

OAI21x1_ASAP7_75t_L g6150 ( 
.A1(n_5874),
.A2(n_5612),
.B(n_5513),
.Y(n_6150)
);

NAND2xp5_ASAP7_75t_L g6151 ( 
.A(n_5857),
.B(n_5555),
.Y(n_6151)
);

OA21x2_ASAP7_75t_L g6152 ( 
.A1(n_6077),
.A2(n_5656),
.B(n_5565),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_5836),
.Y(n_6153)
);

NOR2xp33_ASAP7_75t_L g6154 ( 
.A(n_5812),
.B(n_5554),
.Y(n_6154)
);

AOI21x1_ASAP7_75t_L g6155 ( 
.A1(n_5902),
.A2(n_5730),
.B(n_5617),
.Y(n_6155)
);

AOI22xp33_ASAP7_75t_L g6156 ( 
.A1(n_5967),
.A2(n_5741),
.B1(n_5718),
.B2(n_5600),
.Y(n_6156)
);

OAI21x1_ASAP7_75t_L g6157 ( 
.A1(n_5874),
.A2(n_5582),
.B(n_5577),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5838),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_5840),
.Y(n_6159)
);

INVx3_ASAP7_75t_L g6160 ( 
.A(n_5831),
.Y(n_6160)
);

AOI21x1_ASAP7_75t_L g6161 ( 
.A1(n_6075),
.A2(n_5732),
.B(n_5711),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5844),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_5909),
.Y(n_6163)
);

BUFx3_ASAP7_75t_L g6164 ( 
.A(n_5943),
.Y(n_6164)
);

AO21x1_ASAP7_75t_L g6165 ( 
.A1(n_6088),
.A2(n_5790),
.B(n_5564),
.Y(n_6165)
);

NAND2xp5_ASAP7_75t_L g6166 ( 
.A(n_5826),
.B(n_5555),
.Y(n_6166)
);

OAI21x1_ASAP7_75t_L g6167 ( 
.A1(n_5997),
.A2(n_5584),
.B(n_5571),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5850),
.Y(n_6168)
);

NAND2xp5_ASAP7_75t_L g6169 ( 
.A(n_5826),
.B(n_5555),
.Y(n_6169)
);

OR2x2_ASAP7_75t_L g6170 ( 
.A(n_5886),
.B(n_5653),
.Y(n_6170)
);

NAND2xp5_ASAP7_75t_L g6171 ( 
.A(n_5880),
.B(n_5741),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5909),
.Y(n_6172)
);

AOI22xp33_ASAP7_75t_L g6173 ( 
.A1(n_5856),
.A2(n_5718),
.B1(n_5600),
.B2(n_5489),
.Y(n_6173)
);

OA21x2_ASAP7_75t_L g6174 ( 
.A1(n_6003),
.A2(n_5578),
.B(n_5622),
.Y(n_6174)
);

NAND2xp5_ASAP7_75t_L g6175 ( 
.A(n_6013),
.B(n_5564),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5933),
.Y(n_6176)
);

OA21x2_ASAP7_75t_L g6177 ( 
.A1(n_6075),
.A2(n_5886),
.B(n_5821),
.Y(n_6177)
);

INVx3_ASAP7_75t_L g6178 ( 
.A(n_5831),
.Y(n_6178)
);

BUFx3_ASAP7_75t_L g6179 ( 
.A(n_5928),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_5851),
.Y(n_6180)
);

OAI21x1_ASAP7_75t_L g6181 ( 
.A1(n_5875),
.A2(n_5891),
.B(n_5876),
.Y(n_6181)
);

OA21x2_ASAP7_75t_L g6182 ( 
.A1(n_5920),
.A2(n_5522),
.B(n_5544),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5860),
.Y(n_6183)
);

OAI21x1_ASAP7_75t_L g6184 ( 
.A1(n_5948),
.A2(n_5607),
.B(n_5589),
.Y(n_6184)
);

OAI21x1_ASAP7_75t_L g6185 ( 
.A1(n_5937),
.A2(n_5929),
.B(n_5982),
.Y(n_6185)
);

AO21x2_ASAP7_75t_L g6186 ( 
.A1(n_6033),
.A2(n_5790),
.B(n_5734),
.Y(n_6186)
);

AND2x4_ASAP7_75t_L g6187 ( 
.A(n_6042),
.B(n_5525),
.Y(n_6187)
);

OAI21xp5_ASAP7_75t_L g6188 ( 
.A1(n_6026),
.A2(n_5784),
.B(n_5721),
.Y(n_6188)
);

OAI21x1_ASAP7_75t_L g6189 ( 
.A1(n_5937),
.A2(n_5661),
.B(n_5753),
.Y(n_6189)
);

AO21x1_ASAP7_75t_L g6190 ( 
.A1(n_6043),
.A2(n_5638),
.B(n_5491),
.Y(n_6190)
);

OR2x6_ASAP7_75t_L g6191 ( 
.A(n_5995),
.B(n_5621),
.Y(n_6191)
);

AOI21xp5_ASAP7_75t_L g6192 ( 
.A1(n_5859),
.A2(n_5646),
.B(n_5778),
.Y(n_6192)
);

OAI22xp5_ASAP7_75t_L g6193 ( 
.A1(n_6010),
.A2(n_5603),
.B1(n_5632),
.B2(n_5620),
.Y(n_6193)
);

AND2x2_ASAP7_75t_L g6194 ( 
.A(n_5830),
.B(n_5525),
.Y(n_6194)
);

AND2x4_ASAP7_75t_L g6195 ( 
.A(n_6042),
.B(n_5716),
.Y(n_6195)
);

AOI21x1_ASAP7_75t_L g6196 ( 
.A1(n_5908),
.A2(n_5620),
.B(n_5603),
.Y(n_6196)
);

OAI21x1_ASAP7_75t_L g6197 ( 
.A1(n_5892),
.A2(n_5758),
.B(n_5534),
.Y(n_6197)
);

AND2x4_ASAP7_75t_L g6198 ( 
.A(n_6080),
.B(n_5716),
.Y(n_6198)
);

AND2x2_ASAP7_75t_L g6199 ( 
.A(n_5941),
.B(n_5716),
.Y(n_6199)
);

OAI21x1_ASAP7_75t_L g6200 ( 
.A1(n_5884),
.A2(n_5673),
.B(n_5547),
.Y(n_6200)
);

OAI21x1_ASAP7_75t_SL g6201 ( 
.A1(n_5916),
.A2(n_5782),
.B(n_5789),
.Y(n_6201)
);

OAI21x1_ASAP7_75t_SL g6202 ( 
.A1(n_5950),
.A2(n_108),
.B(n_109),
.Y(n_6202)
);

INVx2_ASAP7_75t_L g6203 ( 
.A(n_5918),
.Y(n_6203)
);

INVx2_ASAP7_75t_SL g6204 ( 
.A(n_5824),
.Y(n_6204)
);

OAI21x1_ASAP7_75t_SL g6205 ( 
.A1(n_5856),
.A2(n_109),
.B(n_110),
.Y(n_6205)
);

OAI21xp5_ASAP7_75t_L g6206 ( 
.A1(n_6026),
.A2(n_5632),
.B(n_5489),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_5965),
.Y(n_6207)
);

OR2x2_ASAP7_75t_L g6208 ( 
.A(n_5810),
.B(n_5588),
.Y(n_6208)
);

INVxp33_ASAP7_75t_L g6209 ( 
.A(n_5962),
.Y(n_6209)
);

NOR2xp33_ASAP7_75t_L g6210 ( 
.A(n_5887),
.B(n_110),
.Y(n_6210)
);

AO21x2_ASAP7_75t_L g6211 ( 
.A1(n_5910),
.A2(n_111),
.B(n_112),
.Y(n_6211)
);

OAI21x1_ASAP7_75t_L g6212 ( 
.A1(n_5947),
.A2(n_2156),
.B(n_2146),
.Y(n_6212)
);

AND2x4_ASAP7_75t_L g6213 ( 
.A(n_6086),
.B(n_115),
.Y(n_6213)
);

OR2x6_ASAP7_75t_L g6214 ( 
.A(n_6023),
.B(n_3260),
.Y(n_6214)
);

OAI21x1_ASAP7_75t_L g6215 ( 
.A1(n_5897),
.A2(n_2156),
.B(n_115),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5863),
.Y(n_6216)
);

AO21x2_ASAP7_75t_L g6217 ( 
.A1(n_5910),
.A2(n_117),
.B(n_118),
.Y(n_6217)
);

OA21x2_ASAP7_75t_L g6218 ( 
.A1(n_5903),
.A2(n_117),
.B(n_120),
.Y(n_6218)
);

OAI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_6068),
.A2(n_121),
.B(n_122),
.Y(n_6219)
);

OR2x2_ASAP7_75t_L g6220 ( 
.A(n_5945),
.B(n_123),
.Y(n_6220)
);

OAI21xp5_ASAP7_75t_L g6221 ( 
.A1(n_6068),
.A2(n_123),
.B(n_124),
.Y(n_6221)
);

AOI21xp5_ASAP7_75t_L g6222 ( 
.A1(n_5859),
.A2(n_124),
.B(n_125),
.Y(n_6222)
);

HB1xp67_ASAP7_75t_L g6223 ( 
.A(n_5841),
.Y(n_6223)
);

AO31x2_ASAP7_75t_L g6224 ( 
.A1(n_6043),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_6224)
);

NOR2x1_ASAP7_75t_R g6225 ( 
.A(n_5999),
.B(n_126),
.Y(n_6225)
);

BUFx6f_ASAP7_75t_L g6226 ( 
.A(n_5811),
.Y(n_6226)
);

AOI21x1_ASAP7_75t_L g6227 ( 
.A1(n_5815),
.A2(n_127),
.B(n_129),
.Y(n_6227)
);

AOI21x1_ASAP7_75t_L g6228 ( 
.A1(n_5820),
.A2(n_130),
.B(n_132),
.Y(n_6228)
);

OAI21x1_ASAP7_75t_SL g6229 ( 
.A1(n_5998),
.A2(n_134),
.B(n_135),
.Y(n_6229)
);

AO21x2_ASAP7_75t_L g6230 ( 
.A1(n_5935),
.A2(n_135),
.B(n_136),
.Y(n_6230)
);

BUFx8_ASAP7_75t_L g6231 ( 
.A(n_5990),
.Y(n_6231)
);

OR2x2_ASAP7_75t_L g6232 ( 
.A(n_5986),
.B(n_136),
.Y(n_6232)
);

OAI21xp5_ASAP7_75t_L g6233 ( 
.A1(n_5979),
.A2(n_137),
.B(n_138),
.Y(n_6233)
);

OAI21x1_ASAP7_75t_SL g6234 ( 
.A1(n_5871),
.A2(n_139),
.B(n_141),
.Y(n_6234)
);

OAI21xp5_ASAP7_75t_L g6235 ( 
.A1(n_6083),
.A2(n_139),
.B(n_141),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_5924),
.Y(n_6236)
);

AOI21xp5_ASAP7_75t_L g6237 ( 
.A1(n_5971),
.A2(n_142),
.B(n_144),
.Y(n_6237)
);

AOI21xp5_ASAP7_75t_SL g6238 ( 
.A1(n_6007),
.A2(n_5960),
.B(n_6017),
.Y(n_6238)
);

OAI21x1_ASAP7_75t_L g6239 ( 
.A1(n_5939),
.A2(n_2156),
.B(n_142),
.Y(n_6239)
);

AO21x2_ASAP7_75t_L g6240 ( 
.A1(n_5968),
.A2(n_144),
.B(n_145),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_5877),
.B(n_145),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_5926),
.Y(n_6242)
);

AO31x2_ASAP7_75t_L g6243 ( 
.A1(n_5975),
.A2(n_148),
.A3(n_146),
.B(n_147),
.Y(n_6243)
);

OAI21x1_ASAP7_75t_L g6244 ( 
.A1(n_6087),
.A2(n_2156),
.B(n_146),
.Y(n_6244)
);

NOR2xp33_ASAP7_75t_L g6245 ( 
.A(n_5887),
.B(n_147),
.Y(n_6245)
);

AO21x2_ASAP7_75t_L g6246 ( 
.A1(n_5837),
.A2(n_5809),
.B(n_6016),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_L g6247 ( 
.A(n_5837),
.B(n_148),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5959),
.Y(n_6248)
);

OAI21x1_ASAP7_75t_L g6249 ( 
.A1(n_6087),
.A2(n_149),
.B(n_150),
.Y(n_6249)
);

CKINVDCx20_ASAP7_75t_R g6250 ( 
.A(n_5819),
.Y(n_6250)
);

OAI21x1_ASAP7_75t_L g6251 ( 
.A1(n_5849),
.A2(n_5940),
.B(n_5895),
.Y(n_6251)
);

OA21x2_ASAP7_75t_L g6252 ( 
.A1(n_5932),
.A2(n_149),
.B(n_151),
.Y(n_6252)
);

OAI21xp5_ASAP7_75t_L g6253 ( 
.A1(n_6083),
.A2(n_152),
.B(n_153),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_5959),
.Y(n_6254)
);

NAND2xp5_ASAP7_75t_L g6255 ( 
.A(n_5985),
.B(n_152),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5813),
.Y(n_6256)
);

AO21x1_ASAP7_75t_L g6257 ( 
.A1(n_6017),
.A2(n_153),
.B(n_154),
.Y(n_6257)
);

NAND3xp33_ASAP7_75t_L g6258 ( 
.A(n_5979),
.B(n_155),
.C(n_156),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5869),
.Y(n_6259)
);

OAI21x1_ASAP7_75t_L g6260 ( 
.A1(n_5849),
.A2(n_155),
.B(n_157),
.Y(n_6260)
);

NAND2x1_ASAP7_75t_L g6261 ( 
.A(n_5862),
.B(n_3260),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_5870),
.Y(n_6262)
);

HB1xp67_ASAP7_75t_L g6263 ( 
.A(n_5841),
.Y(n_6263)
);

OAI21x1_ASAP7_75t_L g6264 ( 
.A1(n_6004),
.A2(n_158),
.B(n_159),
.Y(n_6264)
);

BUFx8_ASAP7_75t_SL g6265 ( 
.A(n_5915),
.Y(n_6265)
);

NOR2xp33_ASAP7_75t_L g6266 ( 
.A(n_5887),
.B(n_158),
.Y(n_6266)
);

AOI21xp5_ASAP7_75t_L g6267 ( 
.A1(n_5971),
.A2(n_160),
.B(n_161),
.Y(n_6267)
);

OR2x6_ASAP7_75t_L g6268 ( 
.A(n_5824),
.B(n_3260),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5904),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5906),
.Y(n_6270)
);

NAND2xp5_ASAP7_75t_L g6271 ( 
.A(n_6008),
.B(n_161),
.Y(n_6271)
);

OAI21x1_ASAP7_75t_L g6272 ( 
.A1(n_5905),
.A2(n_162),
.B(n_165),
.Y(n_6272)
);

INVx1_ASAP7_75t_L g6273 ( 
.A(n_5866),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5894),
.Y(n_6274)
);

AOI21xp5_ASAP7_75t_L g6275 ( 
.A1(n_6085),
.A2(n_162),
.B(n_165),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_5861),
.Y(n_6276)
);

OAI21x1_ASAP7_75t_L g6277 ( 
.A1(n_5890),
.A2(n_5927),
.B(n_5952),
.Y(n_6277)
);

NAND2xp5_ASAP7_75t_L g6278 ( 
.A(n_6008),
.B(n_167),
.Y(n_6278)
);

AND2x2_ASAP7_75t_L g6279 ( 
.A(n_5872),
.B(n_168),
.Y(n_6279)
);

OA21x2_ASAP7_75t_L g6280 ( 
.A1(n_5893),
.A2(n_170),
.B(n_171),
.Y(n_6280)
);

AO21x2_ASAP7_75t_L g6281 ( 
.A1(n_5809),
.A2(n_171),
.B(n_172),
.Y(n_6281)
);

NAND2x1p5_ASAP7_75t_L g6282 ( 
.A(n_5936),
.B(n_3260),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_5867),
.Y(n_6283)
);

OAI21xp5_ASAP7_75t_L g6284 ( 
.A1(n_6085),
.A2(n_173),
.B(n_174),
.Y(n_6284)
);

OAI21x1_ASAP7_75t_L g6285 ( 
.A1(n_5951),
.A2(n_175),
.B(n_176),
.Y(n_6285)
);

AOI21xp5_ASAP7_75t_L g6286 ( 
.A1(n_5992),
.A2(n_178),
.B(n_179),
.Y(n_6286)
);

BUFx6f_ASAP7_75t_L g6287 ( 
.A(n_5811),
.Y(n_6287)
);

NOR2xp67_ASAP7_75t_L g6288 ( 
.A(n_5811),
.B(n_5936),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_5867),
.Y(n_6289)
);

HB1xp67_ASAP7_75t_L g6290 ( 
.A(n_5893),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5867),
.Y(n_6291)
);

OAI21x1_ASAP7_75t_L g6292 ( 
.A1(n_5865),
.A2(n_179),
.B(n_180),
.Y(n_6292)
);

BUFx2_ASAP7_75t_R g6293 ( 
.A(n_5914),
.Y(n_6293)
);

NOR2xp33_ASAP7_75t_L g6294 ( 
.A(n_5913),
.B(n_181),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_5964),
.Y(n_6295)
);

CKINVDCx5p33_ASAP7_75t_R g6296 ( 
.A(n_5824),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5898),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5912),
.Y(n_6298)
);

INVx6_ASAP7_75t_L g6299 ( 
.A(n_5811),
.Y(n_6299)
);

OAI21x1_ASAP7_75t_L g6300 ( 
.A1(n_5865),
.A2(n_182),
.B(n_183),
.Y(n_6300)
);

A2O1A1Ixp33_ASAP7_75t_L g6301 ( 
.A1(n_5992),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_6301)
);

NAND2xp5_ASAP7_75t_L g6302 ( 
.A(n_5953),
.B(n_5966),
.Y(n_6302)
);

OA21x2_ASAP7_75t_L g6303 ( 
.A1(n_6019),
.A2(n_185),
.B(n_187),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5969),
.Y(n_6304)
);

AND2x4_ASAP7_75t_L g6305 ( 
.A(n_5956),
.B(n_185),
.Y(n_6305)
);

AOI21xp5_ASAP7_75t_L g6306 ( 
.A1(n_5848),
.A2(n_187),
.B(n_188),
.Y(n_6306)
);

INVx4_ASAP7_75t_L g6307 ( 
.A(n_5822),
.Y(n_6307)
);

BUFx2_ASAP7_75t_L g6308 ( 
.A(n_5814),
.Y(n_6308)
);

BUFx10_ASAP7_75t_L g6309 ( 
.A(n_5913),
.Y(n_6309)
);

BUFx6f_ASAP7_75t_L g6310 ( 
.A(n_5822),
.Y(n_6310)
);

OAI21x1_ASAP7_75t_L g6311 ( 
.A1(n_5922),
.A2(n_189),
.B(n_190),
.Y(n_6311)
);

AOI21xp5_ASAP7_75t_L g6312 ( 
.A1(n_5848),
.A2(n_189),
.B(n_190),
.Y(n_6312)
);

OA21x2_ASAP7_75t_L g6313 ( 
.A1(n_6021),
.A2(n_191),
.B(n_192),
.Y(n_6313)
);

NAND2x1p5_ASAP7_75t_L g6314 ( 
.A(n_5936),
.B(n_3260),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_5964),
.Y(n_6315)
);

INVx4_ASAP7_75t_L g6316 ( 
.A(n_5913),
.Y(n_6316)
);

CKINVDCx11_ASAP7_75t_R g6317 ( 
.A(n_6001),
.Y(n_6317)
);

INVx4_ASAP7_75t_L g6318 ( 
.A(n_5936),
.Y(n_6318)
);

OAI21xp5_ASAP7_75t_L g6319 ( 
.A1(n_5961),
.A2(n_6071),
.B(n_5923),
.Y(n_6319)
);

NAND3xp33_ASAP7_75t_L g6320 ( 
.A(n_5961),
.B(n_193),
.C(n_194),
.Y(n_6320)
);

INVx3_ASAP7_75t_L g6321 ( 
.A(n_5944),
.Y(n_6321)
);

OAI21x1_ASAP7_75t_L g6322 ( 
.A1(n_5845),
.A2(n_193),
.B(n_194),
.Y(n_6322)
);

OAI21x1_ASAP7_75t_L g6323 ( 
.A1(n_5839),
.A2(n_196),
.B(n_197),
.Y(n_6323)
);

OA21x2_ASAP7_75t_L g6324 ( 
.A1(n_5949),
.A2(n_196),
.B(n_197),
.Y(n_6324)
);

OAI21x1_ASAP7_75t_L g6325 ( 
.A1(n_5949),
.A2(n_198),
.B(n_199),
.Y(n_6325)
);

OAI21x1_ASAP7_75t_L g6326 ( 
.A1(n_5978),
.A2(n_6048),
.B(n_5881),
.Y(n_6326)
);

OR2x2_ASAP7_75t_L g6327 ( 
.A(n_5814),
.B(n_201),
.Y(n_6327)
);

AND2x4_ASAP7_75t_L g6328 ( 
.A(n_5956),
.B(n_202),
.Y(n_6328)
);

AO31x2_ASAP7_75t_L g6329 ( 
.A1(n_6022),
.A2(n_205),
.A3(n_203),
.B(n_204),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_5969),
.Y(n_6330)
);

NAND2x1p5_ASAP7_75t_L g6331 ( 
.A(n_5973),
.B(n_3316),
.Y(n_6331)
);

OAI21x1_ASAP7_75t_L g6332 ( 
.A1(n_5978),
.A2(n_204),
.B(n_205),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_5944),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_6014),
.Y(n_6334)
);

AO21x1_ASAP7_75t_L g6335 ( 
.A1(n_6010),
.A2(n_206),
.B(n_207),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_5953),
.B(n_206),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_5858),
.Y(n_6337)
);

OA21x2_ASAP7_75t_L g6338 ( 
.A1(n_6078),
.A2(n_207),
.B(n_208),
.Y(n_6338)
);

OAI21xp5_ASAP7_75t_L g6339 ( 
.A1(n_6071),
.A2(n_208),
.B(n_209),
.Y(n_6339)
);

INVx2_ASAP7_75t_SL g6340 ( 
.A(n_5832),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6014),
.Y(n_6341)
);

OAI21x1_ASAP7_75t_L g6342 ( 
.A1(n_6048),
.A2(n_210),
.B(n_211),
.Y(n_6342)
);

OAI21x1_ASAP7_75t_L g6343 ( 
.A1(n_6055),
.A2(n_211),
.B(n_212),
.Y(n_6343)
);

NAND2x1p5_ASAP7_75t_L g6344 ( 
.A(n_5973),
.B(n_3316),
.Y(n_6344)
);

OR2x2_ASAP7_75t_L g6345 ( 
.A(n_5814),
.B(n_212),
.Y(n_6345)
);

INVx2_ASAP7_75t_L g6346 ( 
.A(n_5858),
.Y(n_6346)
);

NOR2xp33_ASAP7_75t_L g6347 ( 
.A(n_6209),
.B(n_5980),
.Y(n_6347)
);

AND2x4_ASAP7_75t_L g6348 ( 
.A(n_6288),
.B(n_5973),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_6134),
.Y(n_6349)
);

AOI21xp5_ASAP7_75t_L g6350 ( 
.A1(n_6109),
.A2(n_6063),
.B(n_5960),
.Y(n_6350)
);

OA21x2_ASAP7_75t_L g6351 ( 
.A1(n_6185),
.A2(n_6000),
.B(n_6078),
.Y(n_6351)
);

AND2x4_ASAP7_75t_L g6352 ( 
.A(n_6288),
.B(n_6318),
.Y(n_6352)
);

AND2x2_ASAP7_75t_L g6353 ( 
.A(n_6160),
.B(n_5872),
.Y(n_6353)
);

AND2x4_ASAP7_75t_L g6354 ( 
.A(n_6318),
.B(n_5973),
.Y(n_6354)
);

A2O1A1Ixp33_ASAP7_75t_L g6355 ( 
.A1(n_6319),
.A2(n_6222),
.B(n_6275),
.C(n_6117),
.Y(n_6355)
);

AOI21x1_ASAP7_75t_SL g6356 ( 
.A1(n_6271),
.A2(n_6001),
.B(n_6049),
.Y(n_6356)
);

NAND2xp5_ASAP7_75t_L g6357 ( 
.A(n_6100),
.B(n_6059),
.Y(n_6357)
);

AND2x2_ASAP7_75t_L g6358 ( 
.A(n_6160),
.B(n_6062),
.Y(n_6358)
);

AND2x4_ASAP7_75t_L g6359 ( 
.A(n_6316),
.B(n_6178),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6178),
.B(n_5972),
.Y(n_6360)
);

OR2x2_ASAP7_75t_L g6361 ( 
.A(n_6098),
.B(n_5807),
.Y(n_6361)
);

AOI21xp5_ASAP7_75t_SL g6362 ( 
.A1(n_6103),
.A2(n_6047),
.B(n_6063),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6333),
.B(n_6099),
.Y(n_6363)
);

AOI21xp5_ASAP7_75t_SL g6364 ( 
.A1(n_6103),
.A2(n_6007),
.B(n_6031),
.Y(n_6364)
);

AOI21xp5_ASAP7_75t_SL g6365 ( 
.A1(n_6225),
.A2(n_6031),
.B(n_5987),
.Y(n_6365)
);

AOI21xp5_ASAP7_75t_L g6366 ( 
.A1(n_6319),
.A2(n_5987),
.B(n_6089),
.Y(n_6366)
);

AOI21xp5_ASAP7_75t_SL g6367 ( 
.A1(n_6225),
.A2(n_6090),
.B(n_6089),
.Y(n_6367)
);

OAI22xp5_ASAP7_75t_L g6368 ( 
.A1(n_6320),
.A2(n_6082),
.B1(n_6005),
.B2(n_6054),
.Y(n_6368)
);

AND2x2_ASAP7_75t_L g6369 ( 
.A(n_6107),
.B(n_5972),
.Y(n_6369)
);

CKINVDCx9p33_ASAP7_75t_R g6370 ( 
.A(n_6127),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_6134),
.Y(n_6371)
);

AND2x2_ASAP7_75t_L g6372 ( 
.A(n_6128),
.B(n_6020),
.Y(n_6372)
);

NAND2xp5_ASAP7_75t_SL g6373 ( 
.A(n_6316),
.B(n_6092),
.Y(n_6373)
);

INVxp67_ASAP7_75t_L g6374 ( 
.A(n_6278),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_6095),
.Y(n_6375)
);

OAI22xp5_ASAP7_75t_L g6376 ( 
.A1(n_6320),
.A2(n_6082),
.B1(n_6005),
.B2(n_6054),
.Y(n_6376)
);

AOI221x1_ASAP7_75t_SL g6377 ( 
.A1(n_6258),
.A2(n_6091),
.B1(n_5925),
.B2(n_5938),
.C(n_6049),
.Y(n_6377)
);

AOI21xp5_ASAP7_75t_SL g6378 ( 
.A1(n_6324),
.A2(n_6090),
.B(n_6034),
.Y(n_6378)
);

AND2x2_ASAP7_75t_L g6379 ( 
.A(n_6135),
.B(n_6027),
.Y(n_6379)
);

OR2x2_ASAP7_75t_L g6380 ( 
.A(n_6124),
.B(n_5807),
.Y(n_6380)
);

NAND2xp5_ASAP7_75t_L g6381 ( 
.A(n_6100),
.B(n_6059),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_6308),
.B(n_6012),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6143),
.Y(n_6383)
);

O2A1O1Ixp5_ASAP7_75t_L g6384 ( 
.A1(n_6190),
.A2(n_5942),
.B(n_5888),
.C(n_5901),
.Y(n_6384)
);

A2O1A1Ixp33_ASAP7_75t_L g6385 ( 
.A1(n_6339),
.A2(n_5888),
.B(n_5901),
.C(n_5942),
.Y(n_6385)
);

INVx3_ASAP7_75t_L g6386 ( 
.A(n_6122),
.Y(n_6386)
);

A2O1A1Ixp33_ASAP7_75t_L g6387 ( 
.A1(n_6286),
.A2(n_5925),
.B(n_5835),
.C(n_6084),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_6095),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_L g6389 ( 
.A(n_6123),
.B(n_5970),
.Y(n_6389)
);

OAI22xp5_ASAP7_75t_L g6390 ( 
.A1(n_6258),
.A2(n_5980),
.B1(n_5843),
.B2(n_5835),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_6124),
.B(n_5970),
.Y(n_6391)
);

NAND2xp5_ASAP7_75t_L g6392 ( 
.A(n_6119),
.B(n_6041),
.Y(n_6392)
);

BUFx5_ASAP7_75t_L g6393 ( 
.A(n_6309),
.Y(n_6393)
);

NAND2xp5_ASAP7_75t_L g6394 ( 
.A(n_6119),
.B(n_6046),
.Y(n_6394)
);

A2O1A1Ixp33_ASAP7_75t_L g6395 ( 
.A1(n_6142),
.A2(n_6073),
.B(n_6030),
.C(n_6045),
.Y(n_6395)
);

O2A1O1Ixp5_ASAP7_75t_L g6396 ( 
.A1(n_6335),
.A2(n_5938),
.B(n_6032),
.C(n_6029),
.Y(n_6396)
);

NAND2x1p5_ASAP7_75t_L g6397 ( 
.A(n_6261),
.B(n_5994),
.Y(n_6397)
);

INVx2_ASAP7_75t_L g6398 ( 
.A(n_6321),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6143),
.Y(n_6399)
);

NAND2xp5_ASAP7_75t_L g6400 ( 
.A(n_6223),
.B(n_6092),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6337),
.B(n_6018),
.Y(n_6401)
);

AND2x2_ASAP7_75t_L g6402 ( 
.A(n_6346),
.B(n_5862),
.Y(n_6402)
);

INVxp67_ASAP7_75t_SL g6403 ( 
.A(n_6290),
.Y(n_6403)
);

OAI22xp5_ASAP7_75t_L g6404 ( 
.A1(n_6193),
.A2(n_5862),
.B1(n_6073),
.B2(n_5984),
.Y(n_6404)
);

OAI22xp5_ASAP7_75t_L g6405 ( 
.A1(n_6173),
.A2(n_5984),
.B1(n_5994),
.B2(n_6066),
.Y(n_6405)
);

AOI21x1_ASAP7_75t_SL g6406 ( 
.A1(n_6247),
.A2(n_6044),
.B(n_6035),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_6144),
.Y(n_6407)
);

OR2x2_ASAP7_75t_L g6408 ( 
.A(n_6263),
.B(n_6081),
.Y(n_6408)
);

BUFx12f_ASAP7_75t_L g6409 ( 
.A(n_6317),
.Y(n_6409)
);

AOI21xp5_ASAP7_75t_SL g6410 ( 
.A1(n_6324),
.A2(n_6034),
.B(n_6015),
.Y(n_6410)
);

NOR2xp67_ASAP7_75t_L g6411 ( 
.A(n_6307),
.B(n_6035),
.Y(n_6411)
);

INVx3_ASAP7_75t_SL g6412 ( 
.A(n_6296),
.Y(n_6412)
);

HB1xp67_ASAP7_75t_L g6413 ( 
.A(n_6334),
.Y(n_6413)
);

OAI22xp5_ASAP7_75t_L g6414 ( 
.A1(n_6301),
.A2(n_5984),
.B1(n_5879),
.B2(n_5899),
.Y(n_6414)
);

AOI21x1_ASAP7_75t_SL g6415 ( 
.A1(n_6305),
.A2(n_6328),
.B(n_6169),
.Y(n_6415)
);

OR2x2_ASAP7_75t_L g6416 ( 
.A(n_6101),
.B(n_5934),
.Y(n_6416)
);

OAI22xp5_ASAP7_75t_L g6417 ( 
.A1(n_6233),
.A2(n_6221),
.B1(n_6219),
.B2(n_6238),
.Y(n_6417)
);

HB1xp67_ASAP7_75t_L g6418 ( 
.A(n_6334),
.Y(n_6418)
);

AOI21xp5_ASAP7_75t_SL g6419 ( 
.A1(n_6280),
.A2(n_6052),
.B(n_6015),
.Y(n_6419)
);

OAI22xp5_ASAP7_75t_L g6420 ( 
.A1(n_6192),
.A2(n_6067),
.B1(n_6058),
.B2(n_6011),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_6144),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6146),
.Y(n_6422)
);

BUFx2_ASAP7_75t_L g6423 ( 
.A(n_6226),
.Y(n_6423)
);

AND2x4_ASAP7_75t_L g6424 ( 
.A(n_6305),
.B(n_6328),
.Y(n_6424)
);

NAND2xp5_ASAP7_75t_L g6425 ( 
.A(n_6175),
.B(n_6052),
.Y(n_6425)
);

AND2x2_ASAP7_75t_L g6426 ( 
.A(n_6120),
.B(n_6321),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_6248),
.Y(n_6427)
);

OA21x2_ASAP7_75t_L g6428 ( 
.A1(n_6283),
.A2(n_6044),
.B(n_6053),
.Y(n_6428)
);

NOR2xp67_ASAP7_75t_L g6429 ( 
.A(n_6307),
.B(n_6038),
.Y(n_6429)
);

OAI22xp5_ASAP7_75t_L g6430 ( 
.A1(n_6237),
.A2(n_6058),
.B1(n_6011),
.B2(n_5846),
.Y(n_6430)
);

NOR2xp67_ASAP7_75t_L g6431 ( 
.A(n_6341),
.B(n_6038),
.Y(n_6431)
);

NAND2xp5_ASAP7_75t_L g6432 ( 
.A(n_6341),
.B(n_5934),
.Y(n_6432)
);

OAI22xp5_ASAP7_75t_L g6433 ( 
.A1(n_6267),
.A2(n_6188),
.B1(n_6284),
.B2(n_6233),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6146),
.Y(n_6434)
);

OAI22xp5_ASAP7_75t_L g6435 ( 
.A1(n_6188),
.A2(n_6058),
.B1(n_6069),
.B2(n_5879),
.Y(n_6435)
);

AND2x2_ASAP7_75t_L g6436 ( 
.A(n_6309),
.B(n_6061),
.Y(n_6436)
);

OA21x2_ASAP7_75t_L g6437 ( 
.A1(n_6283),
.A2(n_5921),
.B(n_6076),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6106),
.B(n_6061),
.Y(n_6438)
);

HB1xp67_ASAP7_75t_L g6439 ( 
.A(n_6338),
.Y(n_6439)
);

OA21x2_ASAP7_75t_L g6440 ( 
.A1(n_6289),
.A2(n_5991),
.B(n_5989),
.Y(n_6440)
);

NAND2xp5_ASAP7_75t_L g6441 ( 
.A(n_6208),
.B(n_5919),
.Y(n_6441)
);

OR2x2_ASAP7_75t_L g6442 ( 
.A(n_6151),
.B(n_5919),
.Y(n_6442)
);

OA21x2_ASAP7_75t_L g6443 ( 
.A1(n_6289),
.A2(n_6072),
.B(n_6056),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_6125),
.B(n_5996),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_6254),
.Y(n_6445)
);

OAI22xp5_ASAP7_75t_L g6446 ( 
.A1(n_6235),
.A2(n_6069),
.B1(n_5954),
.B2(n_5852),
.Y(n_6446)
);

OAI22xp5_ASAP7_75t_L g6447 ( 
.A1(n_6156),
.A2(n_6069),
.B1(n_5954),
.B2(n_5852),
.Y(n_6447)
);

O2A1O1Ixp5_ASAP7_75t_L g6448 ( 
.A1(n_6165),
.A2(n_6306),
.B(n_6312),
.C(n_6257),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6153),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6153),
.Y(n_6450)
);

OR2x2_ASAP7_75t_L g6451 ( 
.A(n_6171),
.B(n_5996),
.Y(n_6451)
);

O2A1O1Ixp33_ASAP7_75t_L g6452 ( 
.A1(n_6229),
.A2(n_6074),
.B(n_6025),
.C(n_6079),
.Y(n_6452)
);

NAND2xp5_ASAP7_75t_L g6453 ( 
.A(n_6111),
.B(n_6006),
.Y(n_6453)
);

AND2x4_ASAP7_75t_L g6454 ( 
.A(n_6118),
.B(n_5954),
.Y(n_6454)
);

AOI21x1_ASAP7_75t_SL g6455 ( 
.A1(n_6166),
.A2(n_5896),
.B(n_5977),
.Y(n_6455)
);

OR2x2_ASAP7_75t_L g6456 ( 
.A(n_6132),
.B(n_6006),
.Y(n_6456)
);

HB1xp67_ASAP7_75t_L g6457 ( 
.A(n_6338),
.Y(n_6457)
);

OAI22xp5_ASAP7_75t_L g6458 ( 
.A1(n_6154),
.A2(n_6114),
.B1(n_6293),
.B2(n_6327),
.Y(n_6458)
);

OA21x2_ASAP7_75t_L g6459 ( 
.A1(n_6291),
.A2(n_5957),
.B(n_5883),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6158),
.Y(n_6460)
);

BUFx3_ASAP7_75t_L g6461 ( 
.A(n_6265),
.Y(n_6461)
);

AND2x2_ASAP7_75t_SL g6462 ( 
.A(n_6145),
.B(n_5833),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_6255),
.B(n_5889),
.Y(n_6463)
);

NOR2xp67_ASAP7_75t_L g6464 ( 
.A(n_6121),
.B(n_213),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_6295),
.B(n_5917),
.Y(n_6465)
);

AOI21x1_ASAP7_75t_SL g6466 ( 
.A1(n_6213),
.A2(n_6050),
.B(n_5907),
.Y(n_6466)
);

HB1xp67_ASAP7_75t_L g6467 ( 
.A(n_6132),
.Y(n_6467)
);

OAI22xp5_ASAP7_75t_L g6468 ( 
.A1(n_6345),
.A2(n_6206),
.B1(n_6299),
.B2(n_6191),
.Y(n_6468)
);

CKINVDCx20_ASAP7_75t_R g6469 ( 
.A(n_6139),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_6158),
.Y(n_6470)
);

NAND2xp5_ASAP7_75t_L g6471 ( 
.A(n_6336),
.B(n_5911),
.Y(n_6471)
);

HB1xp67_ASAP7_75t_L g6472 ( 
.A(n_6102),
.Y(n_6472)
);

AOI21xp5_ASAP7_75t_L g6473 ( 
.A1(n_6253),
.A2(n_6040),
.B(n_5976),
.Y(n_6473)
);

AND2x2_ASAP7_75t_L g6474 ( 
.A(n_6315),
.B(n_5882),
.Y(n_6474)
);

OR2x2_ASAP7_75t_L g6475 ( 
.A(n_6259),
.B(n_5988),
.Y(n_6475)
);

INVx2_ASAP7_75t_L g6476 ( 
.A(n_6310),
.Y(n_6476)
);

AND2x4_ASAP7_75t_L g6477 ( 
.A(n_6118),
.B(n_5981),
.Y(n_6477)
);

AOI21xp5_ASAP7_75t_SL g6478 ( 
.A1(n_6280),
.A2(n_213),
.B(n_214),
.Y(n_6478)
);

AOI21xp5_ASAP7_75t_L g6479 ( 
.A1(n_6201),
.A2(n_5983),
.B(n_6009),
.Y(n_6479)
);

OAI22xp5_ASAP7_75t_L g6480 ( 
.A1(n_6299),
.A2(n_5974),
.B1(n_5963),
.B2(n_6024),
.Y(n_6480)
);

NAND2xp5_ASAP7_75t_L g6481 ( 
.A(n_6302),
.B(n_6037),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6159),
.Y(n_6482)
);

OR2x2_ASAP7_75t_L g6483 ( 
.A(n_6259),
.B(n_214),
.Y(n_6483)
);

HB1xp67_ASAP7_75t_L g6484 ( 
.A(n_6102),
.Y(n_6484)
);

BUFx10_ASAP7_75t_L g6485 ( 
.A(n_6210),
.Y(n_6485)
);

OAI22xp5_ASAP7_75t_L g6486 ( 
.A1(n_6191),
.A2(n_6214),
.B1(n_6138),
.B2(n_6204),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_L g6487 ( 
.A(n_6126),
.B(n_6159),
.Y(n_6487)
);

AOI21x1_ASAP7_75t_SL g6488 ( 
.A1(n_6213),
.A2(n_215),
.B(n_216),
.Y(n_6488)
);

HB1xp67_ASAP7_75t_L g6489 ( 
.A(n_6104),
.Y(n_6489)
);

AND2x2_ASAP7_75t_L g6490 ( 
.A(n_6140),
.B(n_215),
.Y(n_6490)
);

NAND2xp5_ASAP7_75t_L g6491 ( 
.A(n_6126),
.B(n_6162),
.Y(n_6491)
);

INVxp67_ASAP7_75t_L g6492 ( 
.A(n_6310),
.Y(n_6492)
);

INVx2_ASAP7_75t_L g6493 ( 
.A(n_6310),
.Y(n_6493)
);

OR2x2_ASAP7_75t_L g6494 ( 
.A(n_6262),
.B(n_216),
.Y(n_6494)
);

OA21x2_ASAP7_75t_L g6495 ( 
.A1(n_6291),
.A2(n_6181),
.B(n_6304),
.Y(n_6495)
);

INVxp33_ASAP7_75t_SL g6496 ( 
.A(n_6276),
.Y(n_6496)
);

AOI21x1_ASAP7_75t_SL g6497 ( 
.A1(n_6194),
.A2(n_217),
.B(n_218),
.Y(n_6497)
);

CKINVDCx20_ASAP7_75t_R g6498 ( 
.A(n_6250),
.Y(n_6498)
);

INVxp33_ASAP7_75t_L g6499 ( 
.A(n_6164),
.Y(n_6499)
);

HB1xp67_ASAP7_75t_L g6500 ( 
.A(n_6104),
.Y(n_6500)
);

A2O1A1Ixp33_ASAP7_75t_L g6501 ( 
.A1(n_6245),
.A2(n_220),
.B(n_217),
.C(n_219),
.Y(n_6501)
);

INVxp67_ASAP7_75t_L g6502 ( 
.A(n_6266),
.Y(n_6502)
);

NAND2xp5_ASAP7_75t_L g6503 ( 
.A(n_6162),
.B(n_219),
.Y(n_6503)
);

OA21x2_ASAP7_75t_L g6504 ( 
.A1(n_6304),
.A2(n_222),
.B(n_223),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_6168),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_6168),
.B(n_6180),
.Y(n_6506)
);

HB1xp67_ASAP7_75t_L g6507 ( 
.A(n_6105),
.Y(n_6507)
);

OA21x2_ASAP7_75t_L g6508 ( 
.A1(n_6330),
.A2(n_223),
.B(n_224),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_L g6509 ( 
.A(n_6180),
.B(n_224),
.Y(n_6509)
);

O2A1O1Ixp5_ASAP7_75t_L g6510 ( 
.A1(n_6141),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_6510)
);

AND2x2_ASAP7_75t_L g6511 ( 
.A(n_6147),
.B(n_225),
.Y(n_6511)
);

AOI21xp5_ASAP7_75t_SL g6512 ( 
.A1(n_6211),
.A2(n_226),
.B(n_227),
.Y(n_6512)
);

AOI21xp5_ASAP7_75t_SL g6513 ( 
.A1(n_6211),
.A2(n_228),
.B(n_229),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_6183),
.Y(n_6514)
);

AOI21xp5_ASAP7_75t_L g6515 ( 
.A1(n_6217),
.A2(n_229),
.B(n_230),
.Y(n_6515)
);

CKINVDCx14_ASAP7_75t_R g6516 ( 
.A(n_6129),
.Y(n_6516)
);

HB1xp67_ASAP7_75t_L g6517 ( 
.A(n_6105),
.Y(n_6517)
);

INVx2_ASAP7_75t_L g6518 ( 
.A(n_6121),
.Y(n_6518)
);

NAND2xp5_ASAP7_75t_L g6519 ( 
.A(n_6183),
.B(n_230),
.Y(n_6519)
);

O2A1O1Ixp5_ASAP7_75t_L g6520 ( 
.A1(n_6155),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_6520)
);

NAND2xp5_ASAP7_75t_L g6521 ( 
.A(n_6216),
.B(n_231),
.Y(n_6521)
);

AOI21xp5_ASAP7_75t_L g6522 ( 
.A1(n_6217),
.A2(n_234),
.B(n_235),
.Y(n_6522)
);

OAI22xp5_ASAP7_75t_L g6523 ( 
.A1(n_6214),
.A2(n_3317),
.B1(n_3351),
.B2(n_3316),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6163),
.B(n_234),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_L g6525 ( 
.A(n_6216),
.B(n_6177),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_L g6526 ( 
.A(n_6177),
.B(n_235),
.Y(n_6526)
);

AND2x4_ASAP7_75t_L g6527 ( 
.A(n_6226),
.B(n_236),
.Y(n_6527)
);

NOR2xp67_ASAP7_75t_L g6528 ( 
.A(n_6137),
.B(n_6226),
.Y(n_6528)
);

OAI31xp33_ASAP7_75t_L g6529 ( 
.A1(n_6294),
.A2(n_239),
.A3(n_237),
.B(n_238),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6236),
.B(n_239),
.Y(n_6530)
);

O2A1O1Ixp5_ASAP7_75t_L g6531 ( 
.A1(n_6161),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_6531)
);

OAI22xp5_ASAP7_75t_L g6532 ( 
.A1(n_6340),
.A2(n_3317),
.B1(n_3351),
.B2(n_3316),
.Y(n_6532)
);

AND2x2_ASAP7_75t_L g6533 ( 
.A(n_6172),
.B(n_242),
.Y(n_6533)
);

BUFx3_ASAP7_75t_L g6534 ( 
.A(n_6179),
.Y(n_6534)
);

AND2x2_ASAP7_75t_L g6535 ( 
.A(n_6207),
.B(n_243),
.Y(n_6535)
);

OA21x2_ASAP7_75t_L g6536 ( 
.A1(n_6330),
.A2(n_244),
.B(n_246),
.Y(n_6536)
);

OAI31xp33_ASAP7_75t_L g6537 ( 
.A1(n_6279),
.A2(n_247),
.A3(n_244),
.B(n_246),
.Y(n_6537)
);

INVx2_ASAP7_75t_L g6538 ( 
.A(n_6137),
.Y(n_6538)
);

O2A1O1Ixp5_ASAP7_75t_L g6539 ( 
.A1(n_6227),
.A2(n_253),
.B(n_247),
.C(n_248),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_6203),
.B(n_254),
.Y(n_6540)
);

OAI22xp5_ASAP7_75t_L g6541 ( 
.A1(n_6303),
.A2(n_3317),
.B1(n_3351),
.B2(n_3316),
.Y(n_6541)
);

AND2x4_ASAP7_75t_L g6542 ( 
.A(n_6287),
.B(n_254),
.Y(n_6542)
);

OR2x2_ASAP7_75t_L g6543 ( 
.A(n_6262),
.B(n_255),
.Y(n_6543)
);

OA21x2_ASAP7_75t_L g6544 ( 
.A1(n_6251),
.A2(n_6115),
.B(n_6326),
.Y(n_6544)
);

HB1xp67_ASAP7_75t_L g6545 ( 
.A(n_6115),
.Y(n_6545)
);

OAI22xp5_ASAP7_75t_L g6546 ( 
.A1(n_6303),
.A2(n_3351),
.B1(n_3368),
.B2(n_3317),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6287),
.Y(n_6547)
);

OAI22xp5_ASAP7_75t_L g6548 ( 
.A1(n_6313),
.A2(n_3368),
.B1(n_3387),
.B2(n_3317),
.Y(n_6548)
);

AOI21xp5_ASAP7_75t_SL g6549 ( 
.A1(n_6281),
.A2(n_255),
.B(n_256),
.Y(n_6549)
);

AND2x2_ASAP7_75t_SL g6550 ( 
.A(n_6252),
.B(n_256),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6176),
.B(n_258),
.Y(n_6551)
);

BUFx2_ASAP7_75t_R g6552 ( 
.A(n_6240),
.Y(n_6552)
);

NOR2xp67_ASAP7_75t_L g6553 ( 
.A(n_6287),
.B(n_259),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6236),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_6274),
.B(n_260),
.Y(n_6555)
);

AND2x2_ASAP7_75t_L g6556 ( 
.A(n_6274),
.B(n_260),
.Y(n_6556)
);

AND2x2_ASAP7_75t_L g6557 ( 
.A(n_6256),
.B(n_261),
.Y(n_6557)
);

BUFx10_ASAP7_75t_L g6558 ( 
.A(n_6268),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6256),
.B(n_261),
.Y(n_6559)
);

AND2x4_ASAP7_75t_L g6560 ( 
.A(n_6198),
.B(n_262),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_6273),
.B(n_262),
.Y(n_6561)
);

AOI221x1_ASAP7_75t_SL g6562 ( 
.A1(n_6242),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_6562)
);

AOI21xp5_ASAP7_75t_L g6563 ( 
.A1(n_6186),
.A2(n_263),
.B(n_265),
.Y(n_6563)
);

A2O1A1Ixp33_ASAP7_75t_L g6564 ( 
.A1(n_6325),
.A2(n_6272),
.B(n_6200),
.C(n_6260),
.Y(n_6564)
);

AND2x2_ASAP7_75t_L g6565 ( 
.A(n_6273),
.B(n_268),
.Y(n_6565)
);

CKINVDCx5p33_ASAP7_75t_R g6566 ( 
.A(n_6231),
.Y(n_6566)
);

AOI221x1_ASAP7_75t_SL g6567 ( 
.A1(n_6242),
.A2(n_272),
.B1(n_268),
.B2(n_269),
.C(n_273),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_6220),
.B(n_272),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6269),
.Y(n_6569)
);

OA21x2_ASAP7_75t_L g6570 ( 
.A1(n_6277),
.A2(n_273),
.B(n_275),
.Y(n_6570)
);

AND2x2_ASAP7_75t_L g6571 ( 
.A(n_6297),
.B(n_6298),
.Y(n_6571)
);

OR2x2_ASAP7_75t_L g6572 ( 
.A(n_6269),
.B(n_276),
.Y(n_6572)
);

BUFx3_ASAP7_75t_L g6573 ( 
.A(n_6231),
.Y(n_6573)
);

NAND2xp5_ASAP7_75t_L g6574 ( 
.A(n_6232),
.B(n_277),
.Y(n_6574)
);

AOI21xp5_ASAP7_75t_SL g6575 ( 
.A1(n_6281),
.A2(n_279),
.B(n_280),
.Y(n_6575)
);

INVx1_ASAP7_75t_SL g6576 ( 
.A(n_6112),
.Y(n_6576)
);

OAI22xp5_ASAP7_75t_L g6577 ( 
.A1(n_6313),
.A2(n_3387),
.B1(n_3421),
.B2(n_3368),
.Y(n_6577)
);

AOI21xp5_ASAP7_75t_L g6578 ( 
.A1(n_6186),
.A2(n_282),
.B(n_283),
.Y(n_6578)
);

NAND2xp5_ASAP7_75t_L g6579 ( 
.A(n_6270),
.B(n_282),
.Y(n_6579)
);

OA21x2_ASAP7_75t_L g6580 ( 
.A1(n_6184),
.A2(n_284),
.B(n_285),
.Y(n_6580)
);

AND2x2_ASAP7_75t_L g6581 ( 
.A(n_6297),
.B(n_286),
.Y(n_6581)
);

INVx1_ASAP7_75t_SL g6582 ( 
.A(n_6112),
.Y(n_6582)
);

OAI22xp5_ASAP7_75t_L g6583 ( 
.A1(n_6282),
.A2(n_3387),
.B1(n_3421),
.B2(n_3368),
.Y(n_6583)
);

INVx1_ASAP7_75t_L g6584 ( 
.A(n_6270),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_6298),
.B(n_287),
.Y(n_6585)
);

O2A1O1Ixp33_ASAP7_75t_L g6586 ( 
.A1(n_6205),
.A2(n_290),
.B(n_288),
.C(n_289),
.Y(n_6586)
);

BUFx3_ASAP7_75t_L g6587 ( 
.A(n_6241),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6199),
.B(n_288),
.Y(n_6588)
);

HB1xp67_ASAP7_75t_L g6589 ( 
.A(n_6252),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_6292),
.Y(n_6590)
);

NOR2xp67_ASAP7_75t_L g6591 ( 
.A(n_6136),
.B(n_291),
.Y(n_6591)
);

OAI21xp5_ASAP7_75t_L g6592 ( 
.A1(n_6384),
.A2(n_6157),
.B(n_6110),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6413),
.Y(n_6593)
);

OR2x2_ASAP7_75t_L g6594 ( 
.A(n_6394),
.B(n_6170),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6418),
.Y(n_6595)
);

INVxp67_ASAP7_75t_L g6596 ( 
.A(n_6439),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6349),
.Y(n_6597)
);

BUFx3_ASAP7_75t_L g6598 ( 
.A(n_6573),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6371),
.Y(n_6599)
);

AND2x2_ASAP7_75t_L g6600 ( 
.A(n_6436),
.B(n_6189),
.Y(n_6600)
);

BUFx3_ASAP7_75t_L g6601 ( 
.A(n_6409),
.Y(n_6601)
);

BUFx2_ASAP7_75t_SL g6602 ( 
.A(n_6553),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6383),
.Y(n_6603)
);

INVx1_ASAP7_75t_SL g6604 ( 
.A(n_6370),
.Y(n_6604)
);

INVx3_ASAP7_75t_L g6605 ( 
.A(n_6348),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6399),
.Y(n_6606)
);

OA21x2_ASAP7_75t_L g6607 ( 
.A1(n_6366),
.A2(n_6108),
.B(n_6300),
.Y(n_6607)
);

OR2x2_ASAP7_75t_L g6608 ( 
.A(n_6403),
.B(n_6374),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6407),
.Y(n_6609)
);

AND2x2_ASAP7_75t_L g6610 ( 
.A(n_6353),
.B(n_6375),
.Y(n_6610)
);

INVx2_ASAP7_75t_L g6611 ( 
.A(n_6495),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6388),
.B(n_6198),
.Y(n_6612)
);

AND2x2_ASAP7_75t_L g6613 ( 
.A(n_6438),
.B(n_6218),
.Y(n_6613)
);

BUFx2_ASAP7_75t_L g6614 ( 
.A(n_6386),
.Y(n_6614)
);

AND2x2_ASAP7_75t_L g6615 ( 
.A(n_6424),
.B(n_6218),
.Y(n_6615)
);

OAI21x1_ASAP7_75t_L g6616 ( 
.A1(n_6415),
.A2(n_6150),
.B(n_6093),
.Y(n_6616)
);

BUFx6f_ASAP7_75t_L g6617 ( 
.A(n_6386),
.Y(n_6617)
);

INVx2_ASAP7_75t_L g6618 ( 
.A(n_6495),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_6424),
.B(n_6113),
.Y(n_6619)
);

HB1xp67_ASAP7_75t_L g6620 ( 
.A(n_6457),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6421),
.Y(n_6621)
);

OAI21x1_ASAP7_75t_L g6622 ( 
.A1(n_6406),
.A2(n_6131),
.B(n_6149),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_6422),
.Y(n_6623)
);

BUFx3_ASAP7_75t_L g6624 ( 
.A(n_6461),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6434),
.Y(n_6625)
);

OR2x2_ASAP7_75t_L g6626 ( 
.A(n_6425),
.B(n_6246),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6449),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6450),
.Y(n_6628)
);

OA21x2_ASAP7_75t_L g6629 ( 
.A1(n_6396),
.A2(n_6097),
.B(n_6212),
.Y(n_6629)
);

OR2x2_ASAP7_75t_L g6630 ( 
.A(n_6389),
.B(n_6246),
.Y(n_6630)
);

BUFx2_ASAP7_75t_L g6631 ( 
.A(n_6516),
.Y(n_6631)
);

BUFx3_ASAP7_75t_L g6632 ( 
.A(n_6566),
.Y(n_6632)
);

AND2x4_ASAP7_75t_L g6633 ( 
.A(n_6528),
.B(n_6187),
.Y(n_6633)
);

INVx2_ASAP7_75t_L g6634 ( 
.A(n_6560),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6460),
.Y(n_6635)
);

INVx5_ASAP7_75t_SL g6636 ( 
.A(n_6527),
.Y(n_6636)
);

OAI21x1_ASAP7_75t_L g6637 ( 
.A1(n_6351),
.A2(n_6130),
.B(n_6116),
.Y(n_6637)
);

OR2x2_ASAP7_75t_L g6638 ( 
.A(n_6357),
.B(n_6224),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6470),
.Y(n_6639)
);

CKINVDCx16_ASAP7_75t_R g6640 ( 
.A(n_6498),
.Y(n_6640)
);

INVx2_ASAP7_75t_L g6641 ( 
.A(n_6560),
.Y(n_6641)
);

HB1xp67_ASAP7_75t_L g6642 ( 
.A(n_6591),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6482),
.Y(n_6643)
);

HB1xp67_ASAP7_75t_L g6644 ( 
.A(n_6591),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_6505),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6514),
.Y(n_6646)
);

AND2x2_ASAP7_75t_L g6647 ( 
.A(n_6382),
.B(n_6268),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6554),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6472),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_6484),
.Y(n_6650)
);

AOI21xp33_ASAP7_75t_L g6651 ( 
.A1(n_6433),
.A2(n_6202),
.B(n_6230),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6489),
.Y(n_6652)
);

BUFx3_ASAP7_75t_L g6653 ( 
.A(n_6412),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6500),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6507),
.Y(n_6655)
);

INVx2_ASAP7_75t_L g6656 ( 
.A(n_6408),
.Y(n_6656)
);

AO21x2_ASAP7_75t_L g6657 ( 
.A1(n_6526),
.A2(n_6240),
.B(n_6228),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6398),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_6544),
.Y(n_6659)
);

OA21x2_ASAP7_75t_L g6660 ( 
.A1(n_6381),
.A2(n_6311),
.B(n_6215),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6359),
.B(n_6329),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_L g6662 ( 
.A(n_6377),
.B(n_6350),
.Y(n_6662)
);

NAND2x1p5_ASAP7_75t_L g6663 ( 
.A(n_6348),
.B(n_6285),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6517),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6359),
.B(n_6329),
.Y(n_6665)
);

BUFx6f_ASAP7_75t_L g6666 ( 
.A(n_6527),
.Y(n_6666)
);

BUFx2_ASAP7_75t_L g6667 ( 
.A(n_6423),
.Y(n_6667)
);

INVx2_ASAP7_75t_L g6668 ( 
.A(n_6544),
.Y(n_6668)
);

AND2x2_ASAP7_75t_L g6669 ( 
.A(n_6358),
.B(n_6329),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6504),
.Y(n_6670)
);

INVx2_ASAP7_75t_L g6671 ( 
.A(n_6504),
.Y(n_6671)
);

OA21x2_ASAP7_75t_L g6672 ( 
.A1(n_6448),
.A2(n_6355),
.B(n_6576),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6545),
.Y(n_6673)
);

INVx3_ASAP7_75t_L g6674 ( 
.A(n_6352),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6569),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_L g6676 ( 
.A(n_6377),
.B(n_6230),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6584),
.Y(n_6677)
);

INVx2_ASAP7_75t_L g6678 ( 
.A(n_6508),
.Y(n_6678)
);

INVx1_ASAP7_75t_SL g6679 ( 
.A(n_6496),
.Y(n_6679)
);

OAI21x1_ASAP7_75t_L g6680 ( 
.A1(n_6351),
.A2(n_6096),
.B(n_6167),
.Y(n_6680)
);

INVx3_ASAP7_75t_L g6681 ( 
.A(n_6352),
.Y(n_6681)
);

OR2x2_ASAP7_75t_L g6682 ( 
.A(n_6453),
.B(n_6224),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_6506),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6508),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_6536),
.Y(n_6685)
);

HB1xp67_ASAP7_75t_L g6686 ( 
.A(n_6589),
.Y(n_6686)
);

AND2x2_ASAP7_75t_L g6687 ( 
.A(n_6426),
.B(n_6187),
.Y(n_6687)
);

INVx3_ASAP7_75t_L g6688 ( 
.A(n_6354),
.Y(n_6688)
);

INVx2_ASAP7_75t_L g6689 ( 
.A(n_6536),
.Y(n_6689)
);

OR2x2_ASAP7_75t_L g6690 ( 
.A(n_6392),
.B(n_6224),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6571),
.Y(n_6691)
);

INVx2_ASAP7_75t_L g6692 ( 
.A(n_6363),
.Y(n_6692)
);

INVx2_ASAP7_75t_SL g6693 ( 
.A(n_6354),
.Y(n_6693)
);

INVx2_ASAP7_75t_L g6694 ( 
.A(n_6570),
.Y(n_6694)
);

INVx2_ASAP7_75t_L g6695 ( 
.A(n_6570),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6483),
.Y(n_6696)
);

OAI21x1_ASAP7_75t_L g6697 ( 
.A1(n_6525),
.A2(n_6344),
.B(n_6331),
.Y(n_6697)
);

HB1xp67_ASAP7_75t_L g6698 ( 
.A(n_6467),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6494),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6369),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6590),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_6543),
.Y(n_6702)
);

AND2x2_ASAP7_75t_L g6703 ( 
.A(n_6476),
.B(n_6314),
.Y(n_6703)
);

BUFx3_ASAP7_75t_L g6704 ( 
.A(n_6542),
.Y(n_6704)
);

INVx2_ASAP7_75t_L g6705 ( 
.A(n_6547),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6572),
.Y(n_6706)
);

AO21x2_ASAP7_75t_L g6707 ( 
.A1(n_6411),
.A2(n_6234),
.B(n_6323),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6487),
.Y(n_6708)
);

INVx3_ASAP7_75t_L g6709 ( 
.A(n_6454),
.Y(n_6709)
);

INVx2_ASAP7_75t_L g6710 ( 
.A(n_6427),
.Y(n_6710)
);

INVx2_ASAP7_75t_L g6711 ( 
.A(n_6445),
.Y(n_6711)
);

AOI22xp33_ASAP7_75t_L g6712 ( 
.A1(n_6368),
.A2(n_6182),
.B1(n_6152),
.B2(n_6197),
.Y(n_6712)
);

NAND2xp5_ASAP7_75t_L g6713 ( 
.A(n_6550),
.B(n_6243),
.Y(n_6713)
);

BUFx3_ASAP7_75t_L g6714 ( 
.A(n_6542),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6491),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6585),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_6555),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_6556),
.Y(n_6718)
);

AO21x1_ASAP7_75t_SL g6719 ( 
.A1(n_6400),
.A2(n_6243),
.B(n_6332),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6557),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_6372),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_6576),
.Y(n_6722)
);

BUFx8_ASAP7_75t_L g6723 ( 
.A(n_6534),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6559),
.Y(n_6724)
);

INVx2_ASAP7_75t_L g6725 ( 
.A(n_6582),
.Y(n_6725)
);

INVx2_ASAP7_75t_L g6726 ( 
.A(n_6582),
.Y(n_6726)
);

INVx3_ASAP7_75t_L g6727 ( 
.A(n_6454),
.Y(n_6727)
);

INVx3_ASAP7_75t_L g6728 ( 
.A(n_6397),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6561),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6380),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6565),
.Y(n_6731)
);

AND2x2_ASAP7_75t_L g6732 ( 
.A(n_6493),
.B(n_6249),
.Y(n_6732)
);

BUFx2_ASAP7_75t_L g6733 ( 
.A(n_6393),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6581),
.Y(n_6734)
);

INVx2_ASAP7_75t_L g6735 ( 
.A(n_6580),
.Y(n_6735)
);

INVx2_ASAP7_75t_L g6736 ( 
.A(n_6580),
.Y(n_6736)
);

INVx2_ASAP7_75t_L g6737 ( 
.A(n_6360),
.Y(n_6737)
);

INVx2_ASAP7_75t_L g6738 ( 
.A(n_6456),
.Y(n_6738)
);

CKINVDCx20_ASAP7_75t_R g6739 ( 
.A(n_6469),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6579),
.Y(n_6740)
);

INVx1_ASAP7_75t_L g6741 ( 
.A(n_6540),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6402),
.B(n_6244),
.Y(n_6742)
);

BUFx2_ASAP7_75t_L g6743 ( 
.A(n_6393),
.Y(n_6743)
);

INVx2_ASAP7_75t_L g6744 ( 
.A(n_6475),
.Y(n_6744)
);

INVx2_ASAP7_75t_L g6745 ( 
.A(n_6428),
.Y(n_6745)
);

INVx2_ASAP7_75t_L g6746 ( 
.A(n_6428),
.Y(n_6746)
);

OA21x2_ASAP7_75t_L g6747 ( 
.A1(n_6395),
.A2(n_6264),
.B(n_6322),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6518),
.Y(n_6748)
);

OR2x6_ASAP7_75t_L g6749 ( 
.A(n_6362),
.B(n_6342),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_6538),
.Y(n_6750)
);

OAI21xp5_ASAP7_75t_L g6751 ( 
.A1(n_6385),
.A2(n_6196),
.B(n_6182),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_6503),
.Y(n_6752)
);

INVx2_ASAP7_75t_L g6753 ( 
.A(n_6401),
.Y(n_6753)
);

INVx2_ASAP7_75t_SL g6754 ( 
.A(n_6393),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6393),
.Y(n_6755)
);

BUFx2_ASAP7_75t_L g6756 ( 
.A(n_6393),
.Y(n_6756)
);

AND2x2_ASAP7_75t_L g6757 ( 
.A(n_6492),
.B(n_6195),
.Y(n_6757)
);

NOR2xp33_ASAP7_75t_L g6758 ( 
.A(n_6499),
.B(n_6152),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_6509),
.Y(n_6759)
);

HB1xp67_ASAP7_75t_L g6760 ( 
.A(n_6552),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6519),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_6521),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6563),
.B(n_6243),
.Y(n_6763)
);

NOR2xp33_ASAP7_75t_L g6764 ( 
.A(n_6347),
.B(n_291),
.Y(n_6764)
);

BUFx2_ASAP7_75t_L g6765 ( 
.A(n_6587),
.Y(n_6765)
);

HB1xp67_ASAP7_75t_L g6766 ( 
.A(n_6411),
.Y(n_6766)
);

OA21x2_ASAP7_75t_L g6767 ( 
.A1(n_6391),
.A2(n_6239),
.B(n_6195),
.Y(n_6767)
);

INVx1_ASAP7_75t_L g6768 ( 
.A(n_6530),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6535),
.Y(n_6769)
);

HB1xp67_ASAP7_75t_L g6770 ( 
.A(n_6464),
.Y(n_6770)
);

INVx1_ASAP7_75t_L g6771 ( 
.A(n_6551),
.Y(n_6771)
);

INVx2_ASAP7_75t_L g6772 ( 
.A(n_6474),
.Y(n_6772)
);

AO21x2_ASAP7_75t_L g6773 ( 
.A1(n_6528),
.A2(n_6343),
.B(n_6094),
.Y(n_6773)
);

INVx2_ASAP7_75t_L g6774 ( 
.A(n_6558),
.Y(n_6774)
);

CKINVDCx6p67_ASAP7_75t_R g6775 ( 
.A(n_6485),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6490),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_6558),
.Y(n_6777)
);

INVx2_ASAP7_75t_L g6778 ( 
.A(n_6416),
.Y(n_6778)
);

BUFx3_ASAP7_75t_L g6779 ( 
.A(n_6485),
.Y(n_6779)
);

INVx2_ASAP7_75t_L g6780 ( 
.A(n_6465),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6379),
.B(n_6148),
.Y(n_6781)
);

INVx1_ASAP7_75t_SL g6782 ( 
.A(n_6462),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_6373),
.B(n_6148),
.Y(n_6783)
);

OR2x6_ASAP7_75t_L g6784 ( 
.A(n_6364),
.B(n_6174),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6511),
.Y(n_6785)
);

INVx1_ASAP7_75t_SL g6786 ( 
.A(n_6588),
.Y(n_6786)
);

CKINVDCx5p33_ASAP7_75t_R g6787 ( 
.A(n_6478),
.Y(n_6787)
);

INVx2_ASAP7_75t_SL g6788 ( 
.A(n_6524),
.Y(n_6788)
);

INVx2_ASAP7_75t_L g6789 ( 
.A(n_6361),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6533),
.Y(n_6790)
);

INVx2_ASAP7_75t_L g6791 ( 
.A(n_6459),
.Y(n_6791)
);

AOI21x1_ASAP7_75t_L g6792 ( 
.A1(n_6464),
.A2(n_6174),
.B(n_6094),
.Y(n_6792)
);

BUFx3_ASAP7_75t_L g6793 ( 
.A(n_6568),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6444),
.Y(n_6794)
);

INVxp67_ASAP7_75t_L g6795 ( 
.A(n_6367),
.Y(n_6795)
);

AO21x2_ASAP7_75t_L g6796 ( 
.A1(n_6432),
.A2(n_6094),
.B(n_6133),
.Y(n_6796)
);

BUFx6f_ASAP7_75t_L g6797 ( 
.A(n_6574),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6410),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6419),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6378),
.Y(n_6800)
);

BUFx2_ASAP7_75t_L g6801 ( 
.A(n_6502),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6451),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_6531),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6459),
.Y(n_6804)
);

OR2x6_ASAP7_75t_L g6805 ( 
.A(n_6512),
.B(n_6133),
.Y(n_6805)
);

INVx3_ASAP7_75t_L g6806 ( 
.A(n_6477),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6437),
.Y(n_6807)
);

INVx2_ASAP7_75t_L g6808 ( 
.A(n_6437),
.Y(n_6808)
);

INVx2_ASAP7_75t_L g6809 ( 
.A(n_6477),
.Y(n_6809)
);

INVx2_ASAP7_75t_SL g6810 ( 
.A(n_6486),
.Y(n_6810)
);

BUFx6f_ASAP7_75t_L g6811 ( 
.A(n_6443),
.Y(n_6811)
);

CKINVDCx14_ASAP7_75t_R g6812 ( 
.A(n_6417),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6520),
.Y(n_6813)
);

HB1xp67_ASAP7_75t_L g6814 ( 
.A(n_6431),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6442),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_6441),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6468),
.B(n_6133),
.Y(n_6817)
);

BUFx8_ASAP7_75t_L g6818 ( 
.A(n_6553),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_SL g6819 ( 
.A(n_6417),
.B(n_3387),
.Y(n_6819)
);

INVx2_ASAP7_75t_L g6820 ( 
.A(n_6443),
.Y(n_6820)
);

INVx2_ASAP7_75t_L g6821 ( 
.A(n_6440),
.Y(n_6821)
);

CKINVDCx11_ASAP7_75t_R g6822 ( 
.A(n_6601),
.Y(n_6822)
);

OA21x2_ASAP7_75t_L g6823 ( 
.A1(n_6662),
.A2(n_6578),
.B(n_6387),
.Y(n_6823)
);

NOR2xp33_ASAP7_75t_L g6824 ( 
.A(n_6601),
.B(n_6458),
.Y(n_6824)
);

OA21x2_ASAP7_75t_L g6825 ( 
.A1(n_6676),
.A2(n_6522),
.B(n_6515),
.Y(n_6825)
);

AND2x4_ASAP7_75t_L g6826 ( 
.A(n_6631),
.B(n_6564),
.Y(n_6826)
);

OA21x2_ASAP7_75t_L g6827 ( 
.A1(n_6795),
.A2(n_6510),
.B(n_6414),
.Y(n_6827)
);

OAI22xp5_ASAP7_75t_L g6828 ( 
.A1(n_6812),
.A2(n_6376),
.B1(n_6390),
.B2(n_6414),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6604),
.B(n_6404),
.Y(n_6829)
);

INVx2_ASAP7_75t_SL g6830 ( 
.A(n_6723),
.Y(n_6830)
);

NAND2xp33_ASAP7_75t_R g6831 ( 
.A(n_6672),
.B(n_6513),
.Y(n_6831)
);

OAI21xp5_ASAP7_75t_L g6832 ( 
.A1(n_6812),
.A2(n_6672),
.B(n_6751),
.Y(n_6832)
);

OA21x2_ASAP7_75t_L g6833 ( 
.A1(n_6795),
.A2(n_6431),
.B(n_6471),
.Y(n_6833)
);

OAI21xp5_ASAP7_75t_L g6834 ( 
.A1(n_6672),
.A2(n_6365),
.B(n_6549),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6614),
.B(n_6405),
.Y(n_6835)
);

AND2x2_ASAP7_75t_L g6836 ( 
.A(n_6765),
.B(n_6463),
.Y(n_6836)
);

AND2x2_ASAP7_75t_L g6837 ( 
.A(n_6704),
.B(n_6420),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6803),
.B(n_6452),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6704),
.B(n_6430),
.Y(n_6839)
);

NOR2xp33_ASAP7_75t_SL g6840 ( 
.A(n_6640),
.B(n_6537),
.Y(n_6840)
);

OR2x2_ASAP7_75t_L g6841 ( 
.A(n_6801),
.B(n_6446),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6714),
.B(n_6481),
.Y(n_6842)
);

NOR2xp33_ASAP7_75t_L g6843 ( 
.A(n_6632),
.B(n_6586),
.Y(n_6843)
);

AOI221xp5_ASAP7_75t_L g6844 ( 
.A1(n_6760),
.A2(n_6435),
.B1(n_6567),
.B2(n_6562),
.C(n_6446),
.Y(n_6844)
);

AND2x4_ASAP7_75t_L g6845 ( 
.A(n_6624),
.B(n_6501),
.Y(n_6845)
);

HB1xp67_ASAP7_75t_L g6846 ( 
.A(n_6770),
.Y(n_6846)
);

NAND4xp25_ASAP7_75t_L g6847 ( 
.A(n_6651),
.B(n_6567),
.C(n_6562),
.D(n_6529),
.Y(n_6847)
);

AND2x2_ASAP7_75t_L g6848 ( 
.A(n_6714),
.B(n_6429),
.Y(n_6848)
);

OAI211xp5_ASAP7_75t_L g6849 ( 
.A1(n_6760),
.A2(n_6575),
.B(n_6529),
.C(n_6537),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_6620),
.Y(n_6850)
);

AND2x2_ASAP7_75t_L g6851 ( 
.A(n_6667),
.B(n_6429),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_6775),
.B(n_6779),
.Y(n_6852)
);

CKINVDCx14_ASAP7_75t_R g6853 ( 
.A(n_6739),
.Y(n_6853)
);

NOR2xp33_ASAP7_75t_L g6854 ( 
.A(n_6632),
.B(n_6447),
.Y(n_6854)
);

OAI22xp5_ASAP7_75t_L g6855 ( 
.A1(n_6784),
.A2(n_6541),
.B1(n_6548),
.B2(n_6546),
.Y(n_6855)
);

AOI21xp5_ASAP7_75t_L g6856 ( 
.A1(n_6787),
.A2(n_6539),
.B(n_6473),
.Y(n_6856)
);

AND2x2_ASAP7_75t_L g6857 ( 
.A(n_6779),
.B(n_6577),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6813),
.B(n_6479),
.Y(n_6858)
);

AO32x2_ASAP7_75t_L g6859 ( 
.A1(n_6810),
.A2(n_6356),
.A3(n_6455),
.B1(n_6532),
.B2(n_6523),
.Y(n_6859)
);

OR2x6_ASAP7_75t_L g6860 ( 
.A(n_6602),
.B(n_6488),
.Y(n_6860)
);

AND2x4_ASAP7_75t_L g6861 ( 
.A(n_6624),
.B(n_6497),
.Y(n_6861)
);

INVx2_ASAP7_75t_SL g6862 ( 
.A(n_6723),
.Y(n_6862)
);

A2O1A1Ixp33_ASAP7_75t_SL g6863 ( 
.A1(n_6758),
.A2(n_6480),
.B(n_6466),
.C(n_6583),
.Y(n_6863)
);

AND2x4_ASAP7_75t_SL g6864 ( 
.A(n_6739),
.B(n_3387),
.Y(n_6864)
);

NAND2xp33_ASAP7_75t_R g6865 ( 
.A(n_6787),
.B(n_292),
.Y(n_6865)
);

NAND2xp5_ASAP7_75t_L g6866 ( 
.A(n_6634),
.B(n_6440),
.Y(n_6866)
);

OAI21xp5_ASAP7_75t_L g6867 ( 
.A1(n_6784),
.A2(n_292),
.B(n_293),
.Y(n_6867)
);

AND2x2_ASAP7_75t_L g6868 ( 
.A(n_6610),
.B(n_294),
.Y(n_6868)
);

AND2x4_ASAP7_75t_L g6869 ( 
.A(n_6598),
.B(n_6653),
.Y(n_6869)
);

O2A1O1Ixp33_ASAP7_75t_SL g6870 ( 
.A1(n_6713),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_6870)
);

AND2x4_ASAP7_75t_L g6871 ( 
.A(n_6598),
.B(n_297),
.Y(n_6871)
);

NOR2xp33_ASAP7_75t_L g6872 ( 
.A(n_6679),
.B(n_297),
.Y(n_6872)
);

CKINVDCx11_ASAP7_75t_R g6873 ( 
.A(n_6617),
.Y(n_6873)
);

NOR2x1_ASAP7_75t_L g6874 ( 
.A(n_6784),
.B(n_299),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6634),
.B(n_299),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6641),
.B(n_300),
.Y(n_6876)
);

AOI22xp5_ASAP7_75t_L g6877 ( 
.A1(n_6749),
.A2(n_304),
.B1(n_301),
.B2(n_303),
.Y(n_6877)
);

A2O1A1Ixp33_ASAP7_75t_L g6878 ( 
.A1(n_6799),
.A2(n_306),
.B(n_301),
.C(n_304),
.Y(n_6878)
);

NOR2x1_ASAP7_75t_SL g6879 ( 
.A(n_6707),
.B(n_307),
.Y(n_6879)
);

NAND2xp5_ASAP7_75t_L g6880 ( 
.A(n_6641),
.B(n_307),
.Y(n_6880)
);

AOI221xp5_ASAP7_75t_L g6881 ( 
.A1(n_6798),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.C(n_311),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6620),
.Y(n_6882)
);

NAND2xp5_ASAP7_75t_L g6883 ( 
.A(n_6786),
.B(n_309),
.Y(n_6883)
);

AND2x4_ASAP7_75t_L g6884 ( 
.A(n_6674),
.B(n_312),
.Y(n_6884)
);

AND2x4_ASAP7_75t_L g6885 ( 
.A(n_6674),
.B(n_312),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6617),
.B(n_313),
.Y(n_6886)
);

AND2x4_ASAP7_75t_L g6887 ( 
.A(n_6653),
.B(n_313),
.Y(n_6887)
);

OAI21xp5_ASAP7_75t_L g6888 ( 
.A1(n_6749),
.A2(n_314),
.B(n_315),
.Y(n_6888)
);

CKINVDCx11_ASAP7_75t_R g6889 ( 
.A(n_6617),
.Y(n_6889)
);

OAI22xp5_ASAP7_75t_L g6890 ( 
.A1(n_6805),
.A2(n_318),
.B1(n_314),
.B2(n_317),
.Y(n_6890)
);

NAND2xp5_ASAP7_75t_L g6891 ( 
.A(n_6788),
.B(n_319),
.Y(n_6891)
);

AO32x2_ASAP7_75t_L g6892 ( 
.A1(n_6693),
.A2(n_322),
.A3(n_320),
.B1(n_321),
.B2(n_324),
.Y(n_6892)
);

AND2x2_ASAP7_75t_L g6893 ( 
.A(n_6617),
.B(n_6681),
.Y(n_6893)
);

NAND2xp5_ASAP7_75t_L g6894 ( 
.A(n_6770),
.B(n_321),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6608),
.B(n_322),
.Y(n_6895)
);

AND2x2_ASAP7_75t_L g6896 ( 
.A(n_6681),
.B(n_324),
.Y(n_6896)
);

AOI21xp5_ASAP7_75t_L g6897 ( 
.A1(n_6819),
.A2(n_325),
.B(n_327),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6686),
.Y(n_6898)
);

AND2x2_ASAP7_75t_L g6899 ( 
.A(n_6687),
.B(n_327),
.Y(n_6899)
);

O2A1O1Ixp33_ASAP7_75t_L g6900 ( 
.A1(n_6749),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_6900)
);

OAI21xp5_ASAP7_75t_L g6901 ( 
.A1(n_6592),
.A2(n_328),
.B(n_329),
.Y(n_6901)
);

NAND3xp33_ASAP7_75t_L g6902 ( 
.A(n_6712),
.B(n_331),
.C(n_332),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6686),
.Y(n_6903)
);

AOI221xp5_ASAP7_75t_L g6904 ( 
.A1(n_6819),
.A2(n_334),
.B1(n_331),
.B2(n_333),
.C(n_336),
.Y(n_6904)
);

AO32x2_ASAP7_75t_L g6905 ( 
.A1(n_6754),
.A2(n_339),
.A3(n_336),
.B1(n_338),
.B2(n_344),
.Y(n_6905)
);

AOI22xp5_ASAP7_75t_L g6906 ( 
.A1(n_6805),
.A2(n_345),
.B1(n_338),
.B2(n_344),
.Y(n_6906)
);

NOR2x1_ASAP7_75t_SL g6907 ( 
.A(n_6707),
.B(n_345),
.Y(n_6907)
);

AND2x2_ASAP7_75t_L g6908 ( 
.A(n_6647),
.B(n_346),
.Y(n_6908)
);

AND2x2_ASAP7_75t_L g6909 ( 
.A(n_6600),
.B(n_346),
.Y(n_6909)
);

A2O1A1Ixp33_ASAP7_75t_L g6910 ( 
.A1(n_6800),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_6910)
);

AOI21xp5_ASAP7_75t_L g6911 ( 
.A1(n_6763),
.A2(n_6805),
.B(n_6782),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6698),
.Y(n_6912)
);

NAND2xp5_ASAP7_75t_L g6913 ( 
.A(n_6776),
.B(n_350),
.Y(n_6913)
);

AND2x4_ASAP7_75t_L g6914 ( 
.A(n_6666),
.B(n_6774),
.Y(n_6914)
);

NAND2xp5_ASAP7_75t_L g6915 ( 
.A(n_6785),
.B(n_352),
.Y(n_6915)
);

OAI22xp5_ASAP7_75t_L g6916 ( 
.A1(n_6712),
.A2(n_6596),
.B1(n_6747),
.B2(n_6671),
.Y(n_6916)
);

AND2x2_ASAP7_75t_L g6917 ( 
.A(n_6636),
.B(n_352),
.Y(n_6917)
);

OR2x2_ASAP7_75t_L g6918 ( 
.A(n_6656),
.B(n_353),
.Y(n_6918)
);

AND2x2_ASAP7_75t_L g6919 ( 
.A(n_6636),
.B(n_6703),
.Y(n_6919)
);

AND2x4_ASAP7_75t_L g6920 ( 
.A(n_6688),
.B(n_355),
.Y(n_6920)
);

OAI221xp5_ASAP7_75t_L g6921 ( 
.A1(n_6747),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.C(n_359),
.Y(n_6921)
);

OR2x2_ASAP7_75t_L g6922 ( 
.A(n_6656),
.B(n_357),
.Y(n_6922)
);

OR2x2_ASAP7_75t_L g6923 ( 
.A(n_6700),
.B(n_359),
.Y(n_6923)
);

OAI21xp5_ASAP7_75t_L g6924 ( 
.A1(n_6747),
.A2(n_360),
.B(n_361),
.Y(n_6924)
);

BUFx12f_ASAP7_75t_L g6925 ( 
.A(n_6818),
.Y(n_6925)
);

OR2x2_ASAP7_75t_L g6926 ( 
.A(n_6700),
.B(n_360),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6698),
.Y(n_6927)
);

AND2x4_ASAP7_75t_L g6928 ( 
.A(n_6688),
.B(n_362),
.Y(n_6928)
);

AO21x2_ASAP7_75t_L g6929 ( 
.A1(n_6596),
.A2(n_363),
.B(n_364),
.Y(n_6929)
);

OA21x2_ASAP7_75t_L g6930 ( 
.A1(n_6611),
.A2(n_364),
.B(n_365),
.Y(n_6930)
);

OR2x2_ASAP7_75t_L g6931 ( 
.A(n_6696),
.B(n_366),
.Y(n_6931)
);

AND2x2_ASAP7_75t_L g6932 ( 
.A(n_6636),
.B(n_367),
.Y(n_6932)
);

AO21x2_ASAP7_75t_L g6933 ( 
.A1(n_6684),
.A2(n_367),
.B(n_368),
.Y(n_6933)
);

OR2x2_ASAP7_75t_L g6934 ( 
.A(n_6699),
.B(n_371),
.Y(n_6934)
);

AOI22xp5_ASAP7_75t_L g6935 ( 
.A1(n_6774),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_6935)
);

INVx1_ASAP7_75t_L g6936 ( 
.A(n_6642),
.Y(n_6936)
);

AND2x4_ASAP7_75t_L g6937 ( 
.A(n_6666),
.B(n_374),
.Y(n_6937)
);

OAI21x1_ASAP7_75t_SL g6938 ( 
.A1(n_6792),
.A2(n_6671),
.B(n_6670),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6642),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_6753),
.B(n_375),
.Y(n_6940)
);

NOR2x1_ASAP7_75t_SL g6941 ( 
.A(n_6719),
.B(n_6657),
.Y(n_6941)
);

AO32x2_ASAP7_75t_L g6942 ( 
.A1(n_6657),
.A2(n_378),
.A3(n_376),
.B1(n_377),
.B2(n_379),
.Y(n_6942)
);

OR2x2_ASAP7_75t_L g6943 ( 
.A(n_6702),
.B(n_376),
.Y(n_6943)
);

AND2x4_ASAP7_75t_L g6944 ( 
.A(n_6605),
.B(n_378),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6753),
.B(n_379),
.Y(n_6945)
);

AOI22xp5_ASAP7_75t_L g6946 ( 
.A1(n_6777),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_6742),
.B(n_381),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6709),
.B(n_382),
.Y(n_6948)
);

AOI21xp5_ASAP7_75t_L g6949 ( 
.A1(n_6685),
.A2(n_383),
.B(n_384),
.Y(n_6949)
);

INVxp67_ASAP7_75t_L g6950 ( 
.A(n_6644),
.Y(n_6950)
);

OAI21xp5_ASAP7_75t_L g6951 ( 
.A1(n_6616),
.A2(n_385),
.B(n_386),
.Y(n_6951)
);

HB1xp67_ASAP7_75t_L g6952 ( 
.A(n_6644),
.Y(n_6952)
);

O2A1O1Ixp5_ASAP7_75t_L g6953 ( 
.A1(n_6670),
.A2(n_391),
.B(n_385),
.C(n_390),
.Y(n_6953)
);

INVxp67_ASAP7_75t_L g6954 ( 
.A(n_6666),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6709),
.B(n_391),
.Y(n_6955)
);

NOR2xp67_ASAP7_75t_L g6956 ( 
.A(n_6728),
.B(n_392),
.Y(n_6956)
);

AND2x2_ASAP7_75t_L g6957 ( 
.A(n_6727),
.B(n_393),
.Y(n_6957)
);

INVx4_ASAP7_75t_L g6958 ( 
.A(n_6666),
.Y(n_6958)
);

HB1xp67_ASAP7_75t_L g6959 ( 
.A(n_6766),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6593),
.Y(n_6960)
);

OR2x2_ASAP7_75t_L g6961 ( 
.A(n_6706),
.B(n_394),
.Y(n_6961)
);

AOI221xp5_ASAP7_75t_L g6962 ( 
.A1(n_6758),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.C(n_397),
.Y(n_6962)
);

INVx2_ASAP7_75t_L g6963 ( 
.A(n_6605),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6727),
.B(n_395),
.Y(n_6964)
);

INVx3_ASAP7_75t_L g6965 ( 
.A(n_6633),
.Y(n_6965)
);

AOI22xp5_ASAP7_75t_L g6966 ( 
.A1(n_6777),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_6966)
);

A2O1A1Ixp33_ASAP7_75t_L g6967 ( 
.A1(n_6764),
.A2(n_6689),
.B(n_6678),
.C(n_6622),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6612),
.B(n_399),
.Y(n_6968)
);

A2O1A1Ixp33_ASAP7_75t_L g6969 ( 
.A1(n_6764),
.A2(n_404),
.B(n_400),
.C(n_402),
.Y(n_6969)
);

OA21x2_ASAP7_75t_L g6970 ( 
.A1(n_6611),
.A2(n_400),
.B(n_404),
.Y(n_6970)
);

AND2x2_ASAP7_75t_L g6971 ( 
.A(n_6737),
.B(n_406),
.Y(n_6971)
);

AND2x4_ASAP7_75t_L g6972 ( 
.A(n_6790),
.B(n_407),
.Y(n_6972)
);

OA21x2_ASAP7_75t_L g6973 ( 
.A1(n_6618),
.A2(n_408),
.B(n_409),
.Y(n_6973)
);

OA21x2_ASAP7_75t_L g6974 ( 
.A1(n_6618),
.A2(n_408),
.B(n_409),
.Y(n_6974)
);

AND2x2_ASAP7_75t_L g6975 ( 
.A(n_6737),
.B(n_414),
.Y(n_6975)
);

AO21x2_ASAP7_75t_L g6976 ( 
.A1(n_6722),
.A2(n_415),
.B(n_416),
.Y(n_6976)
);

AND2x4_ASAP7_75t_L g6977 ( 
.A(n_6633),
.B(n_415),
.Y(n_6977)
);

AND2x4_ASAP7_75t_L g6978 ( 
.A(n_6633),
.B(n_416),
.Y(n_6978)
);

O2A1O1Ixp33_ASAP7_75t_L g6979 ( 
.A1(n_6678),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_6979)
);

AND2x2_ASAP7_75t_L g6980 ( 
.A(n_6721),
.B(n_417),
.Y(n_6980)
);

INVx1_ASAP7_75t_SL g6981 ( 
.A(n_6669),
.Y(n_6981)
);

NOR2xp33_ASAP7_75t_L g6982 ( 
.A(n_6797),
.B(n_419),
.Y(n_6982)
);

OR2x2_ASAP7_75t_L g6983 ( 
.A(n_6793),
.B(n_421),
.Y(n_6983)
);

AND2x2_ASAP7_75t_L g6984 ( 
.A(n_6721),
.B(n_421),
.Y(n_6984)
);

INVx4_ASAP7_75t_L g6985 ( 
.A(n_6797),
.Y(n_6985)
);

INVx2_ASAP7_75t_L g6986 ( 
.A(n_6806),
.Y(n_6986)
);

AO32x1_ASAP7_75t_L g6987 ( 
.A1(n_6689),
.A2(n_425),
.A3(n_422),
.B1(n_423),
.B2(n_427),
.Y(n_6987)
);

OR2x6_ASAP7_75t_L g6988 ( 
.A(n_6797),
.B(n_422),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_SL g6989 ( 
.A(n_6797),
.B(n_3421),
.Y(n_6989)
);

OR2x2_ASAP7_75t_L g6990 ( 
.A(n_6793),
.B(n_423),
.Y(n_6990)
);

NAND2xp5_ASAP7_75t_L g6991 ( 
.A(n_6717),
.B(n_425),
.Y(n_6991)
);

O2A1O1Ixp33_ASAP7_75t_L g6992 ( 
.A1(n_6694),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_6992)
);

OAI221xp5_ASAP7_75t_SL g6993 ( 
.A1(n_6638),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.C(n_431),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6718),
.B(n_430),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6595),
.Y(n_6995)
);

HB1xp67_ASAP7_75t_L g6996 ( 
.A(n_6766),
.Y(n_6996)
);

NOR2xp33_ASAP7_75t_L g6997 ( 
.A(n_6818),
.B(n_431),
.Y(n_6997)
);

AND2x2_ASAP7_75t_L g6998 ( 
.A(n_6757),
.B(n_432),
.Y(n_6998)
);

O2A1O1Ixp33_ASAP7_75t_SL g6999 ( 
.A1(n_6690),
.A2(n_435),
.B(n_433),
.C(n_434),
.Y(n_6999)
);

OA21x2_ASAP7_75t_L g7000 ( 
.A1(n_6659),
.A2(n_437),
.B(n_438),
.Y(n_7000)
);

AND2x4_ASAP7_75t_L g7001 ( 
.A(n_6771),
.B(n_437),
.Y(n_7001)
);

OAI22xp5_ASAP7_75t_L g7002 ( 
.A1(n_6694),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_SL g7003 ( 
.A(n_6728),
.B(n_3421),
.Y(n_7003)
);

AO21x2_ASAP7_75t_L g7004 ( 
.A1(n_6722),
.A2(n_439),
.B(n_440),
.Y(n_7004)
);

HB1xp67_ASAP7_75t_L g7005 ( 
.A(n_6952),
.Y(n_7005)
);

HB1xp67_ASAP7_75t_L g7006 ( 
.A(n_6846),
.Y(n_7006)
);

BUFx2_ASAP7_75t_L g7007 ( 
.A(n_6853),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6936),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_6954),
.B(n_6720),
.Y(n_7009)
);

AND2x2_ASAP7_75t_L g7010 ( 
.A(n_6869),
.B(n_6852),
.Y(n_7010)
);

NOR2x1_ASAP7_75t_L g7011 ( 
.A(n_6874),
.B(n_6725),
.Y(n_7011)
);

BUFx2_ASAP7_75t_L g7012 ( 
.A(n_6925),
.Y(n_7012)
);

AOI22xp33_ASAP7_75t_SL g7013 ( 
.A1(n_6840),
.A2(n_6817),
.B1(n_6695),
.B2(n_6736),
.Y(n_7013)
);

HB1xp67_ASAP7_75t_L g7014 ( 
.A(n_6959),
.Y(n_7014)
);

INVx2_ASAP7_75t_SL g7015 ( 
.A(n_6830),
.Y(n_7015)
);

HB1xp67_ASAP7_75t_L g7016 ( 
.A(n_6996),
.Y(n_7016)
);

INVx2_ASAP7_75t_L g7017 ( 
.A(n_6941),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6939),
.Y(n_7018)
);

INVx2_ASAP7_75t_L g7019 ( 
.A(n_6958),
.Y(n_7019)
);

AND2x2_ASAP7_75t_L g7020 ( 
.A(n_6919),
.B(n_6732),
.Y(n_7020)
);

OAI221xp5_ASAP7_75t_L g7021 ( 
.A1(n_6834),
.A2(n_6695),
.B1(n_6736),
.B2(n_6735),
.C(n_6682),
.Y(n_7021)
);

AND2x2_ASAP7_75t_L g7022 ( 
.A(n_6893),
.B(n_6724),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6862),
.B(n_6729),
.Y(n_7023)
);

INVx2_ASAP7_75t_L g7024 ( 
.A(n_6965),
.Y(n_7024)
);

INVx4_ASAP7_75t_L g7025 ( 
.A(n_6822),
.Y(n_7025)
);

INVx2_ASAP7_75t_SL g7026 ( 
.A(n_6977),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6879),
.Y(n_7027)
);

OR2x2_ASAP7_75t_L g7028 ( 
.A(n_6838),
.B(n_6981),
.Y(n_7028)
);

NAND2xp5_ASAP7_75t_L g7029 ( 
.A(n_6914),
.B(n_6731),
.Y(n_7029)
);

INVx2_ASAP7_75t_L g7030 ( 
.A(n_6907),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6850),
.Y(n_7031)
);

HB1xp67_ASAP7_75t_L g7032 ( 
.A(n_6831),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6882),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6826),
.B(n_6839),
.Y(n_7034)
);

HB1xp67_ASAP7_75t_L g7035 ( 
.A(n_6930),
.Y(n_7035)
);

AND2x2_ASAP7_75t_L g7036 ( 
.A(n_6826),
.B(n_6837),
.Y(n_7036)
);

INVx1_ASAP7_75t_L g7037 ( 
.A(n_6898),
.Y(n_7037)
);

INVxp67_ASAP7_75t_SL g7038 ( 
.A(n_6865),
.Y(n_7038)
);

OR2x2_ASAP7_75t_L g7039 ( 
.A(n_6841),
.B(n_6692),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_L g7040 ( 
.A(n_6956),
.B(n_6734),
.Y(n_7040)
);

AND2x2_ASAP7_75t_L g7041 ( 
.A(n_6835),
.B(n_6619),
.Y(n_7041)
);

NAND2xp5_ASAP7_75t_L g7042 ( 
.A(n_6977),
.B(n_6741),
.Y(n_7042)
);

AND2x2_ASAP7_75t_L g7043 ( 
.A(n_6829),
.B(n_6661),
.Y(n_7043)
);

OR2x2_ASAP7_75t_L g7044 ( 
.A(n_6950),
.B(n_6692),
.Y(n_7044)
);

OR2x2_ASAP7_75t_L g7045 ( 
.A(n_6858),
.B(n_6963),
.Y(n_7045)
);

HB1xp67_ASAP7_75t_L g7046 ( 
.A(n_6930),
.Y(n_7046)
);

AND2x2_ASAP7_75t_L g7047 ( 
.A(n_6845),
.B(n_6665),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_6933),
.Y(n_7048)
);

AND2x2_ASAP7_75t_L g7049 ( 
.A(n_6861),
.B(n_6769),
.Y(n_7049)
);

OR2x2_ASAP7_75t_L g7050 ( 
.A(n_6895),
.B(n_6705),
.Y(n_7050)
);

INVx2_ASAP7_75t_L g7051 ( 
.A(n_6942),
.Y(n_7051)
);

AOI22xp33_ASAP7_75t_SL g7052 ( 
.A1(n_6828),
.A2(n_6735),
.B1(n_6615),
.B2(n_6607),
.Y(n_7052)
);

INVx2_ASAP7_75t_L g7053 ( 
.A(n_6873),
.Y(n_7053)
);

INVx2_ASAP7_75t_L g7054 ( 
.A(n_6942),
.Y(n_7054)
);

AND2x2_ASAP7_75t_L g7055 ( 
.A(n_6824),
.B(n_6705),
.Y(n_7055)
);

CKINVDCx5p33_ASAP7_75t_R g7056 ( 
.A(n_6889),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_L g7057 ( 
.A(n_6978),
.B(n_6740),
.Y(n_7057)
);

HB1xp67_ASAP7_75t_L g7058 ( 
.A(n_6970),
.Y(n_7058)
);

AND2x2_ASAP7_75t_L g7059 ( 
.A(n_6909),
.B(n_6716),
.Y(n_7059)
);

HB1xp67_ASAP7_75t_L g7060 ( 
.A(n_6970),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6903),
.Y(n_7061)
);

OAI22xp5_ASAP7_75t_L g7062 ( 
.A1(n_6844),
.A2(n_6663),
.B1(n_6726),
.B2(n_6725),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6912),
.Y(n_7063)
);

AND2x2_ASAP7_75t_L g7064 ( 
.A(n_6947),
.B(n_6752),
.Y(n_7064)
);

NAND2xp5_ASAP7_75t_L g7065 ( 
.A(n_6978),
.B(n_6759),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_6842),
.B(n_6761),
.Y(n_7066)
);

AND2x2_ASAP7_75t_L g7067 ( 
.A(n_6836),
.B(n_6762),
.Y(n_7067)
);

AND2x4_ASAP7_75t_L g7068 ( 
.A(n_6985),
.B(n_6649),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6942),
.Y(n_7069)
);

NAND2xp5_ASAP7_75t_L g7070 ( 
.A(n_6823),
.B(n_6768),
.Y(n_7070)
);

AND2x4_ASAP7_75t_L g7071 ( 
.A(n_6986),
.B(n_6650),
.Y(n_7071)
);

NOR2xp67_ASAP7_75t_L g7072 ( 
.A(n_6849),
.B(n_6814),
.Y(n_7072)
);

NAND2xp5_ASAP7_75t_SL g7073 ( 
.A(n_6832),
.B(n_6663),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6927),
.Y(n_7074)
);

AOI221xp5_ASAP7_75t_L g7075 ( 
.A1(n_6847),
.A2(n_6916),
.B1(n_6924),
.B2(n_6902),
.C(n_6921),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_6823),
.B(n_6652),
.Y(n_7076)
);

INVxp67_ASAP7_75t_SL g7077 ( 
.A(n_6900),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6980),
.Y(n_7078)
);

AND2x2_ASAP7_75t_L g7079 ( 
.A(n_6998),
.B(n_6613),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6984),
.Y(n_7080)
);

AND2x2_ASAP7_75t_L g7081 ( 
.A(n_6968),
.B(n_6691),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6911),
.B(n_6654),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6929),
.Y(n_7083)
);

OR2x2_ASAP7_75t_L g7084 ( 
.A(n_6880),
.B(n_6655),
.Y(n_7084)
);

INVx2_ASAP7_75t_L g7085 ( 
.A(n_6938),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6877),
.B(n_6664),
.Y(n_7086)
);

AOI221xp5_ASAP7_75t_L g7087 ( 
.A1(n_6856),
.A2(n_6794),
.B1(n_6726),
.B2(n_6673),
.C(n_6738),
.Y(n_7087)
);

BUFx2_ASAP7_75t_L g7088 ( 
.A(n_6988),
.Y(n_7088)
);

HB1xp67_ASAP7_75t_L g7089 ( 
.A(n_6973),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_6988),
.Y(n_7090)
);

AND2x4_ASAP7_75t_L g7091 ( 
.A(n_6848),
.B(n_6733),
.Y(n_7091)
);

OR2x2_ASAP7_75t_L g7092 ( 
.A(n_6918),
.B(n_6658),
.Y(n_7092)
);

INVx2_ASAP7_75t_L g7093 ( 
.A(n_6851),
.Y(n_7093)
);

AOI22xp5_ASAP7_75t_L g7094 ( 
.A1(n_6827),
.A2(n_6658),
.B1(n_6816),
.B2(n_6607),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6973),
.Y(n_7095)
);

INVx2_ASAP7_75t_L g7096 ( 
.A(n_6974),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6940),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6945),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6971),
.Y(n_7099)
);

AND2x2_ASAP7_75t_L g7100 ( 
.A(n_6899),
.B(n_6748),
.Y(n_7100)
);

INVx2_ASAP7_75t_L g7101 ( 
.A(n_6974),
.Y(n_7101)
);

INVxp67_ASAP7_75t_L g7102 ( 
.A(n_6976),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6857),
.B(n_6748),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_6975),
.Y(n_7104)
);

BUFx6f_ASAP7_75t_L g7105 ( 
.A(n_6905),
.Y(n_7105)
);

INVx2_ASAP7_75t_L g7106 ( 
.A(n_7000),
.Y(n_7106)
);

AND2x2_ASAP7_75t_L g7107 ( 
.A(n_6908),
.B(n_6750),
.Y(n_7107)
);

OAI211xp5_ASAP7_75t_L g7108 ( 
.A1(n_6888),
.A2(n_6967),
.B(n_6906),
.C(n_6867),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6922),
.Y(n_7109)
);

OR2x2_ASAP7_75t_L g7110 ( 
.A(n_6894),
.B(n_6594),
.Y(n_7110)
);

INVx3_ASAP7_75t_L g7111 ( 
.A(n_6944),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_6868),
.B(n_6750),
.Y(n_7112)
);

AND2x2_ASAP7_75t_L g7113 ( 
.A(n_6854),
.B(n_6710),
.Y(n_7113)
);

AND2x2_ASAP7_75t_L g7114 ( 
.A(n_6843),
.B(n_6710),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6875),
.Y(n_7115)
);

AOI221xp5_ASAP7_75t_L g7116 ( 
.A1(n_6962),
.A2(n_6993),
.B1(n_6890),
.B2(n_6979),
.C(n_6992),
.Y(n_7116)
);

AND2x2_ASAP7_75t_L g7117 ( 
.A(n_6896),
.B(n_6711),
.Y(n_7117)
);

HB1xp67_ASAP7_75t_L g7118 ( 
.A(n_7000),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_6944),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_6876),
.Y(n_7120)
);

AND2x4_ASAP7_75t_L g7121 ( 
.A(n_6884),
.B(n_6885),
.Y(n_7121)
);

AND2x4_ASAP7_75t_L g7122 ( 
.A(n_6884),
.B(n_6743),
.Y(n_7122)
);

INVx2_ASAP7_75t_L g7123 ( 
.A(n_6885),
.Y(n_7123)
);

INVx3_ASAP7_75t_L g7124 ( 
.A(n_6920),
.Y(n_7124)
);

BUFx2_ASAP7_75t_L g7125 ( 
.A(n_6920),
.Y(n_7125)
);

OR2x2_ASAP7_75t_L g7126 ( 
.A(n_6960),
.B(n_6711),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6948),
.B(n_6756),
.Y(n_7127)
);

INVxp67_ASAP7_75t_R g7128 ( 
.A(n_6917),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6923),
.Y(n_7129)
);

AND2x2_ASAP7_75t_L g7130 ( 
.A(n_6955),
.B(n_6809),
.Y(n_7130)
);

INVx2_ASAP7_75t_SL g7131 ( 
.A(n_6928),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6926),
.Y(n_7132)
);

BUFx3_ASAP7_75t_L g7133 ( 
.A(n_6928),
.Y(n_7133)
);

INVx2_ASAP7_75t_L g7134 ( 
.A(n_7004),
.Y(n_7134)
);

INVx2_ASAP7_75t_L g7135 ( 
.A(n_6833),
.Y(n_7135)
);

AND2x2_ASAP7_75t_L g7136 ( 
.A(n_6957),
.B(n_6809),
.Y(n_7136)
);

HB1xp67_ASAP7_75t_L g7137 ( 
.A(n_6825),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6931),
.Y(n_7138)
);

AO21x2_ASAP7_75t_L g7139 ( 
.A1(n_6863),
.A2(n_6668),
.B(n_6659),
.Y(n_7139)
);

AND2x4_ASAP7_75t_L g7140 ( 
.A(n_6964),
.B(n_6701),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6934),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6833),
.Y(n_7142)
);

AOI22xp33_ASAP7_75t_L g7143 ( 
.A1(n_6825),
.A2(n_6607),
.B1(n_6660),
.B2(n_6773),
.Y(n_7143)
);

HB1xp67_ASAP7_75t_L g7144 ( 
.A(n_6827),
.Y(n_7144)
);

INVx2_ASAP7_75t_SL g7145 ( 
.A(n_6871),
.Y(n_7145)
);

NAND2xp5_ASAP7_75t_L g7146 ( 
.A(n_6949),
.B(n_6683),
.Y(n_7146)
);

AND2x2_ASAP7_75t_L g7147 ( 
.A(n_6932),
.B(n_6802),
.Y(n_7147)
);

OR2x2_ASAP7_75t_L g7148 ( 
.A(n_7038),
.B(n_6995),
.Y(n_7148)
);

AND2x2_ASAP7_75t_L g7149 ( 
.A(n_7007),
.B(n_6886),
.Y(n_7149)
);

AND4x1_ASAP7_75t_L g7150 ( 
.A(n_7011),
.B(n_6881),
.C(n_6953),
.D(n_6901),
.Y(n_7150)
);

AOI22xp33_ASAP7_75t_L g7151 ( 
.A1(n_7075),
.A2(n_6951),
.B1(n_6630),
.B2(n_6783),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_L g7152 ( 
.A(n_7144),
.B(n_6982),
.Y(n_7152)
);

AND2x2_ASAP7_75t_L g7153 ( 
.A(n_7025),
.B(n_6872),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_SL g7154 ( 
.A(n_7121),
.B(n_6897),
.Y(n_7154)
);

NAND3xp33_ASAP7_75t_SL g7155 ( 
.A(n_7013),
.B(n_6904),
.C(n_6969),
.Y(n_7155)
);

NAND2xp5_ASAP7_75t_L g7156 ( 
.A(n_7144),
.B(n_6983),
.Y(n_7156)
);

AND2x2_ASAP7_75t_L g7157 ( 
.A(n_7025),
.B(n_6997),
.Y(n_7157)
);

NOR2xp33_ASAP7_75t_L g7158 ( 
.A(n_7038),
.B(n_6990),
.Y(n_7158)
);

OAI22xp5_ASAP7_75t_L g7159 ( 
.A1(n_7013),
.A2(n_6860),
.B1(n_6910),
.B2(n_6878),
.Y(n_7159)
);

NAND2xp5_ASAP7_75t_L g7160 ( 
.A(n_7032),
.B(n_6999),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_7032),
.B(n_7072),
.Y(n_7161)
);

NAND2xp5_ASAP7_75t_L g7162 ( 
.A(n_7026),
.B(n_6937),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_7125),
.B(n_6870),
.Y(n_7163)
);

AND2x2_ASAP7_75t_L g7164 ( 
.A(n_7012),
.B(n_6859),
.Y(n_7164)
);

OAI21xp5_ASAP7_75t_SL g7165 ( 
.A1(n_7108),
.A2(n_6946),
.B(n_6935),
.Y(n_7165)
);

NOR3xp33_ASAP7_75t_L g7166 ( 
.A(n_7075),
.B(n_6915),
.C(n_6913),
.Y(n_7166)
);

NAND3xp33_ASAP7_75t_L g7167 ( 
.A(n_7087),
.B(n_6966),
.C(n_7002),
.Y(n_7167)
);

NAND3xp33_ASAP7_75t_L g7168 ( 
.A(n_7087),
.B(n_6715),
.C(n_6708),
.Y(n_7168)
);

NAND2xp5_ASAP7_75t_L g7169 ( 
.A(n_7131),
.B(n_6991),
.Y(n_7169)
);

AOI221x1_ASAP7_75t_SL g7170 ( 
.A1(n_7062),
.A2(n_6866),
.B1(n_6994),
.B2(n_6855),
.C(n_6701),
.Y(n_7170)
);

OAI21xp33_ASAP7_75t_L g7171 ( 
.A1(n_7052),
.A2(n_6860),
.B(n_6781),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_L g7172 ( 
.A(n_7111),
.B(n_6943),
.Y(n_7172)
);

AND2x2_ASAP7_75t_L g7173 ( 
.A(n_7128),
.B(n_6859),
.Y(n_7173)
);

OAI221xp5_ASAP7_75t_SL g7174 ( 
.A1(n_7108),
.A2(n_6626),
.B1(n_6738),
.B2(n_6859),
.C(n_6668),
.Y(n_7174)
);

NAND2xp5_ASAP7_75t_L g7175 ( 
.A(n_7111),
.B(n_6961),
.Y(n_7175)
);

OAI21xp5_ASAP7_75t_SL g7176 ( 
.A1(n_7052),
.A2(n_6883),
.B(n_6891),
.Y(n_7176)
);

NAND3xp33_ASAP7_75t_L g7177 ( 
.A(n_7137),
.B(n_6811),
.C(n_6814),
.Y(n_7177)
);

NOR3xp33_ASAP7_75t_L g7178 ( 
.A(n_7021),
.B(n_6755),
.C(n_6972),
.Y(n_7178)
);

OAI221xp5_ASAP7_75t_SL g7179 ( 
.A1(n_7143),
.A2(n_6730),
.B1(n_6778),
.B2(n_6815),
.C(n_6745),
.Y(n_7179)
);

AND2x2_ASAP7_75t_L g7180 ( 
.A(n_7010),
.B(n_7001),
.Y(n_7180)
);

NAND2xp5_ASAP7_75t_L g7181 ( 
.A(n_7124),
.B(n_6887),
.Y(n_7181)
);

AND2x2_ASAP7_75t_L g7182 ( 
.A(n_7034),
.B(n_6755),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_7124),
.B(n_6597),
.Y(n_7183)
);

NAND3xp33_ASAP7_75t_L g7184 ( 
.A(n_7137),
.B(n_6811),
.C(n_6989),
.Y(n_7184)
);

NOR3xp33_ASAP7_75t_SL g7185 ( 
.A(n_7056),
.B(n_7003),
.C(n_6603),
.Y(n_7185)
);

NAND2xp5_ASAP7_75t_L g7186 ( 
.A(n_7077),
.B(n_7027),
.Y(n_7186)
);

OAI22xp5_ASAP7_75t_L g7187 ( 
.A1(n_7105),
.A2(n_6629),
.B1(n_6811),
.B2(n_6660),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_L g7188 ( 
.A(n_7077),
.B(n_6599),
.Y(n_7188)
);

OAI21xp33_ASAP7_75t_SL g7189 ( 
.A1(n_7143),
.A2(n_6616),
.B(n_6680),
.Y(n_7189)
);

NAND3xp33_ASAP7_75t_L g7190 ( 
.A(n_7105),
.B(n_6811),
.C(n_6660),
.Y(n_7190)
);

AND2x2_ASAP7_75t_L g7191 ( 
.A(n_7036),
.B(n_6806),
.Y(n_7191)
);

NAND2xp5_ASAP7_75t_L g7192 ( 
.A(n_7027),
.B(n_6606),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_7005),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_7030),
.B(n_6609),
.Y(n_7194)
);

NAND2xp5_ASAP7_75t_L g7195 ( 
.A(n_7030),
.B(n_6621),
.Y(n_7195)
);

AOI22xp33_ASAP7_75t_L g7196 ( 
.A1(n_7073),
.A2(n_6796),
.B1(n_6629),
.B2(n_6773),
.Y(n_7196)
);

AND2x2_ASAP7_75t_L g7197 ( 
.A(n_7015),
.B(n_6623),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_L g7198 ( 
.A(n_7105),
.B(n_7088),
.Y(n_7198)
);

NAND2xp5_ASAP7_75t_L g7199 ( 
.A(n_7105),
.B(n_6625),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_SL g7200 ( 
.A(n_7121),
.B(n_6778),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_SL g7201 ( 
.A(n_7116),
.B(n_6744),
.Y(n_7201)
);

NOR3xp33_ASAP7_75t_L g7202 ( 
.A(n_7053),
.B(n_6789),
.C(n_6815),
.Y(n_7202)
);

OA21x2_ASAP7_75t_L g7203 ( 
.A1(n_7048),
.A2(n_6746),
.B(n_6745),
.Y(n_7203)
);

AND2x2_ASAP7_75t_L g7204 ( 
.A(n_7055),
.B(n_6627),
.Y(n_7204)
);

NAND2xp5_ASAP7_75t_L g7205 ( 
.A(n_7043),
.B(n_6628),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_7119),
.B(n_6635),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_SL g7207 ( 
.A(n_7116),
.B(n_6744),
.Y(n_7207)
);

NAND3xp33_ASAP7_75t_L g7208 ( 
.A(n_7083),
.B(n_6789),
.C(n_6730),
.Y(n_7208)
);

AOI21x1_ASAP7_75t_L g7209 ( 
.A1(n_7005),
.A2(n_6746),
.B(n_6791),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_7119),
.B(n_6639),
.Y(n_7210)
);

NAND3xp33_ASAP7_75t_L g7211 ( 
.A(n_7083),
.B(n_6645),
.C(n_6643),
.Y(n_7211)
);

OAI21xp5_ASAP7_75t_SL g7212 ( 
.A1(n_7073),
.A2(n_6648),
.B(n_6646),
.Y(n_7212)
);

AND2x2_ASAP7_75t_L g7213 ( 
.A(n_7047),
.B(n_7041),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_L g7214 ( 
.A(n_7123),
.B(n_6675),
.Y(n_7214)
);

NAND4xp25_ASAP7_75t_L g7215 ( 
.A(n_7029),
.B(n_7082),
.C(n_7023),
.D(n_7009),
.Y(n_7215)
);

NAND2xp5_ASAP7_75t_L g7216 ( 
.A(n_7123),
.B(n_6677),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_7145),
.B(n_6780),
.Y(n_7217)
);

NAND4xp25_ASAP7_75t_L g7218 ( 
.A(n_7022),
.B(n_6804),
.C(n_6791),
.D(n_6780),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_SL g7219 ( 
.A(n_7122),
.B(n_6772),
.Y(n_7219)
);

NAND2xp5_ASAP7_75t_SL g7220 ( 
.A(n_7122),
.B(n_6772),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_7024),
.B(n_6864),
.Y(n_7221)
);

OAI221xp5_ASAP7_75t_SL g7222 ( 
.A1(n_7048),
.A2(n_6804),
.B1(n_6808),
.B2(n_6807),
.C(n_6820),
.Y(n_7222)
);

AND2x2_ASAP7_75t_L g7223 ( 
.A(n_7079),
.B(n_6767),
.Y(n_7223)
);

OAI22xp5_ASAP7_75t_L g7224 ( 
.A1(n_7102),
.A2(n_7054),
.B1(n_7069),
.B2(n_7051),
.Y(n_7224)
);

NAND3xp33_ASAP7_75t_L g7225 ( 
.A(n_7076),
.B(n_6629),
.C(n_6807),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7006),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_7020),
.B(n_6767),
.Y(n_7227)
);

AND2x2_ASAP7_75t_L g7228 ( 
.A(n_7049),
.B(n_6767),
.Y(n_7228)
);

NAND2xp5_ASAP7_75t_L g7229 ( 
.A(n_7024),
.B(n_6796),
.Y(n_7229)
);

HB1xp67_ASAP7_75t_L g7230 ( 
.A(n_7006),
.Y(n_7230)
);

NOR3xp33_ASAP7_75t_L g7231 ( 
.A(n_7070),
.B(n_6622),
.C(n_6680),
.Y(n_7231)
);

AOI21xp33_ASAP7_75t_L g7232 ( 
.A1(n_7139),
.A2(n_6808),
.B(n_6820),
.Y(n_7232)
);

AND2x2_ASAP7_75t_L g7233 ( 
.A(n_7130),
.B(n_6892),
.Y(n_7233)
);

NAND2xp5_ASAP7_75t_L g7234 ( 
.A(n_7090),
.B(n_6821),
.Y(n_7234)
);

NAND2xp5_ASAP7_75t_L g7235 ( 
.A(n_7090),
.B(n_6821),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_7133),
.B(n_6697),
.Y(n_7236)
);

AOI22xp33_ASAP7_75t_SL g7237 ( 
.A1(n_7035),
.A2(n_6637),
.B1(n_6987),
.B2(n_6892),
.Y(n_7237)
);

OAI221xp5_ASAP7_75t_SL g7238 ( 
.A1(n_7102),
.A2(n_6987),
.B1(n_6892),
.B2(n_6905),
.C(n_445),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7136),
.B(n_6905),
.Y(n_7239)
);

AND2x2_ASAP7_75t_L g7240 ( 
.A(n_7113),
.B(n_442),
.Y(n_7240)
);

OAI221xp5_ASAP7_75t_SL g7241 ( 
.A1(n_7094),
.A2(n_447),
.B1(n_444),
.B2(n_445),
.C(n_448),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_7133),
.B(n_450),
.Y(n_7242)
);

AND2x2_ASAP7_75t_L g7243 ( 
.A(n_7127),
.B(n_7103),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_7093),
.B(n_7107),
.Y(n_7244)
);

OAI21xp5_ASAP7_75t_SL g7245 ( 
.A1(n_7086),
.A2(n_450),
.B(n_451),
.Y(n_7245)
);

NAND2xp5_ASAP7_75t_L g7246 ( 
.A(n_7093),
.B(n_7068),
.Y(n_7246)
);

OAI22xp5_ASAP7_75t_L g7247 ( 
.A1(n_7051),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7068),
.B(n_456),
.Y(n_7248)
);

OAI221xp5_ASAP7_75t_L g7249 ( 
.A1(n_7146),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_7100),
.B(n_457),
.Y(n_7250)
);

OAI221xp5_ASAP7_75t_L g7251 ( 
.A1(n_7040),
.A2(n_459),
.B1(n_460),
.B2(n_462),
.C(n_463),
.Y(n_7251)
);

AOI21xp5_ASAP7_75t_SL g7252 ( 
.A1(n_7139),
.A2(n_462),
.B(n_464),
.Y(n_7252)
);

NAND4xp25_ASAP7_75t_L g7253 ( 
.A(n_7028),
.B(n_466),
.C(n_464),
.D(n_465),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_L g7254 ( 
.A(n_7019),
.B(n_465),
.Y(n_7254)
);

NAND3xp33_ASAP7_75t_L g7255 ( 
.A(n_7035),
.B(n_468),
.C(n_469),
.Y(n_7255)
);

NAND2xp5_ASAP7_75t_L g7256 ( 
.A(n_7019),
.B(n_471),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_L g7257 ( 
.A(n_7114),
.B(n_472),
.Y(n_7257)
);

OAI22xp5_ASAP7_75t_L g7258 ( 
.A1(n_7054),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_SL g7259 ( 
.A(n_7091),
.B(n_3421),
.Y(n_7259)
);

OAI21xp5_ASAP7_75t_SL g7260 ( 
.A1(n_7115),
.A2(n_473),
.B(n_476),
.Y(n_7260)
);

AND2x2_ASAP7_75t_L g7261 ( 
.A(n_7147),
.B(n_476),
.Y(n_7261)
);

AND2x2_ASAP7_75t_L g7262 ( 
.A(n_7112),
.B(n_477),
.Y(n_7262)
);

OAI22xp33_ASAP7_75t_L g7263 ( 
.A1(n_7069),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_7263)
);

INVx2_ASAP7_75t_L g7264 ( 
.A(n_7014),
.Y(n_7264)
);

AND2x2_ASAP7_75t_L g7265 ( 
.A(n_7081),
.B(n_479),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7014),
.Y(n_7266)
);

OAI211xp5_ASAP7_75t_L g7267 ( 
.A1(n_7046),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_7267)
);

NAND3xp33_ASAP7_75t_L g7268 ( 
.A(n_7046),
.B(n_483),
.C(n_484),
.Y(n_7268)
);

NAND3xp33_ASAP7_75t_L g7269 ( 
.A(n_7058),
.B(n_483),
.C(n_484),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_7016),
.Y(n_7270)
);

NOR2xp33_ASAP7_75t_L g7271 ( 
.A(n_7042),
.B(n_485),
.Y(n_7271)
);

AOI22xp33_ASAP7_75t_SL g7272 ( 
.A1(n_7058),
.A2(n_7089),
.B1(n_7118),
.B2(n_7060),
.Y(n_7272)
);

NAND2xp5_ASAP7_75t_L g7273 ( 
.A(n_7071),
.B(n_7140),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_7071),
.B(n_487),
.Y(n_7274)
);

AOI22xp33_ASAP7_75t_L g7275 ( 
.A1(n_7120),
.A2(n_2397),
.B1(n_2352),
.B2(n_2288),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_L g7276 ( 
.A(n_7140),
.B(n_487),
.Y(n_7276)
);

AOI22xp33_ASAP7_75t_L g7277 ( 
.A1(n_7078),
.A2(n_2397),
.B1(n_2352),
.B2(n_2288),
.Y(n_7277)
);

OAI221xp5_ASAP7_75t_SL g7278 ( 
.A1(n_7134),
.A2(n_488),
.B1(n_490),
.B2(n_491),
.C(n_493),
.Y(n_7278)
);

NAND2xp5_ASAP7_75t_L g7279 ( 
.A(n_7016),
.B(n_488),
.Y(n_7279)
);

NAND3xp33_ASAP7_75t_L g7280 ( 
.A(n_7060),
.B(n_493),
.C(n_494),
.Y(n_7280)
);

AND2x2_ASAP7_75t_L g7281 ( 
.A(n_7067),
.B(n_494),
.Y(n_7281)
);

AND2x2_ASAP7_75t_L g7282 ( 
.A(n_7066),
.B(n_495),
.Y(n_7282)
);

NAND3xp33_ASAP7_75t_L g7283 ( 
.A(n_7089),
.B(n_496),
.C(n_497),
.Y(n_7283)
);

AND2x2_ASAP7_75t_L g7284 ( 
.A(n_7059),
.B(n_496),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_7118),
.B(n_498),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_7230),
.Y(n_7286)
);

AND2x2_ASAP7_75t_L g7287 ( 
.A(n_7157),
.B(n_7117),
.Y(n_7287)
);

INVx1_ASAP7_75t_L g7288 ( 
.A(n_7209),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_7149),
.B(n_7064),
.Y(n_7289)
);

HB1xp67_ASAP7_75t_L g7290 ( 
.A(n_7203),
.Y(n_7290)
);

INVx2_ASAP7_75t_L g7291 ( 
.A(n_7213),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_7264),
.Y(n_7292)
);

BUFx2_ASAP7_75t_SL g7293 ( 
.A(n_7153),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7148),
.Y(n_7294)
);

BUFx2_ASAP7_75t_L g7295 ( 
.A(n_7193),
.Y(n_7295)
);

OR2x2_ASAP7_75t_L g7296 ( 
.A(n_7198),
.B(n_7039),
.Y(n_7296)
);

INVx2_ASAP7_75t_L g7297 ( 
.A(n_7191),
.Y(n_7297)
);

INVx2_ASAP7_75t_L g7298 ( 
.A(n_7243),
.Y(n_7298)
);

HB1xp67_ASAP7_75t_L g7299 ( 
.A(n_7203),
.Y(n_7299)
);

INVx2_ASAP7_75t_L g7300 ( 
.A(n_7180),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_L g7301 ( 
.A(n_7272),
.B(n_7095),
.Y(n_7301)
);

AND2x2_ASAP7_75t_L g7302 ( 
.A(n_7182),
.B(n_7080),
.Y(n_7302)
);

AND2x2_ASAP7_75t_SL g7303 ( 
.A(n_7150),
.B(n_7134),
.Y(n_7303)
);

BUFx3_ASAP7_75t_L g7304 ( 
.A(n_7226),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_7266),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_7270),
.Y(n_7306)
);

BUFx2_ASAP7_75t_L g7307 ( 
.A(n_7273),
.Y(n_7307)
);

NAND2xp5_ASAP7_75t_L g7308 ( 
.A(n_7233),
.B(n_7095),
.Y(n_7308)
);

AND2x2_ASAP7_75t_L g7309 ( 
.A(n_7197),
.B(n_7097),
.Y(n_7309)
);

INVxp67_ASAP7_75t_L g7310 ( 
.A(n_7164),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_L g7311 ( 
.A(n_7239),
.B(n_7096),
.Y(n_7311)
);

NAND2xp5_ASAP7_75t_L g7312 ( 
.A(n_7165),
.B(n_7096),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_7246),
.Y(n_7313)
);

INVx1_ASAP7_75t_SL g7314 ( 
.A(n_7173),
.Y(n_7314)
);

BUFx2_ASAP7_75t_L g7315 ( 
.A(n_7228),
.Y(n_7315)
);

OR2x2_ASAP7_75t_L g7316 ( 
.A(n_7186),
.B(n_7044),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_7158),
.B(n_7101),
.Y(n_7317)
);

AND2x2_ASAP7_75t_L g7318 ( 
.A(n_7240),
.B(n_7098),
.Y(n_7318)
);

AND2x2_ASAP7_75t_L g7319 ( 
.A(n_7281),
.B(n_7099),
.Y(n_7319)
);

AND2x2_ASAP7_75t_L g7320 ( 
.A(n_7202),
.B(n_7104),
.Y(n_7320)
);

NAND2xp5_ASAP7_75t_L g7321 ( 
.A(n_7170),
.B(n_7101),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_7242),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_7265),
.Y(n_7323)
);

INVx2_ASAP7_75t_L g7324 ( 
.A(n_7181),
.Y(n_7324)
);

NOR2x1_ASAP7_75t_L g7325 ( 
.A(n_7252),
.B(n_7135),
.Y(n_7325)
);

AND2x2_ASAP7_75t_L g7326 ( 
.A(n_7282),
.B(n_7091),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_7250),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_7262),
.Y(n_7328)
);

AND2x2_ASAP7_75t_L g7329 ( 
.A(n_7204),
.B(n_7138),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_7284),
.B(n_7141),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7172),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_7261),
.B(n_7109),
.Y(n_7332)
);

BUFx2_ASAP7_75t_L g7333 ( 
.A(n_7162),
.Y(n_7333)
);

INVx2_ASAP7_75t_L g7334 ( 
.A(n_7223),
.Y(n_7334)
);

AND2x2_ASAP7_75t_L g7335 ( 
.A(n_7185),
.B(n_7129),
.Y(n_7335)
);

NAND2xp5_ASAP7_75t_L g7336 ( 
.A(n_7224),
.B(n_7106),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7175),
.Y(n_7337)
);

INVx4_ASAP7_75t_SL g7338 ( 
.A(n_7285),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_7244),
.Y(n_7339)
);

AND2x2_ASAP7_75t_L g7340 ( 
.A(n_7154),
.B(n_7132),
.Y(n_7340)
);

AND2x4_ASAP7_75t_L g7341 ( 
.A(n_7200),
.B(n_7008),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7224),
.B(n_7106),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_7163),
.B(n_7045),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_L g7344 ( 
.A(n_7237),
.B(n_7018),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7178),
.B(n_7017),
.Y(n_7345)
);

INVx2_ASAP7_75t_L g7346 ( 
.A(n_7248),
.Y(n_7346)
);

HB1xp67_ASAP7_75t_L g7347 ( 
.A(n_7190),
.Y(n_7347)
);

NAND2xp5_ASAP7_75t_L g7348 ( 
.A(n_7201),
.B(n_7207),
.Y(n_7348)
);

AND2x2_ASAP7_75t_L g7349 ( 
.A(n_7271),
.B(n_7217),
.Y(n_7349)
);

BUFx3_ASAP7_75t_L g7350 ( 
.A(n_7156),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_7234),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_7235),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7276),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_7274),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_7227),
.Y(n_7355)
);

AND2x4_ASAP7_75t_SL g7356 ( 
.A(n_7166),
.B(n_7031),
.Y(n_7356)
);

AND2x2_ASAP7_75t_L g7357 ( 
.A(n_7169),
.B(n_7017),
.Y(n_7357)
);

AND2x2_ASAP7_75t_L g7358 ( 
.A(n_7161),
.B(n_7057),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_7183),
.Y(n_7359)
);

AND2x4_ASAP7_75t_L g7360 ( 
.A(n_7219),
.B(n_7033),
.Y(n_7360)
);

OAI322xp33_ASAP7_75t_L g7361 ( 
.A1(n_7159),
.A2(n_7142),
.A3(n_7135),
.B1(n_7037),
.B2(n_7061),
.C1(n_7074),
.C2(n_7063),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_7254),
.Y(n_7362)
);

OR2x2_ASAP7_75t_L g7363 ( 
.A(n_7160),
.B(n_7050),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_7256),
.Y(n_7364)
);

HB1xp67_ASAP7_75t_L g7365 ( 
.A(n_7187),
.Y(n_7365)
);

AND2x2_ASAP7_75t_L g7366 ( 
.A(n_7220),
.B(n_7065),
.Y(n_7366)
);

INVxp67_ASAP7_75t_SL g7367 ( 
.A(n_7187),
.Y(n_7367)
);

AND2x4_ASAP7_75t_L g7368 ( 
.A(n_7177),
.B(n_7085),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_7279),
.Y(n_7369)
);

HB1xp67_ASAP7_75t_L g7370 ( 
.A(n_7285),
.Y(n_7370)
);

OR2x2_ASAP7_75t_L g7371 ( 
.A(n_7215),
.B(n_7092),
.Y(n_7371)
);

OR2x2_ASAP7_75t_L g7372 ( 
.A(n_7152),
.B(n_7110),
.Y(n_7372)
);

AND2x2_ASAP7_75t_L g7373 ( 
.A(n_7205),
.B(n_7085),
.Y(n_7373)
);

INVxp67_ASAP7_75t_L g7374 ( 
.A(n_7156),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_7257),
.B(n_7084),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_7279),
.Y(n_7376)
);

AND2x4_ASAP7_75t_SL g7377 ( 
.A(n_7151),
.B(n_7142),
.Y(n_7377)
);

AND2x2_ASAP7_75t_L g7378 ( 
.A(n_7221),
.B(n_7188),
.Y(n_7378)
);

BUFx2_ASAP7_75t_L g7379 ( 
.A(n_7199),
.Y(n_7379)
);

HB1xp67_ASAP7_75t_L g7380 ( 
.A(n_7208),
.Y(n_7380)
);

OR2x2_ASAP7_75t_L g7381 ( 
.A(n_7152),
.B(n_7126),
.Y(n_7381)
);

INVx1_ASAP7_75t_L g7382 ( 
.A(n_7192),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_7194),
.Y(n_7383)
);

INVx2_ASAP7_75t_L g7384 ( 
.A(n_7195),
.Y(n_7384)
);

AND2x2_ASAP7_75t_L g7385 ( 
.A(n_7159),
.B(n_7236),
.Y(n_7385)
);

NAND2xp5_ASAP7_75t_L g7386 ( 
.A(n_7155),
.B(n_498),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_7206),
.Y(n_7387)
);

INVxp67_ASAP7_75t_L g7388 ( 
.A(n_7255),
.Y(n_7388)
);

INVxp67_ASAP7_75t_L g7389 ( 
.A(n_7268),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_7210),
.Y(n_7390)
);

NAND2xp5_ASAP7_75t_L g7391 ( 
.A(n_7167),
.B(n_499),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_7214),
.Y(n_7392)
);

NAND2xp5_ASAP7_75t_L g7393 ( 
.A(n_7176),
.B(n_499),
.Y(n_7393)
);

INVx3_ASAP7_75t_L g7394 ( 
.A(n_7216),
.Y(n_7394)
);

AND2x2_ASAP7_75t_L g7395 ( 
.A(n_7245),
.B(n_500),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7211),
.Y(n_7396)
);

INVx2_ASAP7_75t_L g7397 ( 
.A(n_7229),
.Y(n_7397)
);

INVx3_ASAP7_75t_L g7398 ( 
.A(n_7174),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_7247),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_7247),
.Y(n_7400)
);

AND2x2_ASAP7_75t_L g7401 ( 
.A(n_7171),
.B(n_500),
.Y(n_7401)
);

BUFx3_ASAP7_75t_L g7402 ( 
.A(n_7269),
.Y(n_7402)
);

INVx2_ASAP7_75t_L g7403 ( 
.A(n_7259),
.Y(n_7403)
);

AND2x4_ASAP7_75t_L g7404 ( 
.A(n_7280),
.B(n_503),
.Y(n_7404)
);

BUFx2_ASAP7_75t_L g7405 ( 
.A(n_7290),
.Y(n_7405)
);

INVx2_ASAP7_75t_L g7406 ( 
.A(n_7290),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_7299),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_7299),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_7303),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_7303),
.Y(n_7410)
);

HB1xp67_ASAP7_75t_L g7411 ( 
.A(n_7338),
.Y(n_7411)
);

INVx4_ASAP7_75t_L g7412 ( 
.A(n_7304),
.Y(n_7412)
);

INVx2_ASAP7_75t_L g7413 ( 
.A(n_7288),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_SL g7414 ( 
.A(n_7348),
.B(n_7196),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7295),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_7304),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7296),
.Y(n_7417)
);

NOR3xp33_ASAP7_75t_SL g7418 ( 
.A(n_7361),
.B(n_7222),
.C(n_7179),
.Y(n_7418)
);

INVx2_ASAP7_75t_L g7419 ( 
.A(n_7350),
.Y(n_7419)
);

INVx1_ASAP7_75t_L g7420 ( 
.A(n_7338),
.Y(n_7420)
);

INVxp33_ASAP7_75t_SL g7421 ( 
.A(n_7293),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_7338),
.Y(n_7422)
);

INVx2_ASAP7_75t_L g7423 ( 
.A(n_7350),
.Y(n_7423)
);

BUFx8_ASAP7_75t_L g7424 ( 
.A(n_7286),
.Y(n_7424)
);

HB1xp67_ASAP7_75t_L g7425 ( 
.A(n_7325),
.Y(n_7425)
);

INVx2_ASAP7_75t_SL g7426 ( 
.A(n_7360),
.Y(n_7426)
);

INVx4_ASAP7_75t_SL g7427 ( 
.A(n_7294),
.Y(n_7427)
);

INVx1_ASAP7_75t_L g7428 ( 
.A(n_7329),
.Y(n_7428)
);

BUFx2_ASAP7_75t_L g7429 ( 
.A(n_7341),
.Y(n_7429)
);

OAI21x1_ASAP7_75t_L g7430 ( 
.A1(n_7336),
.A2(n_7225),
.B(n_7184),
.Y(n_7430)
);

INVxp67_ASAP7_75t_SL g7431 ( 
.A(n_7336),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_7309),
.Y(n_7432)
);

INVx2_ASAP7_75t_L g7433 ( 
.A(n_7365),
.Y(n_7433)
);

INVx2_ASAP7_75t_L g7434 ( 
.A(n_7365),
.Y(n_7434)
);

OAI21x1_ASAP7_75t_L g7435 ( 
.A1(n_7342),
.A2(n_7168),
.B(n_7258),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7332),
.Y(n_7436)
);

NOR2xp33_ASAP7_75t_L g7437 ( 
.A(n_7398),
.B(n_7238),
.Y(n_7437)
);

AND2x2_ASAP7_75t_L g7438 ( 
.A(n_7289),
.B(n_7212),
.Y(n_7438)
);

OA21x2_ASAP7_75t_L g7439 ( 
.A1(n_7301),
.A2(n_7232),
.B(n_7231),
.Y(n_7439)
);

BUFx3_ASAP7_75t_L g7440 ( 
.A(n_7287),
.Y(n_7440)
);

INVx2_ASAP7_75t_L g7441 ( 
.A(n_7341),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_7330),
.Y(n_7442)
);

INVx4_ASAP7_75t_SL g7443 ( 
.A(n_7305),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7316),
.Y(n_7444)
);

AND2x2_ASAP7_75t_L g7445 ( 
.A(n_7314),
.B(n_7232),
.Y(n_7445)
);

INVx2_ASAP7_75t_L g7446 ( 
.A(n_7342),
.Y(n_7446)
);

INVxp67_ASAP7_75t_SL g7447 ( 
.A(n_7348),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_7334),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_7334),
.Y(n_7449)
);

OA21x2_ASAP7_75t_L g7450 ( 
.A1(n_7301),
.A2(n_7283),
.B(n_7218),
.Y(n_7450)
);

BUFx6f_ASAP7_75t_L g7451 ( 
.A(n_7386),
.Y(n_7451)
);

NAND2xp5_ASAP7_75t_L g7452 ( 
.A(n_7314),
.B(n_7260),
.Y(n_7452)
);

HB1xp67_ASAP7_75t_L g7453 ( 
.A(n_7315),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_7319),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_L g7455 ( 
.A(n_7398),
.B(n_7267),
.Y(n_7455)
);

OAI21x1_ASAP7_75t_L g7456 ( 
.A1(n_7367),
.A2(n_7258),
.B(n_7253),
.Y(n_7456)
);

NAND3xp33_ASAP7_75t_SL g7457 ( 
.A(n_7386),
.B(n_7249),
.C(n_7251),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7318),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_7302),
.Y(n_7459)
);

NAND2xp5_ASAP7_75t_L g7460 ( 
.A(n_7310),
.B(n_7263),
.Y(n_7460)
);

INVx2_ASAP7_75t_L g7461 ( 
.A(n_7360),
.Y(n_7461)
);

AND2x2_ASAP7_75t_L g7462 ( 
.A(n_7326),
.B(n_7189),
.Y(n_7462)
);

INVx3_ASAP7_75t_L g7463 ( 
.A(n_7368),
.Y(n_7463)
);

HB1xp67_ASAP7_75t_L g7464 ( 
.A(n_7370),
.Y(n_7464)
);

INVxp67_ASAP7_75t_SL g7465 ( 
.A(n_7380),
.Y(n_7465)
);

AND2x2_ASAP7_75t_L g7466 ( 
.A(n_7310),
.B(n_7275),
.Y(n_7466)
);

INVx2_ASAP7_75t_L g7467 ( 
.A(n_7356),
.Y(n_7467)
);

OAI21xp5_ASAP7_75t_SL g7468 ( 
.A1(n_7377),
.A2(n_7277),
.B(n_7241),
.Y(n_7468)
);

AOI21x1_ASAP7_75t_L g7469 ( 
.A1(n_7347),
.A2(n_7278),
.B(n_503),
.Y(n_7469)
);

NAND3xp33_ASAP7_75t_L g7470 ( 
.A(n_7380),
.B(n_505),
.C(n_507),
.Y(n_7470)
);

INVx3_ASAP7_75t_L g7471 ( 
.A(n_7368),
.Y(n_7471)
);

OR2x2_ASAP7_75t_L g7472 ( 
.A(n_7367),
.B(n_508),
.Y(n_7472)
);

INVx2_ASAP7_75t_L g7473 ( 
.A(n_7356),
.Y(n_7473)
);

HB1xp67_ASAP7_75t_L g7474 ( 
.A(n_7370),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7298),
.Y(n_7475)
);

OR2x6_ASAP7_75t_L g7476 ( 
.A(n_7374),
.B(n_7393),
.Y(n_7476)
);

INVx2_ASAP7_75t_L g7477 ( 
.A(n_7347),
.Y(n_7477)
);

INVx2_ASAP7_75t_L g7478 ( 
.A(n_7355),
.Y(n_7478)
);

INVx2_ASAP7_75t_L g7479 ( 
.A(n_7340),
.Y(n_7479)
);

INVx3_ASAP7_75t_L g7480 ( 
.A(n_7377),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_7291),
.Y(n_7481)
);

HB1xp67_ASAP7_75t_L g7482 ( 
.A(n_7366),
.Y(n_7482)
);

INVx3_ASAP7_75t_L g7483 ( 
.A(n_7297),
.Y(n_7483)
);

AND2x2_ASAP7_75t_L g7484 ( 
.A(n_7345),
.B(n_509),
.Y(n_7484)
);

NOR2x1p5_ASAP7_75t_L g7485 ( 
.A(n_7300),
.B(n_509),
.Y(n_7485)
);

INVx2_ASAP7_75t_L g7486 ( 
.A(n_7381),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_7307),
.Y(n_7487)
);

INVx1_ASAP7_75t_L g7488 ( 
.A(n_7333),
.Y(n_7488)
);

HB1xp67_ASAP7_75t_L g7489 ( 
.A(n_7374),
.Y(n_7489)
);

OA21x2_ASAP7_75t_L g7490 ( 
.A1(n_7393),
.A2(n_510),
.B(n_511),
.Y(n_7490)
);

INVx2_ASAP7_75t_L g7491 ( 
.A(n_7320),
.Y(n_7491)
);

INVx2_ASAP7_75t_L g7492 ( 
.A(n_7357),
.Y(n_7492)
);

AND2x2_ASAP7_75t_L g7493 ( 
.A(n_7440),
.B(n_7358),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_7480),
.B(n_7401),
.Y(n_7494)
);

INVx2_ASAP7_75t_L g7495 ( 
.A(n_7405),
.Y(n_7495)
);

NAND2xp5_ASAP7_75t_L g7496 ( 
.A(n_7480),
.B(n_7385),
.Y(n_7496)
);

INVxp67_ASAP7_75t_L g7497 ( 
.A(n_7429),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7405),
.Y(n_7498)
);

INVx3_ASAP7_75t_L g7499 ( 
.A(n_7412),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7440),
.B(n_7438),
.Y(n_7500)
);

OR2x2_ASAP7_75t_L g7501 ( 
.A(n_7426),
.B(n_7308),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_7406),
.Y(n_7502)
);

HB1xp67_ASAP7_75t_L g7503 ( 
.A(n_7406),
.Y(n_7503)
);

HB1xp67_ASAP7_75t_L g7504 ( 
.A(n_7407),
.Y(n_7504)
);

INVx1_ASAP7_75t_L g7505 ( 
.A(n_7453),
.Y(n_7505)
);

INVx2_ASAP7_75t_L g7506 ( 
.A(n_7408),
.Y(n_7506)
);

INVx2_ASAP7_75t_SL g7507 ( 
.A(n_7426),
.Y(n_7507)
);

CKINVDCx20_ASAP7_75t_R g7508 ( 
.A(n_7424),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7411),
.Y(n_7509)
);

AND2x2_ASAP7_75t_L g7510 ( 
.A(n_7438),
.B(n_7335),
.Y(n_7510)
);

AND2x2_ASAP7_75t_L g7511 ( 
.A(n_7467),
.B(n_7343),
.Y(n_7511)
);

OR2x2_ASAP7_75t_L g7512 ( 
.A(n_7480),
.B(n_7308),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_7427),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7427),
.Y(n_7514)
);

AND2x4_ASAP7_75t_L g7515 ( 
.A(n_7427),
.B(n_7292),
.Y(n_7515)
);

AND2x2_ASAP7_75t_L g7516 ( 
.A(n_7467),
.B(n_7378),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7427),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7464),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7421),
.B(n_7311),
.Y(n_7519)
);

INVx1_ASAP7_75t_L g7520 ( 
.A(n_7474),
.Y(n_7520)
);

HB1xp67_ASAP7_75t_L g7521 ( 
.A(n_7445),
.Y(n_7521)
);

INVx2_ASAP7_75t_L g7522 ( 
.A(n_7463),
.Y(n_7522)
);

INVx2_ASAP7_75t_L g7523 ( 
.A(n_7463),
.Y(n_7523)
);

HB1xp67_ASAP7_75t_L g7524 ( 
.A(n_7445),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7463),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_7421),
.B(n_7471),
.Y(n_7526)
);

AND2x2_ASAP7_75t_L g7527 ( 
.A(n_7473),
.B(n_7313),
.Y(n_7527)
);

BUFx2_ASAP7_75t_L g7528 ( 
.A(n_7412),
.Y(n_7528)
);

INVx1_ASAP7_75t_L g7529 ( 
.A(n_7471),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_7471),
.Y(n_7530)
);

AND2x2_ASAP7_75t_L g7531 ( 
.A(n_7473),
.B(n_7323),
.Y(n_7531)
);

NAND2xp5_ASAP7_75t_L g7532 ( 
.A(n_7462),
.B(n_7311),
.Y(n_7532)
);

INVx2_ASAP7_75t_L g7533 ( 
.A(n_7412),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_L g7534 ( 
.A(n_7462),
.B(n_7399),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_7443),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_7428),
.B(n_7482),
.Y(n_7536)
);

NAND2xp5_ASAP7_75t_L g7537 ( 
.A(n_7437),
.B(n_7400),
.Y(n_7537)
);

INVx2_ASAP7_75t_L g7538 ( 
.A(n_7439),
.Y(n_7538)
);

AND2x2_ASAP7_75t_L g7539 ( 
.A(n_7436),
.B(n_7327),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_7443),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7437),
.B(n_7395),
.Y(n_7541)
);

AND2x2_ASAP7_75t_L g7542 ( 
.A(n_7442),
.B(n_7328),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7443),
.Y(n_7543)
);

INVxp67_ASAP7_75t_L g7544 ( 
.A(n_7425),
.Y(n_7544)
);

NOR2xp33_ASAP7_75t_L g7545 ( 
.A(n_7483),
.B(n_7317),
.Y(n_7545)
);

INVx1_ASAP7_75t_L g7546 ( 
.A(n_7443),
.Y(n_7546)
);

INVxp67_ASAP7_75t_L g7547 ( 
.A(n_7489),
.Y(n_7547)
);

NAND2xp5_ASAP7_75t_L g7548 ( 
.A(n_7483),
.B(n_7404),
.Y(n_7548)
);

INVx2_ASAP7_75t_L g7549 ( 
.A(n_7439),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7483),
.Y(n_7550)
);

INVxp67_ASAP7_75t_SL g7551 ( 
.A(n_7409),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7419),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_7409),
.B(n_7404),
.Y(n_7553)
);

AND2x2_ASAP7_75t_L g7554 ( 
.A(n_7454),
.B(n_7324),
.Y(n_7554)
);

INVx2_ASAP7_75t_SL g7555 ( 
.A(n_7424),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_7458),
.B(n_7349),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_7419),
.Y(n_7557)
);

NAND2xp5_ASAP7_75t_L g7558 ( 
.A(n_7410),
.B(n_7312),
.Y(n_7558)
);

NAND2xp5_ASAP7_75t_L g7559 ( 
.A(n_7410),
.B(n_7312),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7439),
.Y(n_7560)
);

AND2x2_ASAP7_75t_L g7561 ( 
.A(n_7459),
.B(n_7375),
.Y(n_7561)
);

NOR2xp33_ASAP7_75t_L g7562 ( 
.A(n_7451),
.B(n_7317),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_7423),
.Y(n_7563)
);

INVx2_ASAP7_75t_L g7564 ( 
.A(n_7441),
.Y(n_7564)
);

NAND2xp5_ASAP7_75t_L g7565 ( 
.A(n_7431),
.B(n_7373),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7432),
.B(n_7479),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7423),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7441),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_7461),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_7503),
.Y(n_7570)
);

INVx1_ASAP7_75t_SL g7571 ( 
.A(n_7508),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7503),
.Y(n_7572)
);

AOI22xp5_ASAP7_75t_L g7573 ( 
.A1(n_7508),
.A2(n_7344),
.B1(n_7414),
.B2(n_7391),
.Y(n_7573)
);

AND2x2_ASAP7_75t_L g7574 ( 
.A(n_7500),
.B(n_7479),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_L g7575 ( 
.A(n_7507),
.B(n_7484),
.Y(n_7575)
);

OAI211xp5_ASAP7_75t_SL g7576 ( 
.A1(n_7537),
.A2(n_7418),
.B(n_7414),
.C(n_7344),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7522),
.Y(n_7577)
);

INVx3_ASAP7_75t_L g7578 ( 
.A(n_7515),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7522),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_7523),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7523),
.Y(n_7581)
);

OR2x2_ASAP7_75t_L g7582 ( 
.A(n_7512),
.B(n_7461),
.Y(n_7582)
);

OAI21xp33_ASAP7_75t_L g7583 ( 
.A1(n_7558),
.A2(n_7321),
.B(n_7455),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_7521),
.Y(n_7584)
);

BUFx2_ASAP7_75t_L g7585 ( 
.A(n_7497),
.Y(n_7585)
);

INVx1_ASAP7_75t_L g7586 ( 
.A(n_7521),
.Y(n_7586)
);

OR2x2_ASAP7_75t_L g7587 ( 
.A(n_7532),
.B(n_7501),
.Y(n_7587)
);

NAND2xp5_ASAP7_75t_L g7588 ( 
.A(n_7555),
.B(n_7484),
.Y(n_7588)
);

AND2x4_ASAP7_75t_SL g7589 ( 
.A(n_7493),
.B(n_7416),
.Y(n_7589)
);

AOI32xp33_ASAP7_75t_L g7590 ( 
.A1(n_7538),
.A2(n_7396),
.A3(n_7321),
.B1(n_7465),
.B2(n_7402),
.Y(n_7590)
);

INVx2_ASAP7_75t_L g7591 ( 
.A(n_7515),
.Y(n_7591)
);

NAND2xp5_ASAP7_75t_L g7592 ( 
.A(n_7524),
.B(n_7451),
.Y(n_7592)
);

INVx2_ASAP7_75t_L g7593 ( 
.A(n_7515),
.Y(n_7593)
);

AND2x2_ASAP7_75t_L g7594 ( 
.A(n_7510),
.B(n_7511),
.Y(n_7594)
);

INVx2_ASAP7_75t_L g7595 ( 
.A(n_7495),
.Y(n_7595)
);

AND2x2_ASAP7_75t_L g7596 ( 
.A(n_7531),
.B(n_7492),
.Y(n_7596)
);

AND2x4_ASAP7_75t_L g7597 ( 
.A(n_7497),
.B(n_7415),
.Y(n_7597)
);

NAND2xp5_ASAP7_75t_L g7598 ( 
.A(n_7524),
.B(n_7451),
.Y(n_7598)
);

INVx1_ASAP7_75t_SL g7599 ( 
.A(n_7528),
.Y(n_7599)
);

NAND2xp5_ASAP7_75t_L g7600 ( 
.A(n_7551),
.B(n_7451),
.Y(n_7600)
);

AND2x2_ASAP7_75t_L g7601 ( 
.A(n_7516),
.B(n_7492),
.Y(n_7601)
);

INVx1_ASAP7_75t_L g7602 ( 
.A(n_7495),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_7504),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7504),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_7551),
.B(n_7433),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_7526),
.Y(n_7606)
);

OR2x2_ASAP7_75t_L g7607 ( 
.A(n_7519),
.B(n_7452),
.Y(n_7607)
);

INVx1_ASAP7_75t_SL g7608 ( 
.A(n_7496),
.Y(n_7608)
);

NAND2xp5_ASAP7_75t_L g7609 ( 
.A(n_7525),
.B(n_7433),
.Y(n_7609)
);

NAND2xp5_ASAP7_75t_L g7610 ( 
.A(n_7529),
.B(n_7434),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_7499),
.Y(n_7611)
);

NAND2xp5_ASAP7_75t_L g7612 ( 
.A(n_7530),
.B(n_7434),
.Y(n_7612)
);

AND2x2_ASAP7_75t_L g7613 ( 
.A(n_7527),
.B(n_7486),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_7499),
.Y(n_7614)
);

AND2x2_ASAP7_75t_L g7615 ( 
.A(n_7536),
.B(n_7486),
.Y(n_7615)
);

NAND2xp5_ASAP7_75t_L g7616 ( 
.A(n_7564),
.B(n_7424),
.Y(n_7616)
);

NOR4xp25_ASAP7_75t_L g7617 ( 
.A(n_7538),
.B(n_7446),
.C(n_7477),
.D(n_7413),
.Y(n_7617)
);

OR2x2_ASAP7_75t_L g7618 ( 
.A(n_7534),
.B(n_7363),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7513),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_7564),
.B(n_7447),
.Y(n_7620)
);

INVx1_ASAP7_75t_SL g7621 ( 
.A(n_7548),
.Y(n_7621)
);

NOR2xp33_ASAP7_75t_L g7622 ( 
.A(n_7494),
.B(n_7388),
.Y(n_7622)
);

NOR2xp33_ASAP7_75t_L g7623 ( 
.A(n_7547),
.B(n_7388),
.Y(n_7623)
);

AND2x4_ASAP7_75t_L g7624 ( 
.A(n_7550),
.B(n_7481),
.Y(n_7624)
);

INVx1_ASAP7_75t_SL g7625 ( 
.A(n_7549),
.Y(n_7625)
);

AND2x2_ASAP7_75t_L g7626 ( 
.A(n_7539),
.B(n_7487),
.Y(n_7626)
);

AND2x2_ASAP7_75t_L g7627 ( 
.A(n_7542),
.B(n_7488),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7514),
.Y(n_7628)
);

OR2x2_ASAP7_75t_L g7629 ( 
.A(n_7559),
.B(n_7460),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_7561),
.B(n_7417),
.Y(n_7630)
);

NAND2xp5_ASAP7_75t_L g7631 ( 
.A(n_7562),
.B(n_7446),
.Y(n_7631)
);

AND2x2_ASAP7_75t_L g7632 ( 
.A(n_7556),
.B(n_7481),
.Y(n_7632)
);

AOI221xp5_ASAP7_75t_L g7633 ( 
.A1(n_7549),
.A2(n_7457),
.B1(n_7477),
.B2(n_7389),
.C(n_7402),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_L g7634 ( 
.A(n_7571),
.B(n_7545),
.Y(n_7634)
);

OR2x2_ASAP7_75t_L g7635 ( 
.A(n_7571),
.B(n_7372),
.Y(n_7635)
);

AND2x4_ASAP7_75t_L g7636 ( 
.A(n_7578),
.B(n_7547),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7578),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7591),
.Y(n_7638)
);

NAND2x1_ASAP7_75t_L g7639 ( 
.A(n_7593),
.B(n_7498),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7592),
.Y(n_7640)
);

NAND2x1p5_ASAP7_75t_L g7641 ( 
.A(n_7585),
.B(n_7505),
.Y(n_7641)
);

INVxp67_ASAP7_75t_L g7642 ( 
.A(n_7598),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_7594),
.Y(n_7643)
);

INVx1_ASAP7_75t_L g7644 ( 
.A(n_7600),
.Y(n_7644)
);

OR2x2_ASAP7_75t_L g7645 ( 
.A(n_7582),
.B(n_7553),
.Y(n_7645)
);

INVxp67_ASAP7_75t_SL g7646 ( 
.A(n_7605),
.Y(n_7646)
);

NAND2xp5_ASAP7_75t_L g7647 ( 
.A(n_7613),
.B(n_7545),
.Y(n_7647)
);

INVx2_ASAP7_75t_SL g7648 ( 
.A(n_7589),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7584),
.Y(n_7649)
);

NOR2xp33_ASAP7_75t_L g7650 ( 
.A(n_7576),
.B(n_7389),
.Y(n_7650)
);

INVxp67_ASAP7_75t_SL g7651 ( 
.A(n_7586),
.Y(n_7651)
);

OAI21xp5_ASAP7_75t_SL g7652 ( 
.A1(n_7573),
.A2(n_7468),
.B(n_7444),
.Y(n_7652)
);

OR2x2_ASAP7_75t_L g7653 ( 
.A(n_7599),
.B(n_7476),
.Y(n_7653)
);

OR2x2_ASAP7_75t_L g7654 ( 
.A(n_7599),
.B(n_7575),
.Y(n_7654)
);

OR2x2_ASAP7_75t_L g7655 ( 
.A(n_7588),
.B(n_7476),
.Y(n_7655)
);

INVx2_ASAP7_75t_SL g7656 ( 
.A(n_7597),
.Y(n_7656)
);

AND2x2_ASAP7_75t_L g7657 ( 
.A(n_7615),
.B(n_7566),
.Y(n_7657)
);

NOR2xp33_ASAP7_75t_L g7658 ( 
.A(n_7583),
.B(n_7491),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_7625),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7625),
.Y(n_7660)
);

AND2x4_ASAP7_75t_L g7661 ( 
.A(n_7596),
.B(n_7518),
.Y(n_7661)
);

OR2x2_ASAP7_75t_L g7662 ( 
.A(n_7587),
.B(n_7476),
.Y(n_7662)
);

INVx2_ASAP7_75t_L g7663 ( 
.A(n_7570),
.Y(n_7663)
);

AND2x4_ASAP7_75t_L g7664 ( 
.A(n_7597),
.B(n_7520),
.Y(n_7664)
);

INVx3_ASAP7_75t_L g7665 ( 
.A(n_7624),
.Y(n_7665)
);

NAND2xp5_ASAP7_75t_L g7666 ( 
.A(n_7574),
.B(n_7562),
.Y(n_7666)
);

OR2x2_ASAP7_75t_L g7667 ( 
.A(n_7616),
.B(n_7476),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7572),
.Y(n_7668)
);

INVx2_ASAP7_75t_L g7669 ( 
.A(n_7624),
.Y(n_7669)
);

AND2x2_ASAP7_75t_L g7670 ( 
.A(n_7601),
.B(n_7554),
.Y(n_7670)
);

NAND2xp5_ASAP7_75t_L g7671 ( 
.A(n_7573),
.B(n_7509),
.Y(n_7671)
);

NAND2xp5_ASAP7_75t_L g7672 ( 
.A(n_7595),
.B(n_7448),
.Y(n_7672)
);

AND2x2_ASAP7_75t_L g7673 ( 
.A(n_7626),
.B(n_7491),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_7632),
.B(n_7449),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7611),
.Y(n_7675)
);

AND2x2_ASAP7_75t_L g7676 ( 
.A(n_7627),
.B(n_7475),
.Y(n_7676)
);

HB1xp67_ASAP7_75t_L g7677 ( 
.A(n_7603),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7604),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7602),
.B(n_7478),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7631),
.Y(n_7680)
);

AOI22x1_ASAP7_75t_L g7681 ( 
.A1(n_7608),
.A2(n_7560),
.B1(n_7472),
.B2(n_7533),
.Y(n_7681)
);

CKINVDCx16_ASAP7_75t_R g7682 ( 
.A(n_7635),
.Y(n_7682)
);

NOR2xp33_ASAP7_75t_L g7683 ( 
.A(n_7656),
.B(n_7583),
.Y(n_7683)
);

INVx2_ASAP7_75t_L g7684 ( 
.A(n_7665),
.Y(n_7684)
);

NAND4xp25_ASAP7_75t_L g7685 ( 
.A(n_7650),
.B(n_7633),
.C(n_7622),
.D(n_7623),
.Y(n_7685)
);

NAND3xp33_ASAP7_75t_SL g7686 ( 
.A(n_7641),
.B(n_7590),
.C(n_7560),
.Y(n_7686)
);

OAI21xp5_ASAP7_75t_SL g7687 ( 
.A1(n_7652),
.A2(n_7630),
.B(n_7621),
.Y(n_7687)
);

NOR2xp33_ASAP7_75t_SL g7688 ( 
.A(n_7657),
.B(n_7618),
.Y(n_7688)
);

AND2x2_ASAP7_75t_L g7689 ( 
.A(n_7673),
.B(n_7379),
.Y(n_7689)
);

OR2x2_ASAP7_75t_L g7690 ( 
.A(n_7639),
.B(n_7478),
.Y(n_7690)
);

OR2x2_ASAP7_75t_L g7691 ( 
.A(n_7665),
.B(n_7371),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_7636),
.Y(n_7692)
);

OAI22xp5_ASAP7_75t_L g7693 ( 
.A1(n_7648),
.A2(n_7391),
.B1(n_7544),
.B2(n_7470),
.Y(n_7693)
);

INVx2_ASAP7_75t_L g7694 ( 
.A(n_7681),
.Y(n_7694)
);

INVx3_ASAP7_75t_L g7695 ( 
.A(n_7636),
.Y(n_7695)
);

OR2x2_ASAP7_75t_L g7696 ( 
.A(n_7634),
.B(n_7450),
.Y(n_7696)
);

INVx2_ASAP7_75t_L g7697 ( 
.A(n_7681),
.Y(n_7697)
);

INVx1_ASAP7_75t_L g7698 ( 
.A(n_7637),
.Y(n_7698)
);

OR2x2_ASAP7_75t_L g7699 ( 
.A(n_7653),
.B(n_7450),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7637),
.Y(n_7700)
);

NAND2xp5_ASAP7_75t_L g7701 ( 
.A(n_7664),
.B(n_7420),
.Y(n_7701)
);

INVx1_ASAP7_75t_L g7702 ( 
.A(n_7664),
.Y(n_7702)
);

AOI32xp33_ASAP7_75t_L g7703 ( 
.A1(n_7670),
.A2(n_7435),
.A3(n_7430),
.B1(n_7456),
.B2(n_7606),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7677),
.Y(n_7704)
);

NOR2xp67_ASAP7_75t_L g7705 ( 
.A(n_7669),
.B(n_7544),
.Y(n_7705)
);

NAND2xp5_ASAP7_75t_L g7706 ( 
.A(n_7661),
.B(n_7422),
.Y(n_7706)
);

AND2x2_ASAP7_75t_L g7707 ( 
.A(n_7643),
.B(n_7331),
.Y(n_7707)
);

NOR2xp67_ASAP7_75t_L g7708 ( 
.A(n_7662),
.B(n_7533),
.Y(n_7708)
);

NOR2xp33_ASAP7_75t_L g7709 ( 
.A(n_7661),
.B(n_7394),
.Y(n_7709)
);

NOR2xp67_ASAP7_75t_L g7710 ( 
.A(n_7659),
.B(n_7517),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7666),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7660),
.Y(n_7712)
);

OAI21xp33_ASAP7_75t_L g7713 ( 
.A1(n_7688),
.A2(n_7685),
.B(n_7687),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_7695),
.Y(n_7714)
);

AND2x2_ASAP7_75t_L g7715 ( 
.A(n_7689),
.B(n_7676),
.Y(n_7715)
);

INVx1_ASAP7_75t_SL g7716 ( 
.A(n_7690),
.Y(n_7716)
);

INVxp67_ASAP7_75t_L g7717 ( 
.A(n_7695),
.Y(n_7717)
);

INVx1_ASAP7_75t_SL g7718 ( 
.A(n_7691),
.Y(n_7718)
);

OAI21xp5_ASAP7_75t_L g7719 ( 
.A1(n_7708),
.A2(n_7430),
.B(n_7435),
.Y(n_7719)
);

HB1xp67_ASAP7_75t_L g7720 ( 
.A(n_7702),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_7701),
.Y(n_7721)
);

INVx2_ASAP7_75t_L g7722 ( 
.A(n_7692),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_7706),
.Y(n_7723)
);

AOI22xp5_ASAP7_75t_L g7724 ( 
.A1(n_7682),
.A2(n_7337),
.B1(n_7339),
.B2(n_7683),
.Y(n_7724)
);

AND2x2_ASAP7_75t_L g7725 ( 
.A(n_7707),
.B(n_7568),
.Y(n_7725)
);

AOI222xp33_ASAP7_75t_L g7726 ( 
.A1(n_7686),
.A2(n_7413),
.B1(n_7671),
.B2(n_7658),
.C1(n_7502),
.C2(n_7541),
.Y(n_7726)
);

INVxp67_ASAP7_75t_SL g7727 ( 
.A(n_7709),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7684),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_7699),
.Y(n_7729)
);

AND2x2_ASAP7_75t_L g7730 ( 
.A(n_7704),
.B(n_7569),
.Y(n_7730)
);

INVx2_ASAP7_75t_SL g7731 ( 
.A(n_7712),
.Y(n_7731)
);

AOI22xp5_ASAP7_75t_L g7732 ( 
.A1(n_7693),
.A2(n_7450),
.B1(n_7642),
.B2(n_7638),
.Y(n_7732)
);

INVx2_ASAP7_75t_L g7733 ( 
.A(n_7698),
.Y(n_7733)
);

NAND2x1_ASAP7_75t_L g7734 ( 
.A(n_7705),
.B(n_7535),
.Y(n_7734)
);

INVxp67_ASAP7_75t_SL g7735 ( 
.A(n_7710),
.Y(n_7735)
);

OR2x6_ASAP7_75t_L g7736 ( 
.A(n_7712),
.B(n_7647),
.Y(n_7736)
);

INVx2_ASAP7_75t_L g7737 ( 
.A(n_7700),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7696),
.Y(n_7738)
);

OAI221xp5_ASAP7_75t_L g7739 ( 
.A1(n_7703),
.A2(n_7651),
.B1(n_7617),
.B2(n_7610),
.C(n_7612),
.Y(n_7739)
);

AO32x1_ASAP7_75t_L g7740 ( 
.A1(n_7694),
.A2(n_7614),
.A3(n_7580),
.B1(n_7581),
.B2(n_7579),
.Y(n_7740)
);

NAND2xp5_ASAP7_75t_L g7741 ( 
.A(n_7735),
.B(n_7577),
.Y(n_7741)
);

OAI22xp33_ASAP7_75t_L g7742 ( 
.A1(n_7732),
.A2(n_7472),
.B1(n_7565),
.B2(n_7609),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7715),
.B(n_7306),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7720),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7740),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_7740),
.Y(n_7746)
);

INVxp67_ASAP7_75t_SL g7747 ( 
.A(n_7734),
.Y(n_7747)
);

NAND2xp33_ASAP7_75t_R g7748 ( 
.A(n_7725),
.B(n_7490),
.Y(n_7748)
);

OAI21xp5_ASAP7_75t_L g7749 ( 
.A1(n_7717),
.A2(n_7620),
.B(n_7674),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7714),
.Y(n_7750)
);

OAI321xp33_ASAP7_75t_L g7751 ( 
.A1(n_7719),
.A2(n_7739),
.A3(n_7713),
.B1(n_7557),
.B2(n_7563),
.C(n_7567),
.Y(n_7751)
);

AOI22xp5_ASAP7_75t_L g7752 ( 
.A1(n_7718),
.A2(n_7675),
.B1(n_7552),
.B2(n_7640),
.Y(n_7752)
);

AO21x1_ASAP7_75t_L g7753 ( 
.A1(n_7729),
.A2(n_7543),
.B(n_7540),
.Y(n_7753)
);

NOR2xp33_ASAP7_75t_L g7754 ( 
.A(n_7716),
.B(n_7394),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7730),
.Y(n_7755)
);

NOR2xp33_ASAP7_75t_L g7756 ( 
.A(n_7722),
.B(n_7369),
.Y(n_7756)
);

O2A1O1Ixp33_ASAP7_75t_L g7757 ( 
.A1(n_7729),
.A2(n_7617),
.B(n_7697),
.C(n_7506),
.Y(n_7757)
);

INVx2_ASAP7_75t_L g7758 ( 
.A(n_7736),
.Y(n_7758)
);

INVx2_ASAP7_75t_L g7759 ( 
.A(n_7736),
.Y(n_7759)
);

OAI21xp5_ASAP7_75t_L g7760 ( 
.A1(n_7724),
.A2(n_7456),
.B(n_7672),
.Y(n_7760)
);

AND2x2_ASAP7_75t_L g7761 ( 
.A(n_7727),
.B(n_7346),
.Y(n_7761)
);

NAND2xp5_ASAP7_75t_L g7762 ( 
.A(n_7726),
.B(n_7619),
.Y(n_7762)
);

AOI322xp5_ASAP7_75t_L g7763 ( 
.A1(n_7728),
.A2(n_7351),
.A3(n_7352),
.B1(n_7646),
.B2(n_7644),
.C1(n_7506),
.C2(n_7359),
.Y(n_7763)
);

NAND2x1p5_ASAP7_75t_L g7764 ( 
.A(n_7731),
.B(n_7654),
.Y(n_7764)
);

OAI22xp5_ASAP7_75t_L g7765 ( 
.A1(n_7721),
.A2(n_7645),
.B1(n_7655),
.B2(n_7607),
.Y(n_7765)
);

INVx2_ASAP7_75t_L g7766 ( 
.A(n_7733),
.Y(n_7766)
);

AOI22xp5_ASAP7_75t_L g7767 ( 
.A1(n_7723),
.A2(n_7322),
.B1(n_7711),
.B2(n_7353),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7737),
.Y(n_7768)
);

NOR2xp67_ASAP7_75t_L g7769 ( 
.A(n_7738),
.B(n_7546),
.Y(n_7769)
);

AOI21xp33_ASAP7_75t_L g7770 ( 
.A1(n_7735),
.A2(n_7629),
.B(n_7667),
.Y(n_7770)
);

AND3x1_ASAP7_75t_L g7771 ( 
.A(n_7713),
.B(n_7663),
.C(n_7678),
.Y(n_7771)
);

AOI22xp5_ASAP7_75t_L g7772 ( 
.A1(n_7718),
.A2(n_7364),
.B1(n_7362),
.B2(n_7354),
.Y(n_7772)
);

NAND2xp33_ASAP7_75t_L g7773 ( 
.A(n_7720),
.B(n_7485),
.Y(n_7773)
);

NAND2xp5_ASAP7_75t_L g7774 ( 
.A(n_7735),
.B(n_7628),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_7735),
.B(n_7376),
.Y(n_7775)
);

AOI311xp33_ASAP7_75t_L g7776 ( 
.A1(n_7770),
.A2(n_7649),
.A3(n_7668),
.B(n_7680),
.C(n_7679),
.Y(n_7776)
);

OAI221xp5_ASAP7_75t_SL g7777 ( 
.A1(n_7763),
.A2(n_7382),
.B1(n_7383),
.B2(n_7680),
.C(n_7668),
.Y(n_7777)
);

NOR2xp33_ASAP7_75t_L g7778 ( 
.A(n_7764),
.B(n_7384),
.Y(n_7778)
);

OAI32xp33_ASAP7_75t_L g7779 ( 
.A1(n_7762),
.A2(n_7397),
.A3(n_7387),
.B1(n_7392),
.B2(n_7390),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7753),
.Y(n_7780)
);

INVx1_ASAP7_75t_L g7781 ( 
.A(n_7747),
.Y(n_7781)
);

INVx3_ASAP7_75t_SL g7782 ( 
.A(n_7761),
.Y(n_7782)
);

NOR2xp33_ASAP7_75t_L g7783 ( 
.A(n_7742),
.B(n_7469),
.Y(n_7783)
);

OAI22xp5_ASAP7_75t_L g7784 ( 
.A1(n_7752),
.A2(n_7403),
.B1(n_7466),
.B2(n_7490),
.Y(n_7784)
);

A2O1A1Ixp33_ASAP7_75t_L g7785 ( 
.A1(n_7757),
.A2(n_7466),
.B(n_7490),
.C(n_513),
.Y(n_7785)
);

INVx1_ASAP7_75t_L g7786 ( 
.A(n_7769),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_7769),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7773),
.Y(n_7788)
);

OAI21xp5_ASAP7_75t_L g7789 ( 
.A1(n_7754),
.A2(n_510),
.B(n_512),
.Y(n_7789)
);

AND2x2_ASAP7_75t_L g7790 ( 
.A(n_7744),
.B(n_7758),
.Y(n_7790)
);

OAI22xp5_ASAP7_75t_L g7791 ( 
.A1(n_7772),
.A2(n_516),
.B1(n_513),
.B2(n_514),
.Y(n_7791)
);

OAI22xp5_ASAP7_75t_L g7792 ( 
.A1(n_7750),
.A2(n_519),
.B1(n_514),
.B2(n_516),
.Y(n_7792)
);

A2O1A1Ixp33_ASAP7_75t_L g7793 ( 
.A1(n_7756),
.A2(n_523),
.B(n_520),
.C(n_521),
.Y(n_7793)
);

AOI21xp5_ASAP7_75t_L g7794 ( 
.A1(n_7741),
.A2(n_521),
.B(n_523),
.Y(n_7794)
);

AOI21xp5_ASAP7_75t_L g7795 ( 
.A1(n_7765),
.A2(n_525),
.B(n_526),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7743),
.Y(n_7796)
);

OAI21xp33_ASAP7_75t_L g7797 ( 
.A1(n_7755),
.A2(n_525),
.B(n_526),
.Y(n_7797)
);

NAND4xp25_ASAP7_75t_L g7798 ( 
.A(n_7749),
.B(n_530),
.C(n_527),
.D(n_528),
.Y(n_7798)
);

OAI211xp5_ASAP7_75t_L g7799 ( 
.A1(n_7760),
.A2(n_531),
.B(n_527),
.C(n_530),
.Y(n_7799)
);

AO221x1_ASAP7_75t_L g7800 ( 
.A1(n_7745),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.C(n_536),
.Y(n_7800)
);

OAI221xp5_ASAP7_75t_L g7801 ( 
.A1(n_7748),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.C(n_537),
.Y(n_7801)
);

NAND2xp5_ASAP7_75t_SL g7802 ( 
.A(n_7759),
.B(n_3450),
.Y(n_7802)
);

OAI21xp5_ASAP7_75t_L g7803 ( 
.A1(n_7774),
.A2(n_538),
.B(n_539),
.Y(n_7803)
);

NAND2xp5_ASAP7_75t_SL g7804 ( 
.A(n_7751),
.B(n_3450),
.Y(n_7804)
);

INVx1_ASAP7_75t_SL g7805 ( 
.A(n_7775),
.Y(n_7805)
);

INVx1_ASAP7_75t_SL g7806 ( 
.A(n_7766),
.Y(n_7806)
);

O2A1O1Ixp33_ASAP7_75t_L g7807 ( 
.A1(n_7746),
.A2(n_538),
.B(n_539),
.C(n_542),
.Y(n_7807)
);

O2A1O1Ixp33_ASAP7_75t_L g7808 ( 
.A1(n_7768),
.A2(n_544),
.B(n_545),
.C(n_546),
.Y(n_7808)
);

AOI22xp33_ASAP7_75t_L g7809 ( 
.A1(n_7767),
.A2(n_3450),
.B1(n_548),
.B2(n_550),
.Y(n_7809)
);

AOI221xp5_ASAP7_75t_L g7810 ( 
.A1(n_7771),
.A2(n_545),
.B1(n_548),
.B2(n_550),
.C(n_551),
.Y(n_7810)
);

AOI211xp5_ASAP7_75t_L g7811 ( 
.A1(n_7779),
.A2(n_7784),
.B(n_7777),
.C(n_7783),
.Y(n_7811)
);

AOI21xp5_ASAP7_75t_L g7812 ( 
.A1(n_7778),
.A2(n_551),
.B(n_553),
.Y(n_7812)
);

A2O1A1Ixp33_ASAP7_75t_L g7813 ( 
.A1(n_7807),
.A2(n_553),
.B(n_554),
.C(n_555),
.Y(n_7813)
);

NAND2xp5_ASAP7_75t_L g7814 ( 
.A(n_7782),
.B(n_554),
.Y(n_7814)
);

OAI211xp5_ASAP7_75t_L g7815 ( 
.A1(n_7810),
.A2(n_555),
.B(n_556),
.C(n_557),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_7786),
.Y(n_7816)
);

AOI221x1_ASAP7_75t_L g7817 ( 
.A1(n_7780),
.A2(n_556),
.B1(n_558),
.B2(n_559),
.C(n_560),
.Y(n_7817)
);

NOR2xp33_ASAP7_75t_L g7818 ( 
.A(n_7798),
.B(n_558),
.Y(n_7818)
);

NOR3xp33_ASAP7_75t_L g7819 ( 
.A(n_7781),
.B(n_560),
.C(n_561),
.Y(n_7819)
);

OAI22xp5_ASAP7_75t_L g7820 ( 
.A1(n_7806),
.A2(n_561),
.B1(n_562),
.B2(n_564),
.Y(n_7820)
);

AOI21xp5_ASAP7_75t_L g7821 ( 
.A1(n_7787),
.A2(n_562),
.B(n_564),
.Y(n_7821)
);

OAI21xp33_ASAP7_75t_SL g7822 ( 
.A1(n_7804),
.A2(n_565),
.B(n_566),
.Y(n_7822)
);

OAI221xp5_ASAP7_75t_L g7823 ( 
.A1(n_7785),
.A2(n_566),
.B1(n_567),
.B2(n_570),
.C(n_571),
.Y(n_7823)
);

OAI211xp5_ASAP7_75t_L g7824 ( 
.A1(n_7799),
.A2(n_567),
.B(n_570),
.C(n_571),
.Y(n_7824)
);

OAI211xp5_ASAP7_75t_SL g7825 ( 
.A1(n_7788),
.A2(n_572),
.B(n_573),
.C(n_574),
.Y(n_7825)
);

AOI221xp5_ASAP7_75t_L g7826 ( 
.A1(n_7801),
.A2(n_575),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_7826)
);

AOI211xp5_ASAP7_75t_L g7827 ( 
.A1(n_7795),
.A2(n_577),
.B(n_580),
.C(n_581),
.Y(n_7827)
);

O2A1O1Ixp5_ASAP7_75t_L g7828 ( 
.A1(n_7802),
.A2(n_581),
.B(n_582),
.C(n_583),
.Y(n_7828)
);

AND2x2_ASAP7_75t_L g7829 ( 
.A(n_7790),
.B(n_584),
.Y(n_7829)
);

OAI21xp5_ASAP7_75t_L g7830 ( 
.A1(n_7805),
.A2(n_584),
.B(n_585),
.Y(n_7830)
);

OAI21xp33_ASAP7_75t_L g7831 ( 
.A1(n_7796),
.A2(n_587),
.B(n_588),
.Y(n_7831)
);

NOR3xp33_ASAP7_75t_SL g7832 ( 
.A(n_7791),
.B(n_589),
.C(n_590),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7800),
.Y(n_7833)
);

AOI22xp5_ASAP7_75t_L g7834 ( 
.A1(n_7797),
.A2(n_7809),
.B1(n_7789),
.B2(n_7794),
.Y(n_7834)
);

AOI322xp5_ASAP7_75t_L g7835 ( 
.A1(n_7776),
.A2(n_589),
.A3(n_591),
.B1(n_592),
.B2(n_595),
.C1(n_596),
.C2(n_597),
.Y(n_7835)
);

AOI21xp33_ASAP7_75t_L g7836 ( 
.A1(n_7808),
.A2(n_592),
.B(n_598),
.Y(n_7836)
);

NOR3xp33_ASAP7_75t_L g7837 ( 
.A(n_7803),
.B(n_598),
.C(n_599),
.Y(n_7837)
);

AOI21xp5_ASAP7_75t_L g7838 ( 
.A1(n_7793),
.A2(n_600),
.B(n_601),
.Y(n_7838)
);

AND2x2_ASAP7_75t_L g7839 ( 
.A(n_7792),
.B(n_600),
.Y(n_7839)
);

AOI22xp33_ASAP7_75t_L g7840 ( 
.A1(n_7781),
.A2(n_3450),
.B1(n_602),
.B2(n_603),
.Y(n_7840)
);

INVxp67_ASAP7_75t_L g7841 ( 
.A(n_7783),
.Y(n_7841)
);

OAI211xp5_ASAP7_75t_SL g7842 ( 
.A1(n_7781),
.A2(n_601),
.B(n_603),
.C(n_604),
.Y(n_7842)
);

AOI22xp5_ASAP7_75t_L g7843 ( 
.A1(n_7778),
.A2(n_3450),
.B1(n_606),
.B2(n_607),
.Y(n_7843)
);

AOI22xp5_ASAP7_75t_L g7844 ( 
.A1(n_7778),
.A2(n_605),
.B1(n_608),
.B2(n_609),
.Y(n_7844)
);

NAND2xp5_ASAP7_75t_L g7845 ( 
.A(n_7829),
.B(n_608),
.Y(n_7845)
);

O2A1O1Ixp33_ASAP7_75t_L g7846 ( 
.A1(n_7813),
.A2(n_609),
.B(n_610),
.C(n_611),
.Y(n_7846)
);

NAND3xp33_ASAP7_75t_L g7847 ( 
.A(n_7835),
.B(n_612),
.C(n_613),
.Y(n_7847)
);

NOR4xp25_ASAP7_75t_L g7848 ( 
.A(n_7833),
.B(n_613),
.C(n_614),
.D(n_616),
.Y(n_7848)
);

OAI21xp5_ASAP7_75t_SL g7849 ( 
.A1(n_7841),
.A2(n_616),
.B(n_617),
.Y(n_7849)
);

AOI21xp33_ASAP7_75t_L g7850 ( 
.A1(n_7816),
.A2(n_618),
.B(n_620),
.Y(n_7850)
);

NOR3xp33_ASAP7_75t_L g7851 ( 
.A(n_7811),
.B(n_618),
.C(n_620),
.Y(n_7851)
);

INVx2_ASAP7_75t_L g7852 ( 
.A(n_7828),
.Y(n_7852)
);

NAND2x1_ASAP7_75t_L g7853 ( 
.A(n_7832),
.B(n_621),
.Y(n_7853)
);

OAI221xp5_ASAP7_75t_L g7854 ( 
.A1(n_7823),
.A2(n_622),
.B1(n_623),
.B2(n_624),
.C(n_626),
.Y(n_7854)
);

OAI211xp5_ASAP7_75t_L g7855 ( 
.A1(n_7817),
.A2(n_622),
.B(n_623),
.C(n_624),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7814),
.Y(n_7856)
);

AOI221xp5_ASAP7_75t_L g7857 ( 
.A1(n_7836),
.A2(n_626),
.B1(n_627),
.B2(n_628),
.C(n_629),
.Y(n_7857)
);

AOI22xp5_ASAP7_75t_L g7858 ( 
.A1(n_7818),
.A2(n_628),
.B1(n_629),
.B2(n_631),
.Y(n_7858)
);

NAND3xp33_ASAP7_75t_L g7859 ( 
.A(n_7827),
.B(n_632),
.C(n_633),
.Y(n_7859)
);

INVx2_ASAP7_75t_L g7860 ( 
.A(n_7839),
.Y(n_7860)
);

O2A1O1Ixp33_ASAP7_75t_L g7861 ( 
.A1(n_7822),
.A2(n_632),
.B(n_633),
.C(n_634),
.Y(n_7861)
);

NAND3xp33_ASAP7_75t_SL g7862 ( 
.A(n_7826),
.B(n_634),
.C(n_636),
.Y(n_7862)
);

OAI21xp33_ASAP7_75t_L g7863 ( 
.A1(n_7834),
.A2(n_638),
.B(n_639),
.Y(n_7863)
);

NAND4xp25_ASAP7_75t_L g7864 ( 
.A(n_7837),
.B(n_639),
.C(n_640),
.D(n_642),
.Y(n_7864)
);

AOI221xp5_ASAP7_75t_L g7865 ( 
.A1(n_7824),
.A2(n_640),
.B1(n_644),
.B2(n_645),
.C(n_646),
.Y(n_7865)
);

O2A1O1Ixp33_ASAP7_75t_L g7866 ( 
.A1(n_7830),
.A2(n_644),
.B(n_647),
.C(n_648),
.Y(n_7866)
);

NOR3xp33_ASAP7_75t_L g7867 ( 
.A(n_7815),
.B(n_7825),
.C(n_7842),
.Y(n_7867)
);

AOI21xp33_ASAP7_75t_L g7868 ( 
.A1(n_7838),
.A2(n_648),
.B(n_649),
.Y(n_7868)
);

NAND3xp33_ASAP7_75t_L g7869 ( 
.A(n_7812),
.B(n_7819),
.C(n_7821),
.Y(n_7869)
);

AOI211xp5_ASAP7_75t_L g7870 ( 
.A1(n_7831),
.A2(n_650),
.B(n_652),
.C(n_653),
.Y(n_7870)
);

AOI221xp5_ASAP7_75t_L g7871 ( 
.A1(n_7820),
.A2(n_7840),
.B1(n_7843),
.B2(n_7844),
.C(n_656),
.Y(n_7871)
);

NAND4xp25_ASAP7_75t_L g7872 ( 
.A(n_7811),
.B(n_652),
.C(n_653),
.D(n_655),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_7845),
.Y(n_7873)
);

NOR3xp33_ASAP7_75t_L g7874 ( 
.A(n_7872),
.B(n_656),
.C(n_658),
.Y(n_7874)
);

AND2x2_ASAP7_75t_L g7875 ( 
.A(n_7848),
.B(n_658),
.Y(n_7875)
);

NAND2xp5_ASAP7_75t_SL g7876 ( 
.A(n_7865),
.B(n_660),
.Y(n_7876)
);

AOI22xp5_ASAP7_75t_L g7877 ( 
.A1(n_7851),
.A2(n_660),
.B1(n_662),
.B2(n_663),
.Y(n_7877)
);

NOR2xp33_ASAP7_75t_L g7878 ( 
.A(n_7864),
.B(n_662),
.Y(n_7878)
);

NAND3xp33_ASAP7_75t_L g7879 ( 
.A(n_7857),
.B(n_663),
.C(n_664),
.Y(n_7879)
);

NAND4xp25_ASAP7_75t_SL g7880 ( 
.A(n_7866),
.B(n_664),
.C(n_665),
.D(n_666),
.Y(n_7880)
);

NOR2x1_ASAP7_75t_L g7881 ( 
.A(n_7855),
.B(n_7849),
.Y(n_7881)
);

INVx2_ASAP7_75t_L g7882 ( 
.A(n_7853),
.Y(n_7882)
);

NAND2xp5_ASAP7_75t_L g7883 ( 
.A(n_7863),
.B(n_666),
.Y(n_7883)
);

NOR2xp33_ASAP7_75t_L g7884 ( 
.A(n_7847),
.B(n_667),
.Y(n_7884)
);

INVx1_ASAP7_75t_L g7885 ( 
.A(n_7861),
.Y(n_7885)
);

AOI211xp5_ASAP7_75t_SL g7886 ( 
.A1(n_7868),
.A2(n_667),
.B(n_668),
.C(n_669),
.Y(n_7886)
);

NAND4xp25_ASAP7_75t_L g7887 ( 
.A(n_7867),
.B(n_668),
.C(n_669),
.D(n_672),
.Y(n_7887)
);

NAND2xp5_ASAP7_75t_L g7888 ( 
.A(n_7870),
.B(n_672),
.Y(n_7888)
);

NOR2xp67_ASAP7_75t_L g7889 ( 
.A(n_7859),
.B(n_673),
.Y(n_7889)
);

AND3x1_ASAP7_75t_L g7890 ( 
.A(n_7852),
.B(n_673),
.C(n_674),
.Y(n_7890)
);

NOR4xp25_ASAP7_75t_L g7891 ( 
.A(n_7862),
.B(n_674),
.C(n_675),
.D(n_676),
.Y(n_7891)
);

NAND2xp5_ASAP7_75t_L g7892 ( 
.A(n_7858),
.B(n_675),
.Y(n_7892)
);

NOR2xp33_ASAP7_75t_L g7893 ( 
.A(n_7854),
.B(n_678),
.Y(n_7893)
);

NAND2xp5_ASAP7_75t_SL g7894 ( 
.A(n_7871),
.B(n_679),
.Y(n_7894)
);

INVx1_ASAP7_75t_L g7895 ( 
.A(n_7846),
.Y(n_7895)
);

NAND3x1_ASAP7_75t_L g7896 ( 
.A(n_7856),
.B(n_680),
.C(n_681),
.Y(n_7896)
);

NAND2xp5_ASAP7_75t_L g7897 ( 
.A(n_7850),
.B(n_680),
.Y(n_7897)
);

NAND3xp33_ASAP7_75t_L g7898 ( 
.A(n_7886),
.B(n_7869),
.C(n_7860),
.Y(n_7898)
);

NAND4xp25_ASAP7_75t_L g7899 ( 
.A(n_7874),
.B(n_681),
.C(n_682),
.D(n_683),
.Y(n_7899)
);

NOR3xp33_ASAP7_75t_L g7900 ( 
.A(n_7894),
.B(n_7885),
.C(n_7882),
.Y(n_7900)
);

NOR2x1_ASAP7_75t_L g7901 ( 
.A(n_7887),
.B(n_682),
.Y(n_7901)
);

AND4x2_ASAP7_75t_L g7902 ( 
.A(n_7881),
.B(n_7891),
.C(n_7880),
.D(n_7890),
.Y(n_7902)
);

NAND4xp25_ASAP7_75t_L g7903 ( 
.A(n_7878),
.B(n_684),
.C(n_685),
.D(n_687),
.Y(n_7903)
);

NAND2xp5_ASAP7_75t_L g7904 ( 
.A(n_7875),
.B(n_688),
.Y(n_7904)
);

AOI211xp5_ASAP7_75t_L g7905 ( 
.A1(n_7884),
.A2(n_691),
.B(n_694),
.C(n_695),
.Y(n_7905)
);

NOR2x1_ASAP7_75t_L g7906 ( 
.A(n_7897),
.B(n_696),
.Y(n_7906)
);

AOI221xp5_ASAP7_75t_L g7907 ( 
.A1(n_7893),
.A2(n_698),
.B1(n_700),
.B2(n_701),
.C(n_702),
.Y(n_7907)
);

AND2x4_ASAP7_75t_L g7908 ( 
.A(n_7889),
.B(n_700),
.Y(n_7908)
);

NOR2xp67_ASAP7_75t_L g7909 ( 
.A(n_7877),
.B(n_703),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7896),
.Y(n_7910)
);

NOR3x1_ASAP7_75t_SL g7911 ( 
.A(n_7873),
.B(n_703),
.C(n_704),
.Y(n_7911)
);

AOI211x1_ASAP7_75t_L g7912 ( 
.A1(n_7879),
.A2(n_704),
.B(n_705),
.C(n_706),
.Y(n_7912)
);

OAI211xp5_ASAP7_75t_L g7913 ( 
.A1(n_7883),
.A2(n_706),
.B(n_2673),
.C(n_2674),
.Y(n_7913)
);

AOI211xp5_ASAP7_75t_SL g7914 ( 
.A1(n_7895),
.A2(n_7888),
.B(n_7892),
.C(n_7876),
.Y(n_7914)
);

AOI21xp33_ASAP7_75t_SL g7915 ( 
.A1(n_7884),
.A2(n_1323),
.B(n_2572),
.Y(n_7915)
);

NOR3xp33_ASAP7_75t_L g7916 ( 
.A(n_7894),
.B(n_2269),
.C(n_2198),
.Y(n_7916)
);

NOR3xp33_ASAP7_75t_L g7917 ( 
.A(n_7894),
.B(n_2269),
.C(n_2198),
.Y(n_7917)
);

NAND4xp25_ASAP7_75t_L g7918 ( 
.A(n_7874),
.B(n_2352),
.C(n_2397),
.D(n_2269),
.Y(n_7918)
);

NOR3xp33_ASAP7_75t_L g7919 ( 
.A(n_7894),
.B(n_1323),
.C(n_2572),
.Y(n_7919)
);

AND2x2_ASAP7_75t_L g7920 ( 
.A(n_7875),
.B(n_2356),
.Y(n_7920)
);

NAND4xp75_ASAP7_75t_L g7921 ( 
.A(n_7890),
.B(n_2572),
.C(n_2899),
.D(n_3338),
.Y(n_7921)
);

NAND2xp5_ASAP7_75t_L g7922 ( 
.A(n_7875),
.B(n_2350),
.Y(n_7922)
);

NOR2xp33_ASAP7_75t_L g7923 ( 
.A(n_7880),
.B(n_2572),
.Y(n_7923)
);

NAND3xp33_ASAP7_75t_SL g7924 ( 
.A(n_7891),
.B(n_2718),
.C(n_2674),
.Y(n_7924)
);

NAND2xp5_ASAP7_75t_L g7925 ( 
.A(n_7875),
.B(n_2350),
.Y(n_7925)
);

NOR2x1_ASAP7_75t_L g7926 ( 
.A(n_7887),
.B(n_2350),
.Y(n_7926)
);

NAND3xp33_ASAP7_75t_L g7927 ( 
.A(n_7886),
.B(n_2674),
.C(n_2710),
.Y(n_7927)
);

AND2x2_ASAP7_75t_L g7928 ( 
.A(n_7901),
.B(n_7908),
.Y(n_7928)
);

INVx1_ASAP7_75t_SL g7929 ( 
.A(n_7904),
.Y(n_7929)
);

INVx4_ASAP7_75t_L g7930 ( 
.A(n_7908),
.Y(n_7930)
);

INVx2_ASAP7_75t_SL g7931 ( 
.A(n_7910),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7911),
.Y(n_7932)
);

AND2x2_ASAP7_75t_L g7933 ( 
.A(n_7906),
.B(n_2350),
.Y(n_7933)
);

NAND2xp5_ASAP7_75t_L g7934 ( 
.A(n_7905),
.B(n_2350),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_7902),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_7912),
.Y(n_7936)
);

NAND2xp5_ASAP7_75t_SL g7937 ( 
.A(n_7907),
.B(n_2674),
.Y(n_7937)
);

AND2x2_ASAP7_75t_L g7938 ( 
.A(n_7909),
.B(n_2342),
.Y(n_7938)
);

OAI221xp5_ASAP7_75t_L g7939 ( 
.A1(n_7899),
.A2(n_2732),
.B1(n_2726),
.B2(n_2718),
.C(n_2710),
.Y(n_7939)
);

NOR2xp33_ASAP7_75t_L g7940 ( 
.A(n_7903),
.B(n_2673),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_7920),
.Y(n_7941)
);

AOI21xp5_ASAP7_75t_L g7942 ( 
.A1(n_7922),
.A2(n_2342),
.B(n_2356),
.Y(n_7942)
);

INVx2_ASAP7_75t_SL g7943 ( 
.A(n_7926),
.Y(n_7943)
);

NAND2xp5_ASAP7_75t_L g7944 ( 
.A(n_7923),
.B(n_2342),
.Y(n_7944)
);

NAND2xp5_ASAP7_75t_L g7945 ( 
.A(n_7914),
.B(n_2342),
.Y(n_7945)
);

INVx1_ASAP7_75t_L g7946 ( 
.A(n_7925),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7921),
.Y(n_7947)
);

AND2x2_ASAP7_75t_L g7948 ( 
.A(n_7900),
.B(n_2342),
.Y(n_7948)
);

INVxp67_ASAP7_75t_L g7949 ( 
.A(n_7898),
.Y(n_7949)
);

INVx1_ASAP7_75t_L g7950 ( 
.A(n_7924),
.Y(n_7950)
);

NOR2x1_ASAP7_75t_L g7951 ( 
.A(n_7927),
.B(n_2356),
.Y(n_7951)
);

NAND2xp5_ASAP7_75t_L g7952 ( 
.A(n_7913),
.B(n_2356),
.Y(n_7952)
);

NAND2xp5_ASAP7_75t_L g7953 ( 
.A(n_7932),
.B(n_7917),
.Y(n_7953)
);

OAI22xp5_ASAP7_75t_L g7954 ( 
.A1(n_7949),
.A2(n_7915),
.B1(n_7916),
.B2(n_7919),
.Y(n_7954)
);

NOR2xp33_ASAP7_75t_L g7955 ( 
.A(n_7930),
.B(n_7918),
.Y(n_7955)
);

NOR2x1_ASAP7_75t_L g7956 ( 
.A(n_7930),
.B(n_2356),
.Y(n_7956)
);

OAI211xp5_ASAP7_75t_L g7957 ( 
.A1(n_7935),
.A2(n_2325),
.B(n_2293),
.C(n_2290),
.Y(n_7957)
);

NOR4xp75_ASAP7_75t_L g7958 ( 
.A(n_7931),
.B(n_2325),
.C(n_2288),
.D(n_2286),
.Y(n_7958)
);

NOR3x1_ASAP7_75t_L g7959 ( 
.A(n_7936),
.B(n_2325),
.C(n_2317),
.Y(n_7959)
);

NAND4xp25_ASAP7_75t_L g7960 ( 
.A(n_7929),
.B(n_2325),
.C(n_2317),
.D(n_2316),
.Y(n_7960)
);

NAND4xp25_ASAP7_75t_L g7961 ( 
.A(n_7940),
.B(n_7928),
.C(n_7952),
.D(n_7945),
.Y(n_7961)
);

OR2x2_ASAP7_75t_L g7962 ( 
.A(n_7934),
.B(n_7941),
.Y(n_7962)
);

NOR3xp33_ASAP7_75t_L g7963 ( 
.A(n_7946),
.B(n_2325),
.C(n_2286),
.Y(n_7963)
);

INVxp33_ASAP7_75t_SL g7964 ( 
.A(n_7948),
.Y(n_7964)
);

AND2x4_ASAP7_75t_L g7965 ( 
.A(n_7933),
.B(n_2673),
.Y(n_7965)
);

NOR3x1_ASAP7_75t_L g7966 ( 
.A(n_7947),
.B(n_2290),
.C(n_2317),
.Y(n_7966)
);

AOI211xp5_ASAP7_75t_L g7967 ( 
.A1(n_7937),
.A2(n_2726),
.B(n_2673),
.C(n_2674),
.Y(n_7967)
);

NAND4xp75_ASAP7_75t_L g7968 ( 
.A(n_7951),
.B(n_2317),
.C(n_2316),
.D(n_2314),
.Y(n_7968)
);

NAND4xp75_ASAP7_75t_L g7969 ( 
.A(n_7950),
.B(n_2317),
.C(n_2316),
.D(n_2314),
.Y(n_7969)
);

INVx1_ASAP7_75t_L g7970 ( 
.A(n_7938),
.Y(n_7970)
);

INVx1_ASAP7_75t_SL g7971 ( 
.A(n_7962),
.Y(n_7971)
);

NAND2xp5_ASAP7_75t_SL g7972 ( 
.A(n_7953),
.B(n_7964),
.Y(n_7972)
);

AOI22xp5_ASAP7_75t_L g7973 ( 
.A1(n_7955),
.A2(n_7943),
.B1(n_7944),
.B2(n_7939),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_7965),
.Y(n_7974)
);

AOI22xp5_ASAP7_75t_L g7975 ( 
.A1(n_7961),
.A2(n_7942),
.B1(n_2732),
.B2(n_2718),
.Y(n_7975)
);

INVx2_ASAP7_75t_L g7976 ( 
.A(n_7965),
.Y(n_7976)
);

INVx2_ASAP7_75t_L g7977 ( 
.A(n_7966),
.Y(n_7977)
);

NOR4xp75_ASAP7_75t_L g7978 ( 
.A(n_7972),
.B(n_7954),
.C(n_7968),
.D(n_7969),
.Y(n_7978)
);

NOR2xp33_ASAP7_75t_L g7979 ( 
.A(n_7971),
.B(n_7970),
.Y(n_7979)
);

NOR2xp33_ASAP7_75t_L g7980 ( 
.A(n_7976),
.B(n_7956),
.Y(n_7980)
);

AOI221xp5_ASAP7_75t_L g7981 ( 
.A1(n_7974),
.A2(n_7960),
.B1(n_7963),
.B2(n_7967),
.C(n_7957),
.Y(n_7981)
);

OAI211xp5_ASAP7_75t_L g7982 ( 
.A1(n_7973),
.A2(n_7958),
.B(n_7959),
.C(n_2316),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_L g7983 ( 
.A(n_7979),
.B(n_7977),
.Y(n_7983)
);

OAI321xp33_ASAP7_75t_L g7984 ( 
.A1(n_7980),
.A2(n_7975),
.A3(n_2732),
.B1(n_2726),
.B2(n_2718),
.C(n_2710),
.Y(n_7984)
);

OR2x2_ASAP7_75t_L g7985 ( 
.A(n_7982),
.B(n_2298),
.Y(n_7985)
);

INVx1_ASAP7_75t_L g7986 ( 
.A(n_7978),
.Y(n_7986)
);

NAND3x1_ASAP7_75t_L g7987 ( 
.A(n_7981),
.B(n_2316),
.C(n_2286),
.Y(n_7987)
);

INVx1_ASAP7_75t_L g7988 ( 
.A(n_7979),
.Y(n_7988)
);

OR2x2_ASAP7_75t_L g7989 ( 
.A(n_7979),
.B(n_2297),
.Y(n_7989)
);

NAND4xp75_ASAP7_75t_L g7990 ( 
.A(n_7979),
.B(n_2293),
.C(n_2290),
.D(n_2288),
.Y(n_7990)
);

AOI221xp5_ASAP7_75t_L g7991 ( 
.A1(n_7979),
.A2(n_2673),
.B1(n_2705),
.B2(n_2710),
.C(n_2718),
.Y(n_7991)
);

AOI221x1_ASAP7_75t_L g7992 ( 
.A1(n_7979),
.A2(n_2314),
.B1(n_2298),
.B2(n_2297),
.C(n_2293),
.Y(n_7992)
);

XNOR2x1_ASAP7_75t_L g7993 ( 
.A(n_7988),
.B(n_2314),
.Y(n_7993)
);

INVx2_ASAP7_75t_L g7994 ( 
.A(n_7989),
.Y(n_7994)
);

OAI22x1_ASAP7_75t_SL g7995 ( 
.A1(n_7986),
.A2(n_2143),
.B1(n_2128),
.B2(n_2298),
.Y(n_7995)
);

INVx2_ASAP7_75t_SL g7996 ( 
.A(n_7983),
.Y(n_7996)
);

INVx2_ASAP7_75t_SL g7997 ( 
.A(n_7985),
.Y(n_7997)
);

INVx1_ASAP7_75t_L g7998 ( 
.A(n_7987),
.Y(n_7998)
);

O2A1O1Ixp33_ASAP7_75t_SL g7999 ( 
.A1(n_7984),
.A2(n_2314),
.B(n_2298),
.C(n_2297),
.Y(n_7999)
);

AND2x2_ASAP7_75t_L g8000 ( 
.A(n_7990),
.B(n_2293),
.Y(n_8000)
);

INVx3_ASAP7_75t_L g8001 ( 
.A(n_7991),
.Y(n_8001)
);

INVx2_ASAP7_75t_L g8002 ( 
.A(n_7992),
.Y(n_8002)
);

INVx2_ASAP7_75t_SL g8003 ( 
.A(n_7988),
.Y(n_8003)
);

INVx1_ASAP7_75t_L g8004 ( 
.A(n_7989),
.Y(n_8004)
);

OAI21xp5_ASAP7_75t_L g8005 ( 
.A1(n_7988),
.A2(n_2143),
.B(n_2128),
.Y(n_8005)
);

NAND3x1_ASAP7_75t_L g8006 ( 
.A(n_7983),
.B(n_2286),
.C(n_2288),
.Y(n_8006)
);

AOI322xp5_ASAP7_75t_L g8007 ( 
.A1(n_7996),
.A2(n_2937),
.A3(n_2930),
.B1(n_2928),
.B2(n_2927),
.C1(n_2969),
.C2(n_2924),
.Y(n_8007)
);

NAND3xp33_ASAP7_75t_L g8008 ( 
.A(n_8003),
.B(n_2290),
.C(n_2293),
.Y(n_8008)
);

AOI322xp5_ASAP7_75t_L g8009 ( 
.A1(n_7997),
.A2(n_2937),
.A3(n_2930),
.B1(n_2928),
.B2(n_2927),
.C1(n_2969),
.C2(n_2924),
.Y(n_8009)
);

AOI22xp5_ASAP7_75t_L g8010 ( 
.A1(n_8004),
.A2(n_2732),
.B1(n_2726),
.B2(n_2710),
.Y(n_8010)
);

AND2x4_ASAP7_75t_L g8011 ( 
.A(n_7994),
.B(n_8000),
.Y(n_8011)
);

INVx2_ASAP7_75t_L g8012 ( 
.A(n_7993),
.Y(n_8012)
);

OAI22xp5_ASAP7_75t_L g8013 ( 
.A1(n_8006),
.A2(n_2732),
.B1(n_2726),
.B2(n_2705),
.Y(n_8013)
);

OAI22xp5_ASAP7_75t_L g8014 ( 
.A1(n_8012),
.A2(n_8001),
.B1(n_7998),
.B2(n_8002),
.Y(n_8014)
);

OAI21xp5_ASAP7_75t_L g8015 ( 
.A1(n_8011),
.A2(n_8005),
.B(n_7999),
.Y(n_8015)
);

OAI21xp5_ASAP7_75t_SL g8016 ( 
.A1(n_8008),
.A2(n_7995),
.B(n_2298),
.Y(n_8016)
);

AND3x1_ASAP7_75t_L g8017 ( 
.A(n_8010),
.B(n_2297),
.C(n_2290),
.Y(n_8017)
);

NOR2xp67_ASAP7_75t_L g8018 ( 
.A(n_8013),
.B(n_2297),
.Y(n_8018)
);

INVx2_ASAP7_75t_L g8019 ( 
.A(n_8017),
.Y(n_8019)
);

OR2x2_ASAP7_75t_L g8020 ( 
.A(n_8014),
.B(n_8007),
.Y(n_8020)
);

INVx4_ASAP7_75t_L g8021 ( 
.A(n_8015),
.Y(n_8021)
);

AOI22xp5_ASAP7_75t_L g8022 ( 
.A1(n_8018),
.A2(n_8009),
.B1(n_2193),
.B2(n_2192),
.Y(n_8022)
);

NOR2xp33_ASAP7_75t_SL g8023 ( 
.A(n_8016),
.B(n_2096),
.Y(n_8023)
);

CKINVDCx5p33_ASAP7_75t_R g8024 ( 
.A(n_8014),
.Y(n_8024)
);

BUFx2_ASAP7_75t_SL g8025 ( 
.A(n_8014),
.Y(n_8025)
);

XNOR2x1_ASAP7_75t_L g8026 ( 
.A(n_8014),
.B(n_2404),
.Y(n_8026)
);

OR2x2_ASAP7_75t_L g8027 ( 
.A(n_8014),
.B(n_2705),
.Y(n_8027)
);

INVx3_ASAP7_75t_L g8028 ( 
.A(n_8017),
.Y(n_8028)
);

NAND2xp5_ASAP7_75t_L g8029 ( 
.A(n_8014),
.B(n_2404),
.Y(n_8029)
);

INVx2_ASAP7_75t_L g8030 ( 
.A(n_8017),
.Y(n_8030)
);

XNOR2xp5_ASAP7_75t_L g8031 ( 
.A(n_8014),
.B(n_2404),
.Y(n_8031)
);

AOI22xp5_ASAP7_75t_L g8032 ( 
.A1(n_8014),
.A2(n_2193),
.B1(n_2192),
.B2(n_2187),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_8025),
.Y(n_8033)
);

AOI21x1_ASAP7_75t_L g8034 ( 
.A1(n_8026),
.A2(n_2404),
.B(n_2368),
.Y(n_8034)
);

AO21x1_ASAP7_75t_L g8035 ( 
.A1(n_8021),
.A2(n_2404),
.B(n_2368),
.Y(n_8035)
);

OAI22x1_ASAP7_75t_L g8036 ( 
.A1(n_8024),
.A2(n_8031),
.B1(n_8027),
.B2(n_8020),
.Y(n_8036)
);

OR2x2_ASAP7_75t_L g8037 ( 
.A(n_8029),
.B(n_2705),
.Y(n_8037)
);

OAI22x1_ASAP7_75t_L g8038 ( 
.A1(n_8019),
.A2(n_2143),
.B1(n_2128),
.B2(n_2105),
.Y(n_8038)
);

INVx1_ASAP7_75t_L g8039 ( 
.A(n_8030),
.Y(n_8039)
);

AOI22xp33_ASAP7_75t_L g8040 ( 
.A1(n_8028),
.A2(n_2096),
.B1(n_2101),
.B2(n_2105),
.Y(n_8040)
);

NAND3xp33_ASAP7_75t_L g8041 ( 
.A(n_8023),
.B(n_2193),
.C(n_2192),
.Y(n_8041)
);

INVx2_ASAP7_75t_L g8042 ( 
.A(n_8037),
.Y(n_8042)
);

OAI22xp5_ASAP7_75t_L g8043 ( 
.A1(n_8033),
.A2(n_8022),
.B1(n_8032),
.B2(n_2105),
.Y(n_8043)
);

AOI311xp33_ASAP7_75t_L g8044 ( 
.A1(n_8039),
.A2(n_2096),
.A3(n_2101),
.B(n_2105),
.C(n_2117),
.Y(n_8044)
);

O2A1O1Ixp33_ASAP7_75t_L g8045 ( 
.A1(n_8035),
.A2(n_2368),
.B(n_2193),
.C(n_2192),
.Y(n_8045)
);

AND2x2_ASAP7_75t_L g8046 ( 
.A(n_8036),
.B(n_2368),
.Y(n_8046)
);

OA22x2_ASAP7_75t_L g8047 ( 
.A1(n_8038),
.A2(n_2193),
.B1(n_2192),
.B2(n_2187),
.Y(n_8047)
);

OAI22xp5_ASAP7_75t_L g8048 ( 
.A1(n_8041),
.A2(n_8034),
.B1(n_8040),
.B2(n_2105),
.Y(n_8048)
);

AOI21xp5_ASAP7_75t_L g8049 ( 
.A1(n_8042),
.A2(n_2368),
.B(n_2187),
.Y(n_8049)
);

XNOR2xp5_ASAP7_75t_L g8050 ( 
.A(n_8046),
.B(n_2096),
.Y(n_8050)
);

OAI21xp5_ASAP7_75t_L g8051 ( 
.A1(n_8043),
.A2(n_2128),
.B(n_2143),
.Y(n_8051)
);

BUFx2_ASAP7_75t_L g8052 ( 
.A(n_8048),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_8050),
.Y(n_8053)
);

OAI22xp5_ASAP7_75t_L g8054 ( 
.A1(n_8052),
.A2(n_8047),
.B1(n_8045),
.B2(n_8044),
.Y(n_8054)
);

OAI21xp33_ASAP7_75t_L g8055 ( 
.A1(n_8051),
.A2(n_2096),
.B(n_2101),
.Y(n_8055)
);

OAI22xp5_ASAP7_75t_L g8056 ( 
.A1(n_8053),
.A2(n_8049),
.B1(n_2117),
.B2(n_2101),
.Y(n_8056)
);

NAND2xp5_ASAP7_75t_L g8057 ( 
.A(n_8054),
.B(n_2187),
.Y(n_8057)
);

OAI22xp33_ASAP7_75t_L g8058 ( 
.A1(n_8057),
.A2(n_8055),
.B1(n_2117),
.B2(n_2101),
.Y(n_8058)
);

AOI22xp33_ASAP7_75t_L g8059 ( 
.A1(n_8056),
.A2(n_2117),
.B1(n_2130),
.B2(n_2136),
.Y(n_8059)
);

NAND2xp5_ASAP7_75t_L g8060 ( 
.A(n_8058),
.B(n_2187),
.Y(n_8060)
);

AND2x2_ASAP7_75t_L g8061 ( 
.A(n_8059),
.B(n_2705),
.Y(n_8061)
);

OR2x2_ASAP7_75t_L g8062 ( 
.A(n_8058),
.B(n_2117),
.Y(n_8062)
);

INVx1_ASAP7_75t_L g8063 ( 
.A(n_8062),
.Y(n_8063)
);

XNOR2xp5_ASAP7_75t_L g8064 ( 
.A(n_8060),
.B(n_2264),
.Y(n_8064)
);

BUFx2_ASAP7_75t_L g8065 ( 
.A(n_8061),
.Y(n_8065)
);

AO21x2_ASAP7_75t_L g8066 ( 
.A1(n_8063),
.A2(n_2128),
.B(n_2143),
.Y(n_8066)
);

AOI221xp5_ASAP7_75t_L g8067 ( 
.A1(n_8065),
.A2(n_2275),
.B1(n_2130),
.B2(n_2136),
.C(n_2143),
.Y(n_8067)
);

NAND2xp5_ASAP7_75t_L g8068 ( 
.A(n_8064),
.B(n_2130),
.Y(n_8068)
);

AOI221xp5_ASAP7_75t_L g8069 ( 
.A1(n_8068),
.A2(n_2275),
.B1(n_2130),
.B2(n_2136),
.C(n_2128),
.Y(n_8069)
);

AOI221xp5_ASAP7_75t_L g8070 ( 
.A1(n_8066),
.A2(n_2275),
.B1(n_2130),
.B2(n_2136),
.C(n_2901),
.Y(n_8070)
);

AOI22xp33_ASAP7_75t_SL g8071 ( 
.A1(n_8070),
.A2(n_8069),
.B1(n_8067),
.B2(n_2275),
.Y(n_8071)
);

AOI211xp5_ASAP7_75t_L g8072 ( 
.A1(n_8071),
.A2(n_2275),
.B(n_2136),
.C(n_2901),
.Y(n_8072)
);


endmodule