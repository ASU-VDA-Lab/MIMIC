module real_jpeg_16933_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_11;
wire n_14;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_13),
.C(n_15),
.Y(n_12)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_3),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_11)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g7 ( 
.A1(n_4),
.A2(n_8),
.B1(n_20),
.B2(n_21),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_5),
.B(n_14),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_18),
.C(n_19),
.Y(n_17)
);


endmodule