module fake_jpeg_23220_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_25),
.B(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_27),
.B1(n_16),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_13),
.Y(n_46)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_4),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_4),
.B(n_6),
.C(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_50),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_22),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_27),
.B(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_20),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_17),
.C(n_32),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_62),
.C(n_12),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_65),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_21),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_51),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_66),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_20),
.B(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_74),
.B1(n_57),
.B2(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_65),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_75),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_29),
.C(n_40),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_59),
.C(n_12),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_54),
.B1(n_58),
.B2(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_63),
.B(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_70),
.B(n_77),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_89),
.B(n_91),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_73),
.B(n_71),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_59),
.B(n_32),
.C(n_34),
.D(n_29),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_82),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_29),
.C(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_6),
.B(n_8),
.Y(n_97)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_98),
.B(n_92),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_100),
.B(n_99),
.C(n_9),
.D(n_15),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_99),
.B1(n_44),
.B2(n_45),
.C(n_21),
.Y(n_103)
);


endmodule