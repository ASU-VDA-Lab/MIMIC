module fake_aes_9748_n_593 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_593);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_593;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g71 ( .A(n_23), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_38), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_54), .Y(n_73) );
INVxp33_ASAP7_75t_SL g74 ( .A(n_46), .Y(n_74) );
INVxp33_ASAP7_75t_SL g75 ( .A(n_44), .Y(n_75) );
BUFx6f_ASAP7_75t_L g76 ( .A(n_67), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_9), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_28), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_62), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_24), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_68), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_66), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_0), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_48), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_5), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_33), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_29), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_57), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_40), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_56), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_17), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_2), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_43), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_0), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_53), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_45), .B(n_34), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_60), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_69), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_11), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_84), .B(n_1), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g118 ( .A(n_79), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_84), .B(n_2), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_102), .B(n_3), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_82), .B(n_3), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_103), .B(n_4), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_73), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_89), .B(n_4), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_114), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_73), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_78), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_90), .B(n_6), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
NAND2xp33_ASAP7_75t_L g144 ( .A(n_80), .B(n_30), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_82), .B(n_6), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_107), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_107), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_86), .B(n_7), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_152), .B(n_111), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_152), .B(n_111), .Y(n_155) );
AO22x2_ASAP7_75t_L g156 ( .A1(n_116), .A2(n_110), .B1(n_97), .B2(n_86), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_132), .B(n_87), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_153), .B(n_110), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_118), .B(n_74), .Y(n_162) );
OR2x2_ASAP7_75t_SL g163 ( .A(n_116), .B(n_97), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_115), .B(n_88), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_101), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_141), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_115), .B(n_88), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_141), .B(n_104), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_141), .B(n_98), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_120), .B(n_127), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_117), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_117), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_117), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_128), .B(n_98), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_118), .B(n_75), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_128), .B(n_93), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_129), .B(n_101), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_119), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_119), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_129), .B(n_94), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_130), .B(n_78), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_127), .B(n_106), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_122), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_122), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_118), .B(n_108), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_130), .B(n_104), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_120), .B(n_100), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_121), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_122), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_124), .Y(n_200) );
AND2x6_ASAP7_75t_L g201 ( .A(n_124), .B(n_106), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_121), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_134), .B(n_105), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_137), .B(n_92), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_123), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_201), .Y(n_208) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_173), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_198), .A2(n_150), .B1(n_126), .B2(n_153), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_205), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_175), .B(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_156), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_156), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_180), .B(n_135), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_173), .Y(n_216) );
BUFx4f_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_169), .B(n_150), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_156), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_180), .B(n_139), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_158), .B(n_135), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_182), .B(n_143), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_200), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_200), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_185), .A2(n_146), .B(n_149), .C(n_143), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_171), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_169), .B(n_126), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_165), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_168), .B(n_149), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_194), .B(n_92), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_203), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_168), .B(n_139), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_191), .B(n_147), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_191), .B(n_147), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_161), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_164), .B(n_131), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_164), .B(n_134), .Y(n_246) );
OR2x2_ASAP7_75t_SL g247 ( .A(n_203), .B(n_105), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_164), .B(n_134), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
NAND3xp33_ASAP7_75t_SL g251 ( .A(n_197), .B(n_95), .C(n_109), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_170), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_197), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_170), .Y(n_255) );
OAI22xp5_ASAP7_75t_SL g256 ( .A1(n_163), .A2(n_77), .B1(n_96), .B2(n_151), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_167), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_162), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_154), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_167), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
AOI22xp33_ASAP7_75t_SL g262 ( .A1(n_238), .A2(n_171), .B1(n_183), .B2(n_155), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_208), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
BUFx2_ASAP7_75t_SL g268 ( .A(n_216), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_213), .A2(n_171), .B1(n_204), .B2(n_170), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_216), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_253), .A2(n_171), .B1(n_179), .B2(n_186), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_214), .A2(n_204), .B1(n_186), .B2(n_179), .Y(n_275) );
INVx4_ASAP7_75t_L g276 ( .A(n_208), .Y(n_276) );
AO22x2_ASAP7_75t_L g277 ( .A1(n_218), .A2(n_186), .B1(n_206), .B2(n_163), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_209), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_259), .B(n_160), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_208), .B(n_206), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_247), .B(n_212), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_258), .B(n_184), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_234), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_204), .B1(n_195), .B2(n_202), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_227), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_243), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_210), .B(n_189), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_215), .A2(n_190), .B(n_196), .Y(n_292) );
CKINVDCx8_ASAP7_75t_R g293 ( .A(n_222), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_234), .Y(n_294) );
INVx5_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_225), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_220), .A2(n_135), .B1(n_140), .B2(n_138), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_234), .B(n_140), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_215), .A2(n_144), .B(n_159), .Y(n_301) );
OR2x6_ASAP7_75t_L g302 ( .A(n_243), .B(n_151), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_239), .B(n_135), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_256), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_304), .A2(n_251), .B1(n_219), .B2(n_231), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_300), .B(n_239), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_285), .B(n_240), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_271), .Y(n_311) );
INVx6_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_300), .B(n_219), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_291), .A2(n_221), .B(n_246), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_274), .A2(n_219), .B1(n_231), .B2(n_217), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_301), .A2(n_159), .B(n_157), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_286), .B(n_241), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_304), .A2(n_231), .B1(n_211), .B2(n_237), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_284), .A2(n_237), .B1(n_222), .B2(n_245), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_267), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_275), .A2(n_217), .B1(n_230), .B2(n_248), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_265), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_262), .B(n_228), .C(n_224), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_294), .A2(n_222), .B1(n_248), .B2(n_224), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_267), .B(n_235), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_265), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_228), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_272), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_282), .A2(n_230), .B1(n_140), .B2(n_142), .C(n_138), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_310), .A2(n_277), .B1(n_293), .B2(n_283), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_316), .B(n_283), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_308), .A2(n_277), .B1(n_222), .B2(n_283), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_315), .A2(n_292), .B(n_303), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_306), .B(n_293), .Y(n_338) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_317), .A2(n_133), .B(n_148), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_313), .B(n_288), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_273), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_329), .A2(n_288), .B1(n_269), .B2(n_298), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_317), .A2(n_133), .B(n_148), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_329), .A2(n_298), .B1(n_264), .B2(n_297), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_327), .B(n_290), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_309), .B(n_280), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_133), .B(n_148), .C(n_151), .Y(n_348) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_325), .A2(n_287), .B(n_138), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_319), .A2(n_264), .B1(n_298), .B2(n_299), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_325), .B(n_174), .C(n_166), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_330), .A2(n_264), .B1(n_299), .B2(n_296), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_322), .A2(n_140), .B1(n_142), .B2(n_302), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_305), .A2(n_142), .B1(n_140), .B2(n_273), .C(n_289), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_313), .A2(n_296), .B1(n_302), .B2(n_289), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_334), .A2(n_320), .B1(n_331), .B2(n_326), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_333), .A2(n_305), .A3(n_307), .B(n_311), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_336), .A2(n_314), .B1(n_307), .B2(n_311), .C(n_323), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_343), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_343), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_339), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_351), .A2(n_328), .B(n_324), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_314), .B(n_123), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_349), .A2(n_281), .B(n_302), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_334), .A2(n_327), .B1(n_321), .B2(n_312), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_333), .A2(n_327), .B1(n_321), .B2(n_302), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_334), .A2(n_327), .B1(n_321), .B2(n_312), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_344), .A2(n_157), .B(n_172), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_337), .A2(n_279), .B(n_243), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_341), .B(n_281), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_347), .B(n_123), .C(n_125), .D(n_12), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_350), .A2(n_276), .B1(n_266), .B2(n_295), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_346), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_276), .B1(n_266), .B2(n_295), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
OAI33xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_125), .A3(n_172), .B1(n_199), .B2(n_192), .B3(n_178), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_125), .B(n_276), .C(n_174), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_352), .A2(n_290), .B1(n_295), .B2(n_249), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_345), .A2(n_229), .B1(n_232), .B2(n_260), .C(n_257), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_346), .B(n_8), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
OAI221xp5_ASAP7_75t_SL g387 ( .A1(n_357), .A2(n_349), .B1(n_342), .B2(n_355), .C(n_340), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_360), .B(n_340), .Y(n_388) );
NAND2xp33_ASAP7_75t_L g389 ( .A(n_370), .B(n_335), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_376), .A2(n_332), .B1(n_340), .B2(n_335), .C(n_354), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
OR2x2_ASAP7_75t_SL g392 ( .A(n_363), .B(n_332), .Y(n_392) );
OAI31xp33_ASAP7_75t_L g393 ( .A1(n_376), .A2(n_346), .A3(n_244), .B(n_254), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_366), .B(n_332), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_358), .A2(n_174), .B1(n_166), .B2(n_192), .C(n_199), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_385), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_357), .A2(n_166), .B(n_174), .C(n_295), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_8), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_166), .B(n_174), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_366), .B(n_61), .Y(n_405) );
AOI31xp33_ASAP7_75t_L g406 ( .A1(n_385), .A2(n_9), .A3(n_13), .B(n_14), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_368), .B(n_13), .Y(n_407) );
AOI33xp33_ASAP7_75t_L g408 ( .A1(n_356), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_18), .B3(n_178), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_378), .B(n_18), .Y(n_410) );
OAI33xp33_ASAP7_75t_L g411 ( .A1(n_386), .A2(n_207), .A3(n_232), .B1(n_250), .B2(n_257), .B3(n_260), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_380), .B(n_166), .C(n_176), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_19), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_279), .B1(n_290), .B2(n_261), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_368), .B(n_20), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_369), .A2(n_250), .B(n_207), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_365), .A2(n_279), .B1(n_261), .B2(n_233), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_371), .B(n_21), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_369), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_363), .B(n_279), .Y(n_422) );
AOI21xp5_ASAP7_75t_SL g423 ( .A1(n_364), .A2(n_254), .B(n_249), .Y(n_423) );
NAND3xp33_ASAP7_75t_SL g424 ( .A(n_382), .B(n_22), .C(n_25), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_193), .B1(n_177), .B2(n_181), .C(n_187), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_375), .B(n_26), .Y(n_426) );
OAI322xp33_ASAP7_75t_SL g427 ( .A1(n_384), .A2(n_27), .A3(n_31), .B1(n_32), .B2(n_35), .C1(n_36), .C2(n_37), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_372), .B(n_39), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_372), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_362), .B(n_41), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_389), .A2(n_381), .B1(n_377), .B2(n_379), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_421), .B(n_362), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_404), .B(n_362), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_406), .A2(n_181), .B1(n_193), .B2(n_188), .C(n_187), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_403), .B(n_373), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_415), .B(n_47), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_383), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_413), .B(n_49), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_394), .B(n_50), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_394), .B(n_55), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_395), .B(n_58), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
OAI322xp33_ASAP7_75t_L g446 ( .A1(n_407), .A2(n_188), .A3(n_193), .B1(n_187), .B2(n_176), .C1(n_177), .C2(n_181), .Y(n_446) );
AOI33xp33_ASAP7_75t_L g447 ( .A1(n_398), .A2(n_59), .A3(n_63), .B1(n_65), .B2(n_176), .B3(n_177), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_407), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_401), .B(n_176), .Y(n_450) );
AND4x1_ASAP7_75t_L g451 ( .A(n_408), .B(n_261), .C(n_244), .D(n_235), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_409), .B(n_177), .Y(n_452) );
NOR2x1p5_ASAP7_75t_SL g453 ( .A(n_431), .B(n_429), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_429), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_430), .B(n_177), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_410), .B(n_181), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_405), .B(n_261), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_388), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_417), .B(n_181), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_417), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_400), .B(n_187), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
NAND3x1_ASAP7_75t_L g464 ( .A(n_408), .B(n_233), .C(n_236), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_426), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_431), .Y(n_468) );
NAND2xp33_ASAP7_75t_R g469 ( .A(n_396), .B(n_233), .Y(n_469) );
INVx6_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_389), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_428), .B(n_188), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_390), .B(n_188), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_422), .B(n_188), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_393), .A2(n_193), .B1(n_236), .B2(n_411), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_416), .B(n_193), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_392), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_387), .B(n_236), .C(n_420), .D(n_399), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_418), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_466), .B(n_422), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_459), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_459), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_471), .B(n_392), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_437), .B(n_402), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_458), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_467), .B(n_423), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_461), .B(n_397), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_443), .B(n_412), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_443), .B(n_423), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_475), .B(n_419), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_463), .B(n_427), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_435), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_435), .B(n_424), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_435), .B(n_425), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_465), .B(n_482), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_439), .B(n_434), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_473), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_470), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_480), .B(n_433), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_433), .B(n_453), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_474), .B(n_468), .Y(n_507) );
AOI32xp33_ASAP7_75t_L g508 ( .A1(n_436), .A2(n_473), .A3(n_440), .B1(n_438), .B2(n_432), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_433), .B(n_454), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_451), .B(n_481), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_455), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_470), .B(n_472), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_472), .B(n_440), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_452), .B(n_478), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_478), .B(n_441), .Y(n_517) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_457), .B(n_440), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_441), .B(n_442), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_446), .A2(n_457), .B(n_479), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_442), .B(n_444), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_444), .B(n_438), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_506), .B(n_447), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_503), .B(n_487), .Y(n_524) );
AOI21xp33_ASAP7_75t_SL g525 ( .A1(n_518), .A2(n_469), .B(n_438), .Y(n_525) );
XOR2x2_ASAP7_75t_L g526 ( .A(n_518), .B(n_464), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_484), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_510), .A2(n_464), .B1(n_479), .B2(n_456), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_501), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_506), .B(n_508), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_502), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_498), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_485), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_497), .B(n_462), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_494), .Y(n_536) );
OAI211xp5_ASAP7_75t_L g537 ( .A1(n_510), .A2(n_477), .B(n_469), .C(n_460), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_520), .A2(n_447), .B(n_476), .Y(n_538) );
AND2x2_ASAP7_75t_SL g539 ( .A(n_506), .B(n_511), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_499), .B(n_493), .C(n_489), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_504), .B(n_500), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_486), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_507), .B(n_511), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_505), .B(n_509), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_505), .B(n_489), .Y(n_546) );
OAI21xp33_ASAP7_75t_SL g547 ( .A1(n_492), .A2(n_495), .B(n_483), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g548 ( .A(n_504), .B(n_505), .Y(n_548) );
BUFx12f_ASAP7_75t_L g549 ( .A(n_516), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_492), .A2(n_522), .B(n_515), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_496), .B(n_490), .Y(n_552) );
AOI211x1_ASAP7_75t_SL g553 ( .A1(n_512), .A2(n_513), .B(n_514), .C(n_519), .Y(n_553) );
XNOR2x1_ASAP7_75t_L g554 ( .A(n_517), .B(n_521), .Y(n_554) );
XNOR2xp5_ASAP7_75t_L g555 ( .A(n_490), .B(n_514), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_510), .A2(n_406), .B(n_497), .C(n_503), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_501), .B(n_487), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_510), .A2(n_464), .B(n_406), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_505), .A2(n_508), .B(n_489), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_501), .B(n_487), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_484), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g563 ( .A1(n_556), .A2(n_530), .B(n_558), .C(n_559), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_541), .B(n_540), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_540), .A2(n_526), .B1(n_535), .B2(n_549), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_543), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_532), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_553), .B(n_552), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_548), .B(n_554), .Y(n_569) );
AOI21xp33_ASAP7_75t_SL g570 ( .A1(n_539), .A2(n_523), .B(n_548), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_535), .B(n_529), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_547), .A2(n_539), .B1(n_528), .B2(n_546), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_524), .A2(n_562), .B1(n_551), .B2(n_546), .C(n_560), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g575 ( .A1(n_565), .A2(n_538), .B(n_537), .C(n_544), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_563), .A2(n_549), .B1(n_536), .B2(n_555), .Y(n_576) );
OAI211xp5_ASAP7_75t_SL g577 ( .A1(n_572), .A2(n_537), .B(n_544), .C(n_557), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_564), .B(n_536), .Y(n_578) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_570), .A2(n_525), .B(n_536), .C(n_555), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_569), .A2(n_554), .B1(n_545), .B2(n_533), .Y(n_580) );
OR3x1_ASAP7_75t_L g581 ( .A(n_566), .B(n_531), .C(n_561), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_576), .B(n_564), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_581), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_575), .B(n_568), .Y(n_584) );
OR4x1_ASAP7_75t_L g585 ( .A(n_579), .B(n_567), .C(n_527), .D(n_550), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g586 ( .A1(n_584), .A2(n_580), .B1(n_578), .B2(n_573), .C1(n_571), .C2(n_577), .Y(n_586) );
OR4x1_ASAP7_75t_L g587 ( .A(n_583), .B(n_542), .C(n_534), .D(n_574), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_587), .Y(n_588) );
AND2x2_ASAP7_75t_SL g589 ( .A(n_587), .B(n_585), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_589), .B(n_582), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_590), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_591), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_592), .A2(n_588), .B(n_586), .Y(n_593) );
endmodule