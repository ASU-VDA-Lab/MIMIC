module real_jpeg_18033_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_27),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_2),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_2),
.B(n_51),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_4),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_25),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_149),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_8),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_8),
.B(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_8),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_8),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_9),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_9),
.B(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22x1_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_12),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_10),
.B(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

AOI31xp33_ASAP7_75t_L g39 ( 
.A1(n_12),
.A2(n_40),
.A3(n_43),
.B(n_49),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_12),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_12),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_12),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_12),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_12),
.B(n_202),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_13),
.B(n_136),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_14),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_170),
.B1(n_282),
.B2(n_283),
.Y(n_17)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_18),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_168),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_128),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g169 ( 
.A(n_20),
.B(n_128),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_66),
.C(n_111),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_21),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_22),
.B(n_39),
.C(n_54),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_29),
.C(n_34),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_23),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_SL g214 ( 
.A(n_24),
.B(n_26),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_24),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_24),
.A2(n_235),
.B1(n_236),
.B2(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_25),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_29),
.Y(n_268)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_54),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_49),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_49),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_59),
.C(n_62),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_61),
.B(n_178),
.C(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2x2_ASAP7_75t_SL g176 ( 
.A(n_62),
.B(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_67),
.B(n_111),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_85),
.C(n_100),
.Y(n_67)
);

XOR2x1_ASAP7_75t_L g272 ( 
.A(n_68),
.B(n_273),
.Y(n_272)
);

XOR2x2_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_76),
.C(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_76),
.A2(n_84),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_76),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_86),
.B(n_101),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_95),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_87),
.A2(n_95),
.B1(n_96),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2x2_ASAP7_75t_L g208 ( 
.A(n_91),
.B(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_96),
.B1(n_139),
.B2(n_143),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_105),
.Y(n_126)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_125),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_122),
.C(n_124),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_118),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_131),
.C(n_132),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_151),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_150),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_170),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_276),
.B(n_281),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_261),
.B(n_275),
.Y(n_172)
);

OAI21x1_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_220),
.B(n_260),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_205),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_205),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.C(n_196),
.Y(n_175)
);

XOR2x1_ASAP7_75t_L g254 ( 
.A(n_176),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_187),
.A2(n_188),
.B1(n_196),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_192),
.Y(n_225)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_214),
.C(n_215),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21x1_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_253),
.B(n_259),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_237),
.B(n_252),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_228),
.C(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_244),
.B(n_251),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_274),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_272),
.Y(n_262)
);

INVxp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.C(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_279),
.Y(n_281)
);


endmodule