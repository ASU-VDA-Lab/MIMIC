module real_jpeg_19011_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_322, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_322;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_0),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_160),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_160),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_26),
.B1(n_35),
.B2(n_160),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_50),
.B(n_60),
.C(n_146),
.D(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_3),
.B(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_48),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_3),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_83),
.B(n_165),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_32),
.B(n_43),
.C(n_197),
.D(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_133),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_3),
.A2(n_31),
.B(n_33),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_26),
.B1(n_35),
.B2(n_179),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_26),
.B1(n_35),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_131),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_131),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_131),
.Y(n_253)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_26),
.B1(n_35),
.B2(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_6),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_7),
.B(n_65),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_7),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_84),
.B1(n_208),
.B2(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_8),
.A2(n_38),
.B1(n_64),
.B2(n_65),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_10),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_10),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_26),
.B1(n_35),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_11),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_93),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_93),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_93),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_109),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_95),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_21),
.B(n_95),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_79),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_22),
.A2(n_71),
.B1(n_72),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_22),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_23),
.A2(n_24),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_57),
.C(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_25),
.A2(n_30),
.B1(n_37),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_25),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_25),
.A2(n_30),
.B1(n_130),
.B2(n_265),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_26),
.A2(n_28),
.B(n_179),
.C(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_30),
.A2(n_34),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_30),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_30),
.A2(n_91),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_44),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_42),
.A2(n_54),
.B1(n_217),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_42),
.A2(n_253),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_48),
.B1(n_52),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_43),
.A2(n_48),
.B1(n_74),
.B2(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_43),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_44),
.B(n_50),
.Y(n_205)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_49),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_54),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_54),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_54),
.A2(n_218),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_58),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_67),
.B1(n_77),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_59),
.A2(n_67),
.B1(n_88),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_59),
.A2(n_67),
.B1(n_159),
.B2(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_59),
.A2(n_195),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_59),
.A2(n_67),
.B1(n_125),
.B2(n_250),
.Y(n_275)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_63),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_60),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_61),
.B(n_65),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_62),
.A2(n_64),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_65),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_67),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_67),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_67),
.B(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_67),
.A2(n_161),
.B(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_90),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_81),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_82),
.A2(n_87),
.B1(n_89),
.B2(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_86),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_83),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_83),
.A2(n_123),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_83),
.A2(n_122),
.B1(n_243),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_84),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_84),
.B(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_85),
.A2(n_171),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_181),
.B(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_85),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_87),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_94),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_137),
.B(n_320),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_134),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_111),
.B(n_134),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_112),
.A2(n_116),
.B1(n_117),
.B2(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_112),
.Y(n_307)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_118),
.A2(n_119),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_128),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_120),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_121),
.B(n_124),
.Y(n_280)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_123),
.B(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_126),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_127),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_132),
.Y(n_257)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_295),
.A3(n_308),
.B1(n_314),
.B2(n_319),
.C(n_322),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_259),
.C(n_291),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_232),
.B(n_258),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_211),
.B(n_231),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_189),
.B(n_210),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_167),
.B(n_188),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_158),
.C(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_176),
.B(n_187),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_174),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_182),
.B(n_186),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_202),
.B2(n_209),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_200),
.B2(n_201),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_201),
.C(n_209),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_198),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_227),
.C(n_229),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_224),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_221),
.C(n_222),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_234),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_247),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_246),
.C(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_241),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_260),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_277),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_277),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.C(n_276),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_276),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_275),
.Y(n_282)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_289),
.B2(n_290),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_281),
.C(n_290),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_286),
.C(n_288),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_284),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_293),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_304),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_296),
.B(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_301),
.C(n_303),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);


endmodule