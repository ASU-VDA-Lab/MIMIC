module fake_jpeg_21115_n_75 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_12),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_1),
.B1(n_8),
.B2(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_8),
.B(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_41),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_42),
.B(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_14),
.B(n_15),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_32),
.B(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_28),
.B(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_24),
.B1(n_34),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_33),
.B1(n_30),
.B2(n_24),
.Y(n_49)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_55),
.B1(n_51),
.B2(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_52),
.B(n_54),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_39),
.C(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_48),
.B1(n_40),
.B2(n_38),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_62),
.B(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_58),
.B1(n_60),
.B2(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_52),
.C(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_46),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_69),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_73),
.Y(n_75)
);


endmodule