module fake_netlist_6_3694_n_96 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_96);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_96;

wire n_52;
wire n_91;
wire n_46;
wire n_88;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_92;
wire n_42;
wire n_90;
wire n_24;
wire n_54;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_25;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AND2x4_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_21),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_18),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_4),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_2),
.B1(n_6),
.B2(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_26),
.B2(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_24),
.B(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_36),
.B1(n_38),
.B2(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_23),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_38),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_R g56 ( 
.A(n_55),
.B(n_26),
.Y(n_56)
);

AO21x2_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_47),
.B(n_32),
.Y(n_57)
);

OAI21x1_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_42),
.B(n_40),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_32),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_40),
.B(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_23),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AND2x4_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_58),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_61),
.B1(n_56),
.B2(n_64),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_54),
.C(n_49),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_61),
.A3(n_67),
.B1(n_68),
.B2(n_27),
.C(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

OAI221xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_61),
.B1(n_66),
.B2(n_53),
.C(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_61),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_70),
.C(n_27),
.Y(n_83)
);

NAND5xp2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_28),
.C(n_72),
.D(n_25),
.E(n_53),
.Y(n_84)
);

NOR3x2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_76),
.C(n_57),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_74),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_82),
.B(n_57),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_57),
.B(n_25),
.Y(n_92)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_25),
.B1(n_74),
.B2(n_66),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_89),
.B(n_88),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_90),
.B(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);


endmodule