module fake_jpeg_15607_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_0),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_33),
.B(n_18),
.Y(n_80)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_2),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_61),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_16),
.A2(n_31),
.B1(n_18),
.B2(n_37),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_17),
.B1(n_31),
.B2(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_17),
.B(n_2),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_66),
.B(n_71),
.Y(n_117)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_20),
.B(n_24),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_78),
.B(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_74),
.B(n_83),
.Y(n_132)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_61),
.C(n_28),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_5),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_98),
.Y(n_131)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_26),
.B1(n_29),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_91),
.Y(n_124)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_26),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_40),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_107)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_35),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_28),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_39),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_133),
.Y(n_142)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_110),
.Y(n_147)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_119),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_99),
.B(n_13),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_38),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_38),
.B1(n_30),
.B2(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_121),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_38),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_134),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_73),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_30),
.B1(n_6),
.B2(n_9),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_30),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_9),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_93),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_68),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_146),
.B(n_148),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_11),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_13),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_70),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_67),
.C(n_97),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_133),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_112),
.B1(n_128),
.B2(n_118),
.Y(n_174)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_65),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_163),
.B(n_166),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_67),
.B(n_90),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_112),
.B(n_107),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_90),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_170),
.C(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_167),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_82),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_88),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_88),
.B(n_95),
.C(n_76),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_140),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g169 ( 
.A(n_117),
.B(n_97),
.C(n_72),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_171),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_72),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_141),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_194),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_165),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_132),
.C(n_137),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_189),
.C(n_191),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_158),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_158),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_117),
.C(n_123),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_108),
.C(n_129),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_110),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_111),
.B(n_115),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_204),
.C(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_165),
.C(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_143),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_207),
.Y(n_220)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_169),
.A3(n_150),
.B1(n_143),
.B2(n_142),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_143),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_162),
.C(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_199),
.B1(n_205),
.B2(n_201),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_199),
.B1(n_202),
.B2(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_189),
.C(n_191),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_193),
.C(n_190),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_187),
.B1(n_174),
.B2(n_195),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_163),
.B1(n_183),
.B2(n_204),
.Y(n_232)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_193),
.B(n_190),
.C(n_148),
.D(n_146),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_223),
.B(n_148),
.C(n_146),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_194),
.B(n_163),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_176),
.B(n_212),
.C(n_200),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_223),
.B1(n_179),
.B2(n_113),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_227),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_203),
.B(n_209),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_232),
.B(n_224),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_216),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_217),
.B(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_151),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_243),
.C(n_233),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_225),
.B(n_216),
.C(n_176),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_242),
.A2(n_236),
.B1(n_228),
.B2(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_242),
.C(n_185),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_249),
.C(n_130),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_181),
.Y(n_252)
);


endmodule