module fake_jpeg_8541_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_68),
.B1(n_27),
.B2(n_33),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_26),
.B1(n_29),
.B2(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_24),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_80),
.Y(n_113)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_29),
.B1(n_27),
.B2(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_77),
.B1(n_83),
.B2(n_18),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_26),
.B1(n_39),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_55),
.B1(n_54),
.B2(n_47),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_25),
.Y(n_105)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_17),
.B1(n_23),
.B2(n_30),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_32),
.B(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_64),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_33),
.B1(n_18),
.B2(n_32),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AND2x4_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_42),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_98),
.B(n_101),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_56),
.C(n_47),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_71),
.B1(n_80),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_20),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_20),
.B(n_42),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_108),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_40),
.C(n_36),
.Y(n_106)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_49),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_43),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_53),
.C(n_91),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_116),
.B1(n_120),
.B2(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_89),
.C(n_34),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_137),
.C(n_138),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_123),
.A2(n_60),
.B(n_28),
.Y(n_173)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_92),
.B1(n_85),
.B2(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_131),
.B1(n_143),
.B2(n_76),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_92),
.B1(n_78),
.B2(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_111),
.B1(n_114),
.B2(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_136),
.B1(n_146),
.B2(n_94),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_141),
.B(n_42),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_65),
.B1(n_67),
.B2(n_84),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_91),
.C(n_43),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_84),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_42),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_34),
.B1(n_36),
.B2(n_46),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_36),
.B1(n_60),
.B2(n_51),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_120),
.B1(n_115),
.B2(n_119),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_161),
.B(n_170),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_154),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_110),
.B1(n_94),
.B2(n_76),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_169),
.B1(n_125),
.B2(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_0),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_157),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_20),
.B(n_30),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_165),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_132),
.B1(n_121),
.B2(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_173),
.B1(n_126),
.B2(n_124),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_166),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_15),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_115),
.C(n_42),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_137),
.C(n_141),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_24),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_181),
.B1(n_150),
.B2(n_30),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_188),
.C(n_190),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_164),
.B(n_155),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_187),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_154),
.C(n_163),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_161),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_142),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_195),
.C(n_42),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_203),
.B(n_208),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_158),
.B(n_156),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_204),
.A2(n_206),
.B(n_209),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_162),
.B1(n_168),
.B2(n_158),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_205),
.A2(n_217),
.B1(n_186),
.B2(n_179),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_200),
.B(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_159),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_24),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_150),
.B1(n_118),
.B2(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_225),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_103),
.B1(n_23),
.B2(n_28),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_224),
.C(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_103),
.B1(n_28),
.B2(n_3),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_103),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_229),
.C(n_216),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_188),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_208),
.C(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_195),
.C(n_180),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_182),
.C(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_237),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_180),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_246),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_179),
.B1(n_183),
.B2(n_64),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_238),
.B1(n_217),
.B2(n_209),
.Y(n_248)
);

XOR2x1_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_24),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_14),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_24),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_15),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_258),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_228),
.C(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_218),
.C(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_256),
.C(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_214),
.C(n_203),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_202),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_201),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_13),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_271),
.C(n_1),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_231),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_270),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_236),
.B(n_244),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_272),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_230),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_2),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_236),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_2),
.C(n_3),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_13),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_263),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_280),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

OAI21x1_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_11),
.B(n_9),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_1),
.B(n_2),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_288),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_291),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_290),
.A2(n_269),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_4),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_264),
.Y(n_294)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_289),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_306),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_271),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_264),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_265),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_300),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_305),
.B(n_302),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_310),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_299),
.B(n_286),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_311),
.C(n_297),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_297),
.B(n_281),
.C(n_279),
.D(n_7),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.C(n_5),
.Y(n_319)
);

OAI221xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_4),
.B1(n_7),
.B2(n_315),
.C(n_305),
.Y(n_320)
);


endmodule