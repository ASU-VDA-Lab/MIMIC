module fake_aes_9430_n_658 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_658);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g89 ( .A(n_19), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_3), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_47), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_55), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_51), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_4), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_11), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_50), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_69), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_79), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_38), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_31), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_83), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_4), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_17), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_73), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_84), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_21), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_25), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_81), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_34), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_62), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_20), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_49), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_0), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_28), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_46), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_14), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_40), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_68), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_59), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_65), .Y(n_132) );
INVxp33_ASAP7_75t_L g133 ( .A(n_72), .Y(n_133) );
NOR2x1_ASAP7_75t_L g134 ( .A(n_90), .B(n_1), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_100), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_97), .B(n_114), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_124), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_107), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_92), .B(n_1), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_133), .B(n_2), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_132), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_96), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_125), .B(n_2), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_101), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_93), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_97), .B(n_5), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_151), .A2(n_111), .B1(n_109), .B2(n_128), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_157), .B(n_158), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_159), .B(n_127), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_159), .B(n_103), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g172 ( .A(n_146), .B(n_111), .C(n_128), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_135), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_157), .B(n_158), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
AND2x6_ASAP7_75t_L g176 ( .A(n_159), .B(n_104), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_160), .B(n_105), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_152), .A2(n_126), .B1(n_108), .B2(n_110), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_142), .A2(n_109), .B1(n_91), .B2(n_123), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_146), .B(n_115), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_157), .B(n_95), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_160), .B(n_106), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_144), .B(n_119), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_149), .B(n_130), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_149), .B(n_130), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_166), .B(n_152), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_169), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_179), .A2(n_139), .B1(n_156), .B2(n_154), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_179), .B(n_154), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_162), .A2(n_156), .B(n_136), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_162), .B(n_95), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_171), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_180), .A2(n_136), .B(n_120), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_161), .Y(n_205) );
NAND3xp33_ASAP7_75t_SL g206 ( .A(n_172), .B(n_138), .C(n_137), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_178), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_185), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_190), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_191), .B(n_98), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_193), .B(n_98), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_169), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_185), .A2(n_134), .B1(n_155), .B2(n_150), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_168), .B(n_129), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_187), .B(n_112), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
OAI21xp33_ASAP7_75t_L g218 ( .A1(n_167), .A2(n_134), .B(n_150), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_190), .B(n_112), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_163), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_169), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_168), .B(n_147), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_183), .Y(n_226) );
AND3x1_ASAP7_75t_L g227 ( .A(n_189), .B(n_121), .C(n_122), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_164), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_190), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_165), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_174), .B(n_116), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_168), .B(n_155), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_176), .B(n_155), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_183), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
INVxp67_ASAP7_75t_L g238 ( .A(n_194), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_194), .B(n_179), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_221), .B(n_185), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_229), .B(n_182), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_195), .Y(n_242) );
INVxp67_ASAP7_75t_SL g243 ( .A(n_209), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_196), .B(n_185), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_199), .B(n_185), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_205), .B(n_185), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_203), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_205), .B(n_176), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_232), .B(n_184), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_201), .A2(n_150), .B(n_117), .C(n_192), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_208), .A2(n_179), .B1(n_176), .B2(n_113), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_199), .A2(n_89), .B(n_118), .C(n_145), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_208), .Y(n_257) );
CKINVDCx11_ASAP7_75t_R g258 ( .A(n_234), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_224), .B(n_176), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_212), .Y(n_261) );
AO22x1_ASAP7_75t_L g262 ( .A1(n_212), .A2(n_176), .B1(n_123), .B2(n_116), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_210), .A2(n_165), .B(n_186), .Y(n_266) );
AO21x1_ASAP7_75t_L g267 ( .A1(n_204), .A2(n_188), .B(n_170), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_234), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_224), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_216), .A2(n_148), .B(n_145), .C(n_175), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_216), .B(n_188), .Y(n_271) );
CKINVDCx8_ASAP7_75t_R g272 ( .A(n_198), .Y(n_272) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_226), .A2(n_188), .B(n_170), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_211), .A2(n_186), .B(n_175), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_234), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_235), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_224), .B(n_140), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g279 ( .A(n_206), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_267), .A2(n_213), .B(n_227), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_242), .B(n_198), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_267), .A2(n_218), .B(n_173), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_273), .A2(n_173), .B(n_236), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_237), .B(n_245), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_237), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_273), .A2(n_236), .B(n_235), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_231), .B(n_230), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_250), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_222), .B(n_225), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_258), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_250), .B(n_198), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_233), .B(n_214), .Y(n_293) );
O2A1O1Ixp5_ASAP7_75t_L g294 ( .A1(n_244), .A2(n_219), .B(n_202), .C(n_233), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_263), .B(n_233), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_238), .B(n_215), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_263), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_275), .A2(n_231), .B(n_230), .Y(n_298) );
AO21x1_ASAP7_75t_L g299 ( .A1(n_274), .A2(n_220), .B(n_143), .Y(n_299) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_261), .Y(n_300) );
INVx4_ASAP7_75t_SL g301 ( .A(n_261), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_245), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_254), .B(n_140), .C(n_143), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_243), .B(n_200), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_252), .A2(n_220), .B(n_140), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_274), .A2(n_192), .B(n_143), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_239), .B(n_200), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_248), .A2(n_200), .B(n_198), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_239), .B(n_228), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_261), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_SL g313 ( .A1(n_259), .A2(n_145), .B(n_148), .C(n_45), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_289), .A2(n_247), .B1(n_240), .B2(n_251), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_285), .B(n_277), .Y(n_317) );
AO31x2_ASAP7_75t_L g318 ( .A1(n_299), .A2(n_277), .A3(n_278), .B(n_246), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_286), .B(n_251), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_293), .A2(n_249), .B1(n_253), .B2(n_279), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_291), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_293), .A2(n_276), .B1(n_268), .B2(n_241), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_302), .A2(n_265), .B1(n_242), .B2(n_276), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_296), .A2(n_268), .B1(n_269), .B2(n_265), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_296), .A2(n_260), .B1(n_264), .B2(n_270), .C(n_257), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_271), .B(n_145), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_289), .A2(n_257), .B1(n_271), .B2(n_255), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_285), .B(n_262), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_295), .A2(n_272), .B1(n_262), .B2(n_255), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g332 ( .A(n_302), .B(n_255), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_302), .B(n_228), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_308), .A2(n_228), .B(n_217), .Y(n_335) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_294), .A2(n_217), .B(n_228), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_272), .B1(n_228), .B2(n_217), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_297), .B(n_217), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_310), .B(n_217), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_297), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_304), .B1(n_307), .B2(n_311), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_319), .B(n_290), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_317), .B(n_280), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_317), .B(n_280), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_343), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_343), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_319), .B(n_280), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_338), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_284), .B(n_299), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_324), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_338), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_340), .B(n_287), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_340), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_320), .B(n_290), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_334), .B(n_311), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_339), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_332), .B(n_301), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_330), .B(n_287), .Y(n_371) );
OR2x2_ASAP7_75t_SL g372 ( .A(n_341), .B(n_287), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_352), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
O2A1O1Ixp5_ASAP7_75t_L g375 ( .A1(n_370), .A2(n_325), .B(n_331), .C(n_294), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_347), .B(n_330), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_347), .B(n_287), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_348), .B(n_287), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_348), .B(n_318), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_349), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_371), .B(n_318), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_371), .B(n_318), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_350), .A2(n_321), .B(n_326), .C(n_329), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_352), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_351), .B(n_355), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_318), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_370), .B(n_332), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_357), .B(n_318), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_353), .B(n_318), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_358), .B(n_325), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_358), .B(n_344), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_345), .A2(n_316), .B1(n_323), .B2(n_327), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_361), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_367), .B(n_344), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_362), .B(n_307), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_362), .A2(n_304), .B1(n_303), .B2(n_322), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_353), .B(n_333), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_349), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_345), .A2(n_328), .A3(n_337), .B(n_292), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_367), .B(n_333), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_385), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_383), .B(n_5), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_404), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_402), .B(n_359), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_404), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_388), .Y(n_413) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_397), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_376), .B(n_359), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_402), .B(n_372), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_376), .B(n_363), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_403), .B(n_379), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_374), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_379), .B(n_372), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_390), .B(n_364), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_388), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_399), .Y(n_429) );
AND2x4_ASAP7_75t_SL g430 ( .A(n_399), .B(n_370), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_368), .B(n_354), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_346), .B1(n_366), .B2(n_305), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_392), .B(n_364), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_381), .B(n_363), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_395), .A2(n_346), .B1(n_366), .B2(n_305), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_397), .B(n_6), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_396), .B(n_354), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_392), .B(n_354), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_381), .B(n_363), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_382), .B(n_363), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_397), .B(n_6), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_374), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_397), .B(n_360), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_382), .B(n_360), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_398), .B(n_386), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_389), .B(n_360), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_398), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_389), .B(n_365), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_377), .B(n_365), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_400), .B(n_7), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_408), .B(n_377), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_434), .B(n_394), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_434), .B(n_394), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
AND3x2_ASAP7_75t_L g461 ( .A(n_437), .B(n_406), .C(n_387), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_416), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_421), .B(n_393), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_421), .B(n_393), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_415), .B(n_378), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_415), .B(n_378), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_448), .B(n_387), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_448), .B(n_407), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_427), .B(n_406), .Y(n_474) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_445), .B(n_414), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_409), .A2(n_407), .B1(n_305), .B2(n_380), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_417), .B(n_380), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_417), .B(n_405), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_428), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_430), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_425), .B(n_405), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_419), .B(n_405), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_412), .Y(n_485) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_414), .B(n_365), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_430), .B(n_368), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_428), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_419), .B(n_368), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_425), .B(n_369), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_422), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_430), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_456), .B(n_7), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_444), .B(n_435), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_427), .B(n_375), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_435), .B(n_356), .Y(n_498) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_444), .B(n_369), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_442), .B(n_369), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_356), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_440), .B(n_356), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_411), .B(n_356), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_438), .B(n_356), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_442), .B(n_305), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_443), .B(n_284), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_413), .B(n_148), .C(n_284), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_443), .B(n_8), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_455), .B(n_8), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_9), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_441), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_438), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_455), .B(n_282), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_441), .Y(n_515) );
NAND3xp33_ASAP7_75t_SL g516 ( .A(n_495), .B(n_433), .C(n_436), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_463), .B(n_452), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_495), .B(n_449), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_463), .B(n_452), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_482), .A2(n_413), .B(n_454), .C(n_423), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_494), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_482), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_464), .B(n_429), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g524 ( .A1(n_511), .A2(n_410), .B(n_447), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_471), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_467), .B(n_451), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_461), .A2(n_412), .B1(n_426), .B2(n_431), .Y(n_528) );
OAI32xp33_ASAP7_75t_L g529 ( .A1(n_509), .A2(n_453), .A3(n_439), .B1(n_446), .B2(n_450), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_461), .A2(n_453), .B1(n_450), .B2(n_446), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_457), .B(n_143), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_486), .A2(n_300), .B(n_313), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_470), .B(n_282), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_475), .B(n_301), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_470), .B(n_282), .Y(n_535) );
OAI322xp33_ASAP7_75t_L g536 ( .A1(n_474), .A2(n_143), .A3(n_153), .B1(n_148), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_462), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_496), .B(n_487), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_468), .B(n_9), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_496), .B(n_143), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_496), .B(n_153), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_474), .A2(n_300), .B(n_336), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_469), .B(n_10), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g547 ( .A1(n_497), .A2(n_10), .B(n_11), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_458), .B(n_153), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_472), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_510), .A2(n_306), .B1(n_342), .B2(n_153), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g552 ( .A1(n_497), .A2(n_12), .B(n_13), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_480), .Y(n_553) );
OAI32xp33_ASAP7_75t_L g554 ( .A1(n_459), .A2(n_314), .A3(n_312), .B1(n_283), .B2(n_342), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_506), .A2(n_153), .B1(n_314), .B2(n_312), .Y(n_555) );
AOI21xp5_ASAP7_75t_SL g556 ( .A1(n_487), .A2(n_283), .B(n_314), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_484), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_481), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_487), .B(n_15), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_492), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_508), .A2(n_335), .B(n_298), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_473), .B(n_15), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_499), .A2(n_312), .B1(n_281), .B2(n_292), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_504), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_483), .B(n_16), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_476), .A2(n_153), .B1(n_17), .B2(n_18), .C(n_16), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_476), .B(n_309), .C(n_281), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_527), .B(n_479), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_523), .B(n_478), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_516), .B(n_508), .C(n_491), .D(n_506), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_548), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_538), .B(n_515), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_530), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
XNOR2x2_ASAP7_75t_SL g576 ( .A(n_528), .B(n_499), .Y(n_576) );
AOI31xp33_ASAP7_75t_L g577 ( .A1(n_520), .A2(n_513), .A3(n_507), .B(n_498), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_549), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_560), .B(n_515), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_541), .B(n_507), .C(n_514), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_522), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_557), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_517), .Y(n_583) );
XOR2xp5_ASAP7_75t_L g584 ( .A(n_540), .B(n_489), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_518), .B(n_514), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_519), .B(n_498), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_538), .A2(n_500), .B(n_512), .C(n_472), .Y(n_587) );
NOR2xp67_ASAP7_75t_L g588 ( .A(n_525), .B(n_512), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_526), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_542), .B(n_493), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_550), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
AO22x2_ASAP7_75t_L g594 ( .A1(n_539), .A2(n_493), .B1(n_490), .B2(n_505), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_543), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_546), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_564), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_545), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_534), .A2(n_490), .B(n_306), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_567), .B(n_309), .C(n_292), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_566), .A2(n_18), .B(n_306), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_552), .A2(n_23), .B(n_24), .Y(n_603) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_563), .B(n_292), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_597), .A2(n_533), .B1(n_535), .B2(n_559), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_582), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_571), .A2(n_524), .B1(n_552), .B2(n_547), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_572), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_578), .B(n_565), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_575), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_571), .A2(n_529), .B1(n_524), .B2(n_536), .C(n_561), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_577), .A2(n_564), .B(n_568), .C(n_554), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_551), .B1(n_562), .B2(n_558), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_598), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_578), .B(n_583), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_586), .B(n_562), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_585), .A2(n_555), .B1(n_544), .B2(n_532), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_589), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_573), .A2(n_556), .B1(n_292), .B2(n_301), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_593), .Y(n_620) );
OAI311xp33_ASAP7_75t_L g621 ( .A1(n_576), .A2(n_26), .A3(n_27), .B1(n_29), .C1(n_30), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_603), .B(n_298), .C(n_288), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_590), .B(n_574), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_587), .A2(n_306), .B(n_298), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_581), .A2(n_32), .B(n_33), .C(n_35), .Y(n_625) );
NOR2x1_ASAP7_75t_SL g626 ( .A(n_579), .B(n_301), .Y(n_626) );
AOI311xp33_ASAP7_75t_L g627 ( .A1(n_613), .A2(n_601), .A3(n_595), .B(n_596), .C(n_602), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_611), .B(n_580), .C(n_602), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_615), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_SL g630 ( .A1(n_612), .A2(n_570), .B(n_569), .C(n_588), .Y(n_630) );
AOI211xp5_ASAP7_75t_SL g631 ( .A1(n_621), .A2(n_599), .B(n_591), .C(n_604), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_623), .A2(n_594), .B1(n_584), .B2(n_592), .C(n_600), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_625), .B(n_594), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_608), .A2(n_288), .B(n_301), .Y(n_634) );
OAI211xp5_ASAP7_75t_SL g635 ( .A1(n_608), .A2(n_36), .B(n_37), .C(n_43), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g636 ( .A1(n_607), .A2(n_288), .A3(n_301), .B1(n_52), .B2(n_56), .Y(n_636) );
OA22x2_ASAP7_75t_L g637 ( .A1(n_605), .A2(n_44), .B1(n_48), .B2(n_61), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_606), .A2(n_616), .B1(n_620), .B2(n_618), .C(n_614), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_609), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_627), .A2(n_617), .B1(n_610), .B2(n_619), .C(n_622), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_629), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_639), .B(n_624), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_633), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_630), .A2(n_626), .B(n_64), .C(n_67), .Y(n_644) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_628), .B(n_63), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_638), .B(n_70), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_641), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_643), .B(n_632), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_640), .B(n_644), .C(n_646), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_642), .B(n_631), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_649), .A2(n_644), .B1(n_645), .B2(n_636), .C(n_637), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_650), .A2(n_635), .B(n_634), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_651), .A2(n_648), .B1(n_647), .B2(n_75), .Y(n_653) );
OAI22xp5_ASAP7_75t_SL g654 ( .A1(n_652), .A2(n_88), .B1(n_74), .B2(n_76), .Y(n_654) );
AND3x4_ASAP7_75t_L g655 ( .A(n_653), .B(n_71), .C(n_77), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_655), .A2(n_654), .B1(n_80), .B2(n_82), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_656), .B(n_78), .C(n_85), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_86), .B(n_87), .Y(n_658) );
endmodule