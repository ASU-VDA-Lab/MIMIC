module fake_jpeg_30620_n_359 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_8),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_53),
.Y(n_118)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_57),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_8),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_19),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_30),
.Y(n_97)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_21),
.Y(n_78)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_31),
.B1(n_18),
.B2(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_87),
.B1(n_90),
.B2(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_43),
.B1(n_37),
.B2(n_31),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_105),
.B1(n_63),
.B2(n_62),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_28),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_18),
.B1(n_29),
.B2(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_18),
.B1(n_29),
.B2(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_37),
.B1(n_30),
.B2(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_4),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_41),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_41),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_118),
.C(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_41),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_41),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_102),
.Y(n_146)
);

NAND2x1p5_ASAP7_75t_L g124 ( 
.A(n_60),
.B(n_34),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_59),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_136),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_0),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_80),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_34),
.B1(n_54),
.B2(n_51),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_134),
.A2(n_143),
.B1(n_144),
.B2(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_140),
.C(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_34),
.A3(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_96),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_34),
.C(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_156),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_34),
.B1(n_7),
.B2(n_10),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_79),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_77),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_94),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_4),
.B(n_5),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_153),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_7),
.C(n_11),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_166),
.C(n_86),
.Y(n_190)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_82),
.B(n_14),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_7),
.B1(n_14),
.B2(n_5),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_148),
.B1(n_156),
.B2(n_125),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_5),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_6),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_117),
.Y(n_181)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_103),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_140),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_196),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_117),
.B1(n_88),
.B2(n_94),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_184),
.B(n_204),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_103),
.B(n_96),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_179),
.B(n_181),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_SL g186 ( 
.A(n_129),
.B(n_108),
.C(n_123),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_123),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_95),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_197),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_119),
.CI(n_104),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_106),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_119),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_131),
.B(n_106),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_152),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_145),
.A2(n_108),
.B1(n_104),
.B2(n_86),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_147),
.B1(n_130),
.B2(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_107),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_133),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_107),
.B(n_130),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_207),
.A2(n_232),
.B1(n_234),
.B2(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_138),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_166),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_136),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_193),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_172),
.A2(n_136),
.B(n_163),
.C(n_144),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_184),
.B(n_182),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_229),
.B(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_162),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_137),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_160),
.B1(n_150),
.B2(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_172),
.A2(n_128),
.B1(n_155),
.B2(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_153),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_198),
.Y(n_263)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_132),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_199),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_168),
.B1(n_202),
.B2(n_188),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_184),
.B(n_175),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_261),
.B(n_214),
.Y(n_268)
);

AOI221xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_234),
.B1(n_212),
.B2(n_210),
.C(n_213),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_195),
.B1(n_168),
.B2(n_182),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_252),
.B1(n_260),
.B2(n_264),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_195),
.B1(n_203),
.B2(n_190),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_175),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_209),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_205),
.C(n_176),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_219),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_205),
.B1(n_176),
.B2(n_183),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_214),
.A2(n_200),
.B(n_198),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_209),
.B(n_230),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_229),
.C(n_233),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_266),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_177),
.B1(n_200),
.B2(n_165),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_222),
.B(n_171),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_222),
.A3(n_231),
.B1(n_224),
.B2(n_223),
.C1(n_221),
.C2(n_232),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_271),
.B(n_279),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_211),
.B1(n_223),
.B2(n_238),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_252),
.B1(n_247),
.B2(n_251),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_256),
.C(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_287),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_278),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_238),
.B(n_220),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_280),
.A2(n_282),
.B1(n_286),
.B2(n_245),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_243),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_228),
.B1(n_215),
.B2(n_227),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_235),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_237),
.B1(n_171),
.B2(n_193),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_164),
.B(n_240),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_251),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_244),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_266),
.C(n_246),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_282),
.C(n_273),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_242),
.B1(n_253),
.B2(n_263),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_293),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_294),
.A2(n_301),
.B1(n_305),
.B2(n_280),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_255),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_270),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_261),
.B1(n_255),
.B2(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_244),
.B1(n_245),
.B2(n_254),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_268),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_293),
.B(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_293),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_311),
.B(n_314),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_312),
.B(n_317),
.Y(n_330)
);

AOI321xp33_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_281),
.A3(n_277),
.B1(n_287),
.B2(n_289),
.C(n_270),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_296),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_288),
.C(n_276),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_321),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_318),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_272),
.C(n_278),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_283),
.B(n_254),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_295),
.B(n_293),
.C(n_307),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_265),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_303),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_301),
.B1(n_303),
.B2(n_298),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_325),
.A2(n_320),
.B1(n_321),
.B2(n_300),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_327),
.Y(n_340)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_331),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_298),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_311),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_330),
.A2(n_317),
.B(n_316),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_339),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_341),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_315),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_314),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_337),
.A2(n_331),
.B(n_323),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_344),
.A2(n_346),
.B(n_342),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_332),
.B1(n_324),
.B2(n_323),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_348),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_SL g346 ( 
.A1(n_343),
.A2(n_323),
.B(n_297),
.C(n_328),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_340),
.A2(n_297),
.B(n_328),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_341),
.B(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_351),
.B(n_354),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_353),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_347),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_356),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_355),
.B(n_352),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_346),
.Y(n_359)
);


endmodule