module real_jpeg_21578_n_17 (n_8, n_0, n_2, n_348, n_10, n_9, n_12, n_349, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_348;
input n_10;
input n_9;
input n_12;
input n_349;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_0),
.A2(n_22),
.B1(n_66),
.B2(n_67),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_0),
.A2(n_22),
.B1(n_49),
.B2(n_50),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_1),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_102),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_102),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_2),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_50),
.B(n_62),
.C(n_87),
.D(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_3),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_108),
.B(n_110),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_3),
.A2(n_32),
.B(n_43),
.C(n_144),
.D(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_3),
.B(n_32),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_3),
.B(n_36),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_31),
.B(n_33),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_125),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_107),
.Y(n_246)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_6),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_59),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_7),
.B(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_7),
.B(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_109),
.B1(n_155),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_8),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_10),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_90),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_11),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_156),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_156),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_156),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_341),
.B(n_344),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_76),
.B(n_340),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_20),
.B(n_37),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_20),
.B(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_20),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_26),
.B1(n_36),
.B2(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_23),
.A2(n_28),
.B(n_125),
.C(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_26),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_207),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_26),
.A2(n_34),
.B(n_36),
.Y(n_343)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_27),
.A2(n_30),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_27),
.A2(n_30),
.B1(n_215),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_27),
.A2(n_206),
.B(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_27),
.A2(n_30),
.B1(n_56),
.B2(n_290),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_30),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_30),
.A2(n_216),
.B(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_36),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_71),
.C(n_73),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_38),
.A2(n_39),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_54),
.C(n_60),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_40),
.A2(n_41),
.B1(n_60),
.B2(n_315),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_42),
.A2(n_52),
.B1(n_165),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_42),
.A2(n_201),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_42),
.A2(n_51),
.B1(n_52),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_48),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_43),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_43),
.A2(n_48),
.B1(n_243),
.B2(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_43),
.A2(n_48),
.B1(n_262),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_44),
.B(n_50),
.Y(n_152)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_47),
.A2(n_49),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_52),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_52),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_52),
.A2(n_166),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_54),
.A2(n_55),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_60),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_60),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_70),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_69),
.B1(n_101),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_61),
.A2(n_142),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_61),
.A2(n_69),
.B1(n_198),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_61),
.A2(n_69),
.B1(n_228),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_61),
.A2(n_69),
.B1(n_237),
.B2(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_62),
.A2(n_65),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx9p33_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_66),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_69),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_69),
.A2(n_103),
.B(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_70),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_71),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_333),
.B(n_339),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_306),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_348),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_254),
.A3(n_294),
.B1(n_300),
.B2(n_305),
.C(n_349),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_209),
.C(n_250),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_180),
.B(n_208),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_159),
.B(n_179),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_136),
.B(n_158),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_112),
.B(n_135),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_88),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_108),
.A2(n_119),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_108),
.A2(n_191),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_108),
.A2(n_119),
.B1(n_226),
.B2(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_108),
.A2(n_127),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_111),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_122),
.B(n_134),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_120),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_125),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_133),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_128),
.B(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_157),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_148),
.C(n_157),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_153),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_175),
.C(n_177),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_172),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_169),
.C(n_170),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_195),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_194),
.C(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_210),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_230),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_211),
.B(n_230),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.C(n_229),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_227),
.Y(n_239)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_248),
.B2(n_249),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_238),
.C(n_249),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_236),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_244),
.C(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_255),
.B(n_272),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.C(n_271),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_256),
.A2(n_257),
.B1(n_265),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_261),
.C(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_267),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_285),
.B(n_289),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_268),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_269),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_292),
.B2(n_293),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_284),
.C(n_293),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_282),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_280),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_281),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_282),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_308),
.B1(n_317),
.B2(n_330),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_319),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_319),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.C(n_318),
.Y(n_307)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_310),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_315),
.C(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_321),
.C(n_325),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_313),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_338),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_343),
.B(n_346),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);


endmodule