module fake_jpeg_29827_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_18),
.C(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_1),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_13),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_0),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_64),
.B(n_3),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_49),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_44),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_79),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_80),
.B(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_3),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_83),
.B1(n_7),
.B2(n_9),
.Y(n_90)
);

AO22x2_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_44),
.B1(n_21),
.B2(n_22),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_37),
.B(n_12),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_4),
.C(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_89),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_10),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_95),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_17),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.C(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_104),
.B1(n_97),
.B2(n_88),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_99),
.B(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_102),
.A3(n_90),
.B1(n_93),
.B2(n_98),
.C1(n_94),
.C2(n_26),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_102),
.Y(n_110)
);


endmodule