module fake_jpeg_17156_n_38 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_13),
.B1(n_9),
.B2(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_0),
.B2(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_18),
.B1(n_14),
.B2(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_21),
.B1(n_5),
.B2(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_24),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_23),
.Y(n_37)
);

NOR2x1_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_3),
.Y(n_38)
);


endmodule