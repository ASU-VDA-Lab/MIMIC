module fake_ariane_1359_n_1057 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1057);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1057;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_479;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_559;
wire n_331;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_715;
wire n_512;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_1044;
wire n_751;
wire n_1027;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_182),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_7),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_99),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_161),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_239),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_133),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_68),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_116),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_212),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_155),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_42),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_52),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_173),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_198),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_226),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_163),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_54),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_41),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_84),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_171),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_124),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_235),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_5),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_137),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_128),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_145),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_67),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_14),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_71),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_59),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_233),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_197),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_19),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_243),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_130),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_181),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_82),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_83),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_189),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_200),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_242),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_151),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_230),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_0),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_0),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_1),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_1),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

BUFx8_ASAP7_75t_SL g323 ( 
.A(n_276),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_2),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

CKINVDCx6p67_ASAP7_75t_R g328 ( 
.A(n_261),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_2),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_3),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_253),
.B(n_3),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_4),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_4),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_5),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_256),
.B(n_53),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_270),
.B(n_6),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_263),
.B(n_6),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_264),
.B(n_7),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_55),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_258),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_276),
.Y(n_347)
);

BUFx8_ASAP7_75t_SL g348 ( 
.A(n_284),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_267),
.B(n_8),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_275),
.B(n_8),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_9),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_255),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_316),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_278),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_L g360 ( 
.A1(n_340),
.A2(n_287),
.B1(n_312),
.B2(n_284),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_312),
.B1(n_287),
.B2(n_294),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_288),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_333),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_281),
.B1(n_255),
.B2(n_313),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_336),
.A2(n_281),
.B1(n_313),
.B2(n_290),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_340),
.A2(n_298),
.B1(n_304),
.B2(n_277),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_336),
.A2(n_308),
.B1(n_311),
.B2(n_305),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_315),
.A2(n_266),
.B1(n_268),
.B2(n_265),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_273),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_274),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_280),
.B1(n_283),
.B2(n_279),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_286),
.B1(n_289),
.B2(n_285),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_292),
.B1(n_295),
.B2(n_291),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

BUFx6f_ASAP7_75t_SL g379 ( 
.A(n_323),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_339),
.A2(n_299),
.B1(n_300),
.B2(n_296),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g383 ( 
.A1(n_329),
.A2(n_303),
.B1(n_306),
.B2(n_302),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_353),
.A2(n_309),
.B1(n_310),
.B2(n_307),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_12),
.Y(n_385)
);

AO22x2_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_13),
.Y(n_387)
);

OR2x6_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_15),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.B(n_16),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_17),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_18),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_19),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_337),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_318),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_R g398 ( 
.A1(n_321),
.A2(n_352),
.B1(n_348),
.B2(n_26),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_324),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_27),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_342),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_326),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

AND2x2_ASAP7_75t_SL g407 ( 
.A(n_361),
.B(n_320),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_320),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_404),
.A2(n_335),
.B(n_330),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_400),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_342),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_326),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_358),
.B(n_387),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_351),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_326),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_351),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_351),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_320),
.Y(n_424)
);

INVx3_ASAP7_75t_R g425 ( 
.A(n_379),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_394),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

OR2x6_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_320),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_367),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_381),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_379),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_405),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_368),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_365),
.B(n_355),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_361),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

NAND2x1p5_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_395),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_343),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_369),
.B(n_344),
.Y(n_446)
);

BUFx4f_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_327),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_360),
.B(n_355),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_365),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_355),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_386),
.B(n_349),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

INVx4_ASAP7_75t_SL g460 ( 
.A(n_405),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_383),
.B(n_327),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_375),
.B(n_349),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_402),
.B(n_28),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_399),
.B(n_345),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_358),
.B(n_325),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_358),
.B(n_325),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_345),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

NAND2x1p5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_325),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_410),
.A2(n_341),
.B(n_345),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_345),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_410),
.A2(n_341),
.B(n_345),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_30),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_30),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_345),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_31),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_432),
.B(n_424),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_407),
.B(n_345),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_420),
.B(n_341),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_341),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_31),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_448),
.B(n_32),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_32),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_414),
.B(n_341),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_452),
.B(n_33),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_426),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_414),
.B(n_341),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_33),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_445),
.B(n_341),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_341),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_430),
.B(n_314),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_437),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_460),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_427),
.B(n_314),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_466),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_415),
.B(n_454),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_462),
.A2(n_443),
.B(n_431),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_449),
.B(n_34),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_34),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_466),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_415),
.B(n_325),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_458),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_470),
.B(n_314),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_314),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_464),
.B(n_35),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_421),
.B(n_314),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_422),
.B(n_35),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_422),
.B(n_317),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_467),
.B(n_317),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_416),
.B(n_317),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_36),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_444),
.B(n_459),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_461),
.B(n_36),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_463),
.B(n_37),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_451),
.B(n_37),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_522),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_500),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_474),
.B(n_447),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_465),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_442),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_484),
.B(n_456),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_469),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_495),
.B(n_507),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_457),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_541),
.B(n_438),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_523),
.B(n_447),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_500),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_474),
.B(n_425),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_474),
.B(n_317),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_474),
.B(n_522),
.Y(n_569)
);

BUFx2_ASAP7_75t_SL g570 ( 
.A(n_517),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_492),
.B(n_317),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_531),
.B(n_38),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_495),
.B(n_38),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_495),
.B(n_39),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_482),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_486),
.B(n_39),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_528),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_507),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_496),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_487),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_488),
.B(n_325),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_317),
.Y(n_587)
);

NAND2x1_ASAP7_75t_SL g588 ( 
.A(n_536),
.B(n_40),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_486),
.B(n_40),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_494),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_507),
.B(n_41),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_527),
.B(n_42),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_531),
.B(n_43),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_497),
.B(n_44),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_528),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_527),
.B(n_44),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_497),
.B(n_45),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_497),
.B(n_45),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_492),
.B(n_46),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_482),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_46),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_519),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_503),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_574),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_566),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

INVx6_ASAP7_75t_L g611 ( 
.A(n_566),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_548),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_566),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_565),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_603),
.A2(n_536),
.B1(n_492),
.B2(n_544),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_565),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_593),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_528),
.Y(n_623)
);

BUFx4f_ASAP7_75t_SL g624 ( 
.A(n_576),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_557),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

BUFx2_ASAP7_75t_SL g629 ( 
.A(n_593),
.Y(n_629)
);

CKINVDCx6p67_ASAP7_75t_R g630 ( 
.A(n_564),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

BUFx2_ASAP7_75t_R g632 ( 
.A(n_551),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_574),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_555),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_582),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_590),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_568),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_547),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_515),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_568),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_593),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_555),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_560),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_560),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_577),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

CKINVDCx8_ASAP7_75t_R g649 ( 
.A(n_570),
.Y(n_649)
);

INVx6_ASAP7_75t_L g650 ( 
.A(n_568),
.Y(n_650)
);

BUFx2_ASAP7_75t_SL g651 ( 
.A(n_597),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_577),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_536),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_558),
.A2(n_544),
.B1(n_481),
.B2(n_543),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_589),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_605),
.Y(n_656)
);

NOR2x1_ASAP7_75t_SL g657 ( 
.A(n_584),
.B(n_505),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_584),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_548),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_582),
.Y(n_660)
);

INVx8_ASAP7_75t_L g661 ( 
.A(n_567),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_596),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_583),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_583),
.Y(n_665)
);

BUFx12f_ASAP7_75t_L g666 ( 
.A(n_589),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_589),
.B(n_542),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_600),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_607),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_652),
.A2(n_488),
.B1(n_538),
.B2(n_481),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_625),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_635),
.B(n_540),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_617),
.A2(n_481),
.B1(n_543),
.B2(n_542),
.Y(n_673)
);

CKINVDCx11_ASAP7_75t_R g674 ( 
.A(n_621),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_622),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_SL g676 ( 
.A1(n_643),
.A2(n_542),
.B1(n_543),
.B2(n_540),
.Y(n_676)
);

CKINVDCx11_ASAP7_75t_R g677 ( 
.A(n_621),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_642),
.A2(n_586),
.B(n_501),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_652),
.A2(n_488),
.B1(n_538),
.B2(n_540),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

CKINVDCx6p67_ASAP7_75t_R g681 ( 
.A(n_608),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_617),
.A2(n_525),
.B1(n_538),
.B2(n_534),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_654),
.A2(n_525),
.B1(n_534),
.B2(n_600),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_609),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_659),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_624),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_668),
.A2(n_525),
.B1(n_482),
.B2(n_597),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_635),
.A2(n_573),
.B1(n_575),
.B2(n_591),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_654),
.A2(n_580),
.B1(n_598),
.B2(n_595),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_610),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_615),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_608),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_643),
.A2(n_499),
.B1(n_597),
.B2(n_545),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_637),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_656),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_660),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_644),
.A2(n_645),
.B1(n_667),
.B2(n_668),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_SL g700 ( 
.A1(n_651),
.A2(n_599),
.B1(n_571),
.B2(n_526),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_613),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_653),
.A2(n_505),
.B1(n_501),
.B2(n_545),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_647),
.A2(n_520),
.B1(n_594),
.B2(n_572),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_628),
.A2(n_509),
.B(n_501),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_647),
.A2(n_520),
.B1(n_503),
.B2(n_592),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_666),
.A2(n_520),
.B1(n_606),
.B2(n_592),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_631),
.Y(n_708)
);

OAI21xp33_ASAP7_75t_SL g709 ( 
.A1(n_659),
.A2(n_588),
.B(n_480),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_649),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_665),
.Y(n_711)
);

OAI22x1_ASAP7_75t_SL g712 ( 
.A1(n_614),
.A2(n_624),
.B1(n_632),
.B2(n_612),
.Y(n_712)
);

INVx6_ASAP7_75t_L g713 ( 
.A(n_639),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_631),
.B(n_579),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_634),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_648),
.A2(n_526),
.B1(n_509),
.B2(n_485),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_636),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

INVx6_ASAP7_75t_L g719 ( 
.A(n_639),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_664),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_611),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_713),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_684),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_682),
.A2(n_666),
.B1(n_618),
.B2(n_655),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_713),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_694),
.A2(n_688),
.B1(n_676),
.B2(n_675),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_683),
.A2(n_649),
.B1(n_630),
.B2(n_659),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_672),
.B(n_699),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_682),
.A2(n_618),
.B1(n_630),
.B2(n_493),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_683),
.A2(n_526),
.B1(n_612),
.B2(n_640),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_673),
.A2(n_640),
.B1(n_490),
.B2(n_502),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_673),
.A2(n_493),
.B1(n_640),
.B2(n_485),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_698),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_687),
.A2(n_493),
.B1(n_485),
.B2(n_606),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_716),
.A2(n_491),
.B1(n_661),
.B2(n_524),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_670),
.A2(n_529),
.B1(n_623),
.B2(n_524),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_689),
.A2(n_679),
.B1(n_699),
.B2(n_700),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_690),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_710),
.B(n_631),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_703),
.A2(n_623),
.B1(n_472),
.B2(n_511),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_686),
.B(n_614),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_708),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_703),
.A2(n_706),
.B1(n_707),
.B2(n_671),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_709),
.A2(n_571),
.B1(n_491),
.B2(n_537),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_706),
.A2(n_623),
.B1(n_472),
.B2(n_511),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_611),
.Y(n_746)
);

OAI21xp33_ASAP7_75t_L g747 ( 
.A1(n_689),
.A2(n_539),
.B(n_513),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_707),
.A2(n_472),
.B1(n_515),
.B2(n_664),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_691),
.A2(n_661),
.B1(n_633),
.B2(n_631),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_692),
.B(n_611),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_702),
.A2(n_602),
.B1(n_579),
.B2(n_662),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_711),
.A2(n_472),
.B1(n_515),
.B2(n_550),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_674),
.A2(n_472),
.B1(n_556),
.B2(n_550),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_SL g754 ( 
.A1(n_680),
.A2(n_480),
.B(n_478),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_695),
.A2(n_571),
.B1(n_537),
.B2(n_633),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_685),
.A2(n_680),
.B1(n_681),
.B2(n_678),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_677),
.A2(n_472),
.B1(n_559),
.B2(n_556),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_697),
.A2(n_571),
.B1(n_633),
.B2(n_661),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_718),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_669),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_715),
.A2(n_472),
.B1(n_559),
.B2(n_571),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_721),
.B(n_504),
.Y(n_762)
);

OAI21xp33_ASAP7_75t_L g763 ( 
.A1(n_704),
.A2(n_539),
.B(n_513),
.Y(n_763)
);

OAI22x1_ASAP7_75t_SL g764 ( 
.A1(n_712),
.A2(n_633),
.B1(n_530),
.B2(n_638),
.Y(n_764)
);

BUFx12f_ASAP7_75t_L g765 ( 
.A(n_693),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_696),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_713),
.B(n_504),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_685),
.A2(n_602),
.B1(n_662),
.B2(n_663),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_705),
.B(n_627),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_717),
.A2(n_535),
.B1(n_627),
.B2(n_518),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_701),
.B(n_663),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_719),
.A2(n_530),
.B1(n_518),
.B2(n_701),
.Y(n_776)
);

INVx5_ASAP7_75t_SL g777 ( 
.A(n_708),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_719),
.B(n_530),
.Y(n_778)
);

OA222x2_ASAP7_75t_L g779 ( 
.A1(n_720),
.A2(n_535),
.B1(n_567),
.B2(n_628),
.C1(n_619),
.C2(n_587),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_719),
.A2(n_518),
.B1(n_512),
.B2(n_508),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_708),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_737),
.A2(n_508),
.B1(n_512),
.B2(n_604),
.Y(n_782)
);

OA21x2_ASAP7_75t_L g783 ( 
.A1(n_747),
.A2(n_533),
.B(n_532),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_726),
.A2(n_508),
.B1(n_512),
.B2(n_604),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_657),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_726),
.A2(n_604),
.B1(n_708),
.B2(n_518),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_738),
.B(n_714),
.Y(n_787)
);

OAI222xp33_ASAP7_75t_L g788 ( 
.A1(n_743),
.A2(n_714),
.B1(n_521),
.B2(n_477),
.C1(n_587),
.C2(n_567),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_728),
.A2(n_478),
.B1(n_521),
.B2(n_477),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_723),
.B(n_628),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_732),
.A2(n_735),
.B1(n_729),
.B2(n_730),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_750),
.B(n_733),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_735),
.A2(n_650),
.B1(n_619),
.B2(n_641),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_724),
.A2(n_477),
.B1(n_514),
.B2(n_587),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_740),
.A2(n_477),
.B1(n_514),
.B2(n_510),
.Y(n_795)
);

OA21x2_ASAP7_75t_L g796 ( 
.A1(n_763),
.A2(n_533),
.B(n_532),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_759),
.B(n_616),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_734),
.A2(n_736),
.B1(n_731),
.B2(n_760),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_727),
.A2(n_650),
.B1(n_514),
.B2(n_561),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_771),
.A2(n_514),
.B1(n_510),
.B2(n_650),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_745),
.A2(n_510),
.B1(n_584),
.B2(n_616),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_766),
.B(n_770),
.Y(n_802)
);

AOI221xp5_ASAP7_75t_L g803 ( 
.A1(n_762),
.A2(n_473),
.B1(n_479),
.B2(n_498),
.C(n_506),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_753),
.A2(n_510),
.B1(n_584),
.B2(n_616),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_757),
.A2(n_510),
.B1(n_626),
.B2(n_616),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_766),
.B(n_47),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_SL g807 ( 
.A1(n_776),
.A2(n_47),
.B(n_48),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_768),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_748),
.A2(n_626),
.B1(n_483),
.B2(n_489),
.Y(n_809)
);

NAND3xp33_ASAP7_75t_L g810 ( 
.A(n_756),
.B(n_626),
.C(n_638),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_773),
.A2(n_626),
.B1(n_483),
.B2(n_489),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_752),
.A2(n_498),
.B1(n_506),
.B2(n_561),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_778),
.B(n_479),
.C(n_473),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_767),
.B(n_638),
.Y(n_814)
);

AOI222xp33_ASAP7_75t_L g815 ( 
.A1(n_764),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.C1(n_51),
.C2(n_52),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_779),
.A2(n_658),
.B1(n_646),
.B2(n_641),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_772),
.A2(n_561),
.B1(n_546),
.B2(n_578),
.Y(n_817)
);

OA21x2_ASAP7_75t_L g818 ( 
.A1(n_754),
.A2(n_519),
.B(n_332),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_742),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_780),
.A2(n_658),
.B1(n_646),
.B2(n_641),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_775),
.A2(n_758),
.B1(n_765),
.B2(n_749),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_770),
.B(n_49),
.Y(n_822)
);

OAI221xp5_ASAP7_75t_L g823 ( 
.A1(n_744),
.A2(n_658),
.B1(n_646),
.B2(n_641),
.C(n_638),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_781),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_739),
.B(n_646),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_758),
.A2(n_581),
.B1(n_578),
.B2(n_546),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_749),
.A2(n_581),
.B1(n_578),
.B2(n_546),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_744),
.A2(n_581),
.B1(n_658),
.B2(n_519),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_755),
.A2(n_346),
.B1(n_334),
.B2(n_332),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_755),
.A2(n_346),
.B1(n_334),
.B2(n_332),
.Y(n_830)
);

OAI222xp33_ASAP7_75t_L g831 ( 
.A1(n_746),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.C1(n_57),
.C2(n_58),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_739),
.B(n_331),
.Y(n_832)
);

OAI222xp33_ASAP7_75t_L g833 ( 
.A1(n_722),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.C1(n_63),
.C2(n_64),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_802),
.B(n_742),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_832),
.A2(n_751),
.B(n_769),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_815),
.A2(n_741),
.B1(n_774),
.B2(n_725),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_785),
.B(n_742),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_785),
.B(n_742),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_819),
.B(n_777),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_806),
.B(n_777),
.Y(n_840)
);

OAI221xp5_ASAP7_75t_L g841 ( 
.A1(n_807),
.A2(n_782),
.B1(n_786),
.B2(n_821),
.C(n_791),
.Y(n_841)
);

AND4x1_ASAP7_75t_L g842 ( 
.A(n_810),
.B(n_761),
.C(n_777),
.D(n_69),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_L g843 ( 
.A(n_831),
.B(n_65),
.C(n_66),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_SL g844 ( 
.A1(n_799),
.A2(n_332),
.B(n_331),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_806),
.B(n_331),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_822),
.B(n_331),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_787),
.B(n_799),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_819),
.B(n_802),
.Y(n_848)
);

AOI211xp5_ASAP7_75t_L g849 ( 
.A1(n_833),
.A2(n_346),
.B(n_334),
.C(n_332),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_822),
.B(n_70),
.C(n_72),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_808),
.B(n_331),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_814),
.B(n_73),
.Y(n_852)
);

AOI221xp5_ASAP7_75t_L g853 ( 
.A1(n_798),
.A2(n_346),
.B1(n_334),
.B2(n_332),
.C(n_331),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_790),
.B(n_784),
.C(n_797),
.Y(n_854)
);

NAND4xp25_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_74),
.C(n_75),
.D(n_76),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_824),
.B(n_77),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_808),
.B(n_334),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_824),
.B(n_334),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_793),
.B(n_346),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_825),
.B(n_346),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_783),
.B(n_78),
.C(n_79),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_818),
.B(n_80),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_783),
.B(n_247),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_SL g864 ( 
.A1(n_828),
.A2(n_81),
.B(n_85),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_783),
.A2(n_789),
.B1(n_795),
.B2(n_794),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_783),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_827),
.B(n_86),
.Y(n_867)
);

OAI221xp5_ASAP7_75t_L g868 ( 
.A1(n_800),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_868)
);

OAI221xp5_ASAP7_75t_SL g869 ( 
.A1(n_829),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_SL g870 ( 
.A1(n_816),
.A2(n_95),
.B(n_96),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_796),
.B(n_97),
.C(n_98),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_796),
.B(n_246),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_796),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_818),
.B(n_100),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_823),
.B(n_102),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_796),
.B(n_103),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_818),
.B(n_813),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_801),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_818),
.B(n_107),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_811),
.A2(n_108),
.B(n_109),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_805),
.B(n_245),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_817),
.B(n_110),
.C(n_111),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_820),
.B(n_112),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_788),
.B(n_113),
.C(n_114),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_826),
.B(n_115),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_809),
.B(n_117),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_812),
.B(n_118),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_851),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_843),
.A2(n_804),
.B1(n_803),
.B2(n_122),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_855),
.B(n_120),
.C(n_121),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_848),
.B(n_123),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_851),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_834),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_847),
.B(n_125),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_873),
.A2(n_126),
.B(n_127),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_834),
.B(n_129),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_847),
.B(n_131),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_837),
.B(n_132),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_SL g901 ( 
.A1(n_841),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_901)
);

AOI221xp5_ASAP7_75t_L g902 ( 
.A1(n_836),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.C(n_141),
.Y(n_902)
);

AO22x1_ASAP7_75t_L g903 ( 
.A1(n_884),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_857),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_836),
.A2(n_880),
.B1(n_867),
.B2(n_885),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_838),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_867),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_870),
.A2(n_875),
.B1(n_885),
.B2(n_864),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_850),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_845),
.B(n_153),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_866),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_839),
.B(n_154),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_854),
.B(n_156),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_863),
.A2(n_157),
.B(n_158),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_877),
.B(n_160),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_840),
.Y(n_916)
);

NAND4xp75_ASAP7_75t_L g917 ( 
.A(n_883),
.B(n_162),
.C(n_164),
.D(n_165),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_849),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_846),
.B(n_172),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_883),
.A2(n_888),
.B1(n_852),
.B2(n_881),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_861),
.B(n_174),
.C(n_175),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_865),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_862),
.B(n_179),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_835),
.B(n_184),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_889),
.B(n_862),
.Y(n_925)
);

NOR2x1_ASAP7_75t_SL g926 ( 
.A(n_892),
.B(n_844),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_904),
.Y(n_927)
);

NAND4xp75_ASAP7_75t_SL g928 ( 
.A(n_898),
.B(n_852),
.C(n_888),
.D(n_874),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_911),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_915),
.B(n_872),
.Y(n_931)
);

XNOR2xp5_ASAP7_75t_L g932 ( 
.A(n_916),
.B(n_842),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_905),
.A2(n_865),
.B1(n_887),
.B2(n_886),
.Y(n_933)
);

NAND4xp75_ASAP7_75t_L g934 ( 
.A(n_908),
.B(n_876),
.C(n_856),
.D(n_853),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_920),
.B(n_913),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_915),
.B(n_860),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_911),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_894),
.B(n_879),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_906),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_893),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_889),
.B(n_859),
.Y(n_941)
);

NAND4xp75_ASAP7_75t_SL g942 ( 
.A(n_898),
.B(n_871),
.C(n_869),
.D(n_882),
.Y(n_942)
);

XOR2x2_ASAP7_75t_L g943 ( 
.A(n_905),
.B(n_868),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_891),
.A2(n_878),
.B1(n_187),
.B2(n_188),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_902),
.B(n_878),
.C(n_191),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_924),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_899),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_897),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_897),
.B(n_186),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_923),
.B(n_192),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_912),
.Y(n_952)
);

XOR2x2_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_932),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_929),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_929),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_943),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_935),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_930),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_949),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_927),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_940),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_949),
.B(n_923),
.Y(n_962)
);

XOR2xp5_ASAP7_75t_L g963 ( 
.A(n_928),
.B(n_900),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_947),
.B(n_896),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_939),
.B(n_937),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_944),
.A2(n_921),
.B1(n_895),
.B2(n_919),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_930),
.Y(n_967)
);

OA22x2_ASAP7_75t_L g968 ( 
.A1(n_957),
.A2(n_933),
.B1(n_952),
.B2(n_925),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_956),
.A2(n_935),
.B1(n_950),
.B2(n_946),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_954),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_962),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_963),
.A2(n_945),
.B1(n_931),
.B2(n_934),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_960),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_953),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_961),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_954),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_955),
.Y(n_977)
);

OAI22x1_ASAP7_75t_L g978 ( 
.A1(n_955),
.A2(n_939),
.B1(n_925),
.B2(n_938),
.Y(n_978)
);

XNOR2x1_ASAP7_75t_L g979 ( 
.A(n_953),
.B(n_942),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_973),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_973),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_975),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_975),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_971),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_979),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

OAI322xp33_ASAP7_75t_L g987 ( 
.A1(n_985),
.A2(n_956),
.A3(n_974),
.B1(n_968),
.B2(n_972),
.C1(n_964),
.C2(n_977),
.Y(n_987)
);

OA22x2_ASAP7_75t_L g988 ( 
.A1(n_985),
.A2(n_978),
.B1(n_970),
.B2(n_976),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

OA22x2_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_983),
.B1(n_984),
.B2(n_986),
.Y(n_990)
);

OA22x2_ASAP7_75t_L g991 ( 
.A1(n_981),
.A2(n_956),
.B1(n_964),
.B2(n_959),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_956),
.B1(n_969),
.B2(n_966),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_990),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_989),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_988),
.A2(n_967),
.B(n_958),
.C(n_922),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_987),
.A2(n_966),
.B1(n_959),
.B2(n_962),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_992),
.B(n_958),
.Y(n_997)
);

NOR2x1_ASAP7_75t_L g998 ( 
.A(n_993),
.B(n_965),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_996),
.A2(n_966),
.B1(n_890),
.B2(n_901),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_994),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_995),
.B(n_967),
.Y(n_1001)
);

NOR4xp25_ASAP7_75t_L g1002 ( 
.A(n_993),
.B(n_922),
.C(n_907),
.D(n_951),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_992),
.A2(n_966),
.B1(n_903),
.B2(n_907),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_965),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1001),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_1003),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_1004),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_1006),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1005),
.Y(n_1012)
);

NOR4xp25_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_1002),
.C(n_910),
.D(n_938),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_1005),
.B(n_909),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1009),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_1004),
.A2(n_918),
.B1(n_896),
.B2(n_925),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_1011),
.A2(n_930),
.B1(n_936),
.B2(n_917),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1010),
.A2(n_896),
.B1(n_914),
.B2(n_941),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1012),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1015),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1017),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1016),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1014),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1014),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1013),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1011),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1023),
.Y(n_1028)
);

OAI22x1_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_941),
.B1(n_926),
.B2(n_948),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1022),
.A2(n_914),
.B1(n_948),
.B2(n_944),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1024),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_1024),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1021),
.Y(n_1033)
);

AND4x2_ASAP7_75t_L g1034 ( 
.A(n_1020),
.B(n_196),
.C(n_199),
.D(n_201),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1026),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_1025),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1018),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_1019),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_1023),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1033),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1032),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_1037),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1036),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1040),
.A2(n_1038),
.B1(n_1030),
.B2(n_1035),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1043),
.A2(n_1029),
.B1(n_1039),
.B2(n_1032),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1044),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1046),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1048),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1047),
.Y(n_1052)
);

XNOR2xp5_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_1045),
.Y(n_1053)
);

AO22x2_ASAP7_75t_L g1054 ( 
.A1(n_1051),
.A2(n_1041),
.B1(n_1042),
.B2(n_1049),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1054),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1055),
.A2(n_1052),
.B1(n_1053),
.B2(n_231),
.C(n_232),
.Y(n_1056)
);

AOI211xp5_ASAP7_75t_L g1057 ( 
.A1(n_1056),
.A2(n_237),
.B(n_238),
.C(n_240),
.Y(n_1057)
);


endmodule