module real_aes_2081_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_753, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_752, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_753;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_752;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g151 ( .A(n_0), .B(n_125), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_1), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_2), .B(n_109), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_3), .B(n_127), .Y(n_444) );
INVx1_ASAP7_75t_L g116 ( .A(n_4), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_5), .B(n_109), .Y(n_178) );
NAND2xp33_ASAP7_75t_SL g221 ( .A(n_6), .B(n_115), .Y(n_221) );
INVx1_ASAP7_75t_L g213 ( .A(n_7), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_8), .Y(n_725) );
AND2x2_ASAP7_75t_L g176 ( .A(n_9), .B(n_133), .Y(n_176) );
AND2x2_ASAP7_75t_L g446 ( .A(n_10), .B(n_129), .Y(n_446) );
AND2x2_ASAP7_75t_L g456 ( .A(n_11), .B(n_219), .Y(n_456) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_13), .B(n_127), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_14), .Y(n_416) );
AOI221x1_ASAP7_75t_L g216 ( .A1(n_15), .A2(n_118), .B1(n_217), .B2(n_219), .C(n_220), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_16), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_17), .B(n_109), .Y(n_501) );
INVx1_ASAP7_75t_L g419 ( .A(n_18), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_19), .A2(n_87), .B1(n_109), .B2(n_162), .Y(n_460) );
AOI221xp5_ASAP7_75t_SL g140 ( .A1(n_20), .A2(n_36), .B1(n_109), .B2(n_118), .C(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_21), .A2(n_118), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_22), .B(n_125), .Y(n_181) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_23), .A2(n_86), .B(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g134 ( .A(n_23), .B(n_86), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_24), .B(n_127), .Y(n_126) );
INVxp67_ASAP7_75t_L g215 ( .A(n_25), .Y(n_215) );
AND2x2_ASAP7_75t_L g202 ( .A(n_26), .B(n_139), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_27), .A2(n_118), .B(n_150), .Y(n_149) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_28), .A2(n_219), .B(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_29), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_30), .B(n_127), .Y(n_142) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_31), .A2(n_99), .B1(n_719), .B2(n_729), .C1(n_741), .C2(n_745), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_31), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_31), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_32), .A2(n_118), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_33), .B(n_127), .Y(n_516) );
AND2x2_ASAP7_75t_L g115 ( .A(n_34), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g119 ( .A(n_34), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g170 ( .A(n_34), .Y(n_170) );
OR2x6_ASAP7_75t_L g417 ( .A(n_35), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_37), .B(n_109), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_38), .A2(n_78), .B1(n_118), .B2(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_39), .B(n_127), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_40), .B(n_109), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_41), .B(n_125), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_42), .A2(n_118), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g154 ( .A(n_43), .B(n_139), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_44), .B(n_125), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_45), .B(n_139), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_46), .B(n_109), .Y(n_493) );
INVx1_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVx1_ASAP7_75t_L g122 ( .A(n_47), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_48), .B(n_127), .Y(n_454) );
AND2x2_ASAP7_75t_L g483 ( .A(n_49), .B(n_139), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_50), .B(n_109), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_51), .B(n_125), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_52), .B(n_125), .Y(n_515) );
AND2x2_ASAP7_75t_L g193 ( .A(n_53), .B(n_139), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_54), .B(n_109), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_55), .B(n_127), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_56), .B(n_109), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_57), .A2(n_118), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_58), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_59), .B(n_125), .Y(n_190) );
AND2x2_ASAP7_75t_L g507 ( .A(n_60), .B(n_133), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_61), .A2(n_118), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_62), .B(n_127), .Y(n_182) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_63), .B(n_129), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_64), .B(n_125), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_65), .B(n_125), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_66), .A2(n_89), .B1(n_118), .B2(n_168), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_67), .B(n_127), .Y(n_504) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
INVx1_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_69), .B(n_125), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_70), .A2(n_100), .B1(n_708), .B2(n_709), .C1(n_715), .C2(n_718), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_70), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_71), .A2(n_118), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_72), .A2(n_118), .B(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_73), .A2(n_118), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g518 ( .A(n_74), .B(n_133), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_75), .B(n_139), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_76), .A2(n_80), .B1(n_109), .B2(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_77), .B(n_109), .Y(n_191) );
INVx1_ASAP7_75t_L g420 ( .A(n_79), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_81), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_82), .B(n_125), .Y(n_143) );
AND2x2_ASAP7_75t_L g437 ( .A(n_83), .B(n_129), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_84), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_85), .A2(n_118), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_88), .B(n_127), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_90), .A2(n_118), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_91), .B(n_127), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_92), .B(n_109), .Y(n_153) );
INVxp67_ASAP7_75t_L g218 ( .A(n_93), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_94), .B(n_127), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_95), .A2(n_118), .B(n_123), .Y(n_117) );
BUFx2_ASAP7_75t_L g506 ( .A(n_96), .Y(n_506) );
BUFx2_ASAP7_75t_L g726 ( .A(n_97), .Y(n_726) );
BUFx2_ASAP7_75t_SL g749 ( .A(n_97), .Y(n_749) );
AOI22xp5_ASAP7_75t_SL g100 ( .A1(n_101), .A2(n_415), .B1(n_421), .B2(n_705), .Y(n_100) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_101), .A2(n_421), .B1(n_711), .B2(n_714), .Y(n_710) );
INVx3_ASAP7_75t_SL g733 ( .A(n_101), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_101), .Y(n_734) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_307), .Y(n_101) );
NOR3xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_235), .C(n_285), .Y(n_102) );
OAI211xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_155), .B(n_203), .C(n_224), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_135), .Y(n_104) );
AND2x2_ASAP7_75t_L g234 ( .A(n_105), .B(n_136), .Y(n_234) );
INVx1_ASAP7_75t_L g365 ( .A(n_105), .Y(n_365) );
NOR2x1p5_ASAP7_75t_L g397 ( .A(n_105), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g208 ( .A(n_106), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g256 ( .A(n_106), .Y(n_256) );
OR2x2_ASAP7_75t_L g260 ( .A(n_106), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_106), .B(n_138), .Y(n_272) );
OR2x2_ASAP7_75t_L g294 ( .A(n_106), .B(n_138), .Y(n_294) );
AND2x4_ASAP7_75t_L g300 ( .A(n_106), .B(n_264), .Y(n_300) );
OR2x2_ASAP7_75t_L g317 ( .A(n_106), .B(n_210), .Y(n_317) );
INVx1_ASAP7_75t_L g352 ( .A(n_106), .Y(n_352) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_106), .Y(n_374) );
OR2x2_ASAP7_75t_L g388 ( .A(n_106), .B(n_321), .Y(n_388) );
AND2x4_ASAP7_75t_SL g392 ( .A(n_106), .B(n_210), .Y(n_392) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_132), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_117), .B(n_129), .Y(n_107) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_115), .Y(n_109) );
INVx1_ASAP7_75t_L g222 ( .A(n_110), .Y(n_222) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
AND2x6_ASAP7_75t_L g125 ( .A(n_111), .B(n_120), .Y(n_125) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g127 ( .A(n_113), .B(n_122), .Y(n_127) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx5_ASAP7_75t_L g128 ( .A(n_115), .Y(n_128) );
AND2x2_ASAP7_75t_L g121 ( .A(n_116), .B(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx3_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
INVx2_ASAP7_75t_L g172 ( .A(n_120), .Y(n_172) );
AND2x4_ASAP7_75t_L g168 ( .A(n_121), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B(n_128), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_125), .B(n_506), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_128), .A2(n_142), .B(n_143), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_128), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_128), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_128), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_128), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_128), .A2(n_435), .B(n_436), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_128), .A2(n_443), .B(n_444), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_128), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_128), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_128), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_128), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_128), .A2(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_SL g159 ( .A(n_129), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_129), .A2(n_501), .B(n_502), .Y(n_500) );
BUFx4f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_L g147 ( .A(n_130), .Y(n_147) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_131), .B(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g183 ( .A(n_131), .B(n_134), .Y(n_183) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g344 ( .A(n_136), .B(n_300), .Y(n_344) );
AND2x2_ASAP7_75t_L g391 ( .A(n_136), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_145), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g207 ( .A(n_138), .Y(n_207) );
AND2x2_ASAP7_75t_L g254 ( .A(n_138), .B(n_145), .Y(n_254) );
INVx2_ASAP7_75t_L g261 ( .A(n_138), .Y(n_261) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_138), .Y(n_382) );
BUFx3_ASAP7_75t_L g398 ( .A(n_138), .Y(n_398) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_144), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_139), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_139), .A2(n_432), .B(n_433), .Y(n_431) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_139), .A2(n_460), .B(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_145), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g321 ( .A(n_145), .B(n_261), .Y(n_321) );
INVx1_ASAP7_75t_L g339 ( .A(n_145), .Y(n_339) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_145), .Y(n_355) );
INVx1_ASAP7_75t_L g377 ( .A(n_145), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_145), .B(n_256), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_145), .B(n_210), .Y(n_414) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_154), .Y(n_146) );
INVx4_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_147), .A2(n_450), .B(n_456), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_174), .Y(n_156) );
AND2x4_ASAP7_75t_L g228 ( .A(n_157), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g239 ( .A(n_157), .Y(n_239) );
AND2x2_ASAP7_75t_L g244 ( .A(n_157), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g279 ( .A(n_157), .B(n_184), .Y(n_279) );
AND2x2_ASAP7_75t_L g289 ( .A(n_157), .B(n_185), .Y(n_289) );
OR2x2_ASAP7_75t_L g369 ( .A(n_157), .B(n_284), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g399 ( .A1(n_157), .A2(n_312), .A3(n_351), .B1(n_384), .B2(n_400), .C1(n_401), .C2(n_402), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_157), .B(n_382), .Y(n_400) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g233 ( .A(n_158), .Y(n_233) );
AOI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_173), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_167), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_162), .A2(n_168), .B1(n_212), .B2(n_214), .Y(n_211) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_166), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2x1p5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_174), .A2(n_346), .B1(n_350), .B2(n_353), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_174), .A2(n_406), .B(n_407), .C(n_410), .Y(n_405) );
AND2x4_ASAP7_75t_SL g174 ( .A(n_175), .B(n_184), .Y(n_174) );
AND2x4_ASAP7_75t_L g227 ( .A(n_175), .B(n_195), .Y(n_227) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_175), .Y(n_231) );
INVx5_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
INVx2_ASAP7_75t_L g252 ( .A(n_175), .Y(n_252) );
AND2x2_ASAP7_75t_L g275 ( .A(n_175), .B(n_185), .Y(n_275) );
AND2x2_ASAP7_75t_L g304 ( .A(n_175), .B(n_194), .Y(n_304) );
OR2x2_ASAP7_75t_L g313 ( .A(n_175), .B(n_233), .Y(n_313) );
OR2x2_ASAP7_75t_L g328 ( .A(n_175), .B(n_242), .Y(n_328) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_183), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_183), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_183), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_183), .B(n_218), .Y(n_217) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_183), .B(n_221), .C(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_183), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_183), .A2(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_184), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_SL g312 ( .A(n_184), .Y(n_312) );
AND2x2_ASAP7_75t_L g335 ( .A(n_184), .B(n_243), .Y(n_335) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_194), .Y(n_184) );
INVx2_ASAP7_75t_L g229 ( .A(n_185), .Y(n_229) );
AND2x2_ASAP7_75t_L g232 ( .A(n_185), .B(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g246 ( .A(n_185), .B(n_195), .Y(n_246) );
INVx1_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_185), .B(n_195), .Y(n_284) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_185), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_185), .B(n_243), .Y(n_359) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_192), .A2(n_196), .B(n_202), .Y(n_195) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_192), .A2(n_196), .B(n_202), .Y(n_242) );
AOI21x1_ASAP7_75t_L g439 ( .A1(n_192), .A2(n_440), .B(n_446), .Y(n_439) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_195), .Y(n_265) );
AND2x2_ASAP7_75t_L g349 ( .A(n_195), .B(n_233), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_201), .Y(n_196) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_205), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x6_ASAP7_75t_SL g413 ( .A(n_206), .B(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_207), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_207), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g361 ( .A(n_207), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_208), .A2(n_270), .B1(n_273), .B2(n_280), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_209), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g305 ( .A(n_209), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_209), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_209), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_223), .Y(n_209) );
AND2x2_ASAP7_75t_L g255 ( .A(n_210), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g264 ( .A(n_210), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_210), .A2(n_271), .B1(n_323), .B2(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g330 ( .A(n_210), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_210), .B(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_210), .B(n_254), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_210), .B(n_261), .Y(n_403) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_216), .Y(n_210) );
INVx3_ASAP7_75t_L g511 ( .A(n_219), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_230), .B(n_234), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
NAND4xp25_ASAP7_75t_SL g273 ( .A(n_226), .B(n_274), .C(n_276), .D(n_278), .Y(n_273) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_227), .B(n_334), .Y(n_363) );
AND2x2_ASAP7_75t_L g390 ( .A(n_227), .B(n_228), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_227), .B(n_250), .Y(n_401) );
INVx1_ASAP7_75t_L g266 ( .A(n_228), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_228), .A2(n_291), .B1(n_302), .B2(n_305), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_228), .B(n_241), .C(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_228), .B(n_243), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_228), .B(n_251), .Y(n_394) );
AND2x2_ASAP7_75t_L g326 ( .A(n_229), .B(n_233), .Y(n_326) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_229), .Y(n_387) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g282 ( .A(n_231), .Y(n_282) );
INVx1_ASAP7_75t_L g372 ( .A(n_232), .Y(n_372) );
AND2x2_ASAP7_75t_L g379 ( .A(n_232), .B(n_243), .Y(n_379) );
BUFx2_ASAP7_75t_L g334 ( .A(n_233), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g235 ( .A(n_236), .B(n_257), .C(n_269), .Y(n_235) );
OAI31xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_244), .A3(n_247), .B(n_253), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_237), .A2(n_291), .B1(n_295), .B2(n_296), .Y(n_290) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
OR2x2_ASAP7_75t_L g276 ( .A(n_239), .B(n_277), .Y(n_276) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_239), .B(n_303), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_240), .A2(n_342), .B(n_372), .C(n_373), .Y(n_371) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_241), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_242), .B(n_250), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_242), .B(n_275), .Y(n_295) );
AND2x2_ASAP7_75t_L g412 ( .A(n_245), .B(n_334), .Y(n_412) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_252), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_251), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g343 ( .A(n_251), .B(n_326), .Y(n_343) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_252), .B(n_326), .Y(n_332) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g324 ( .A(n_254), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_255), .B(n_355), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_265), .A3(n_266), .B1(n_267), .B2(n_752), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_258), .A2(n_343), .B1(n_379), .B2(n_380), .C(n_383), .Y(n_378) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_261), .Y(n_306) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g271 ( .A(n_263), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g376 ( .A(n_264), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_265), .B(n_287), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_267), .A2(n_310), .B1(n_314), .B2(n_318), .C(n_322), .Y(n_309) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI211xp5_ASAP7_75t_L g285 ( .A1(n_272), .A2(n_286), .B(n_290), .C(n_301), .Y(n_285) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_278), .A2(n_288), .A3(n_337), .B1(n_384), .B2(n_385), .C1(n_386), .C2(n_388), .Y(n_383) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_281), .A2(n_411), .B(n_413), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g367 ( .A1(n_287), .A2(n_368), .B(n_370), .C(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g409 ( .A(n_294), .B(n_375), .Y(n_409) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_300), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g384 ( .A(n_300), .Y(n_384) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI31xp33_ASAP7_75t_L g340 ( .A1(n_304), .A2(n_341), .A3(n_343), .B(n_344), .Y(n_340) );
NOR2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_366), .Y(n_307) );
NAND5xp2_ASAP7_75t_L g308 ( .A(n_309), .B(n_329), .C(n_340), .D(n_345), .E(n_356), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_312), .A2(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_333), .C(n_336), .Y(n_329) );
INVxp33_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g358 ( .A(n_334), .B(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_337), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_358), .A2(n_363), .B(n_364), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_378), .C(n_389), .D(n_405), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_376), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g406 ( .A(n_388), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_393), .B2(n_395), .C(n_399), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_415), .Y(n_713) );
AND2x6_ASAP7_75t_SL g415 ( .A(n_416), .B(n_417), .Y(n_415) );
OR2x6_ASAP7_75t_SL g706 ( .A(n_416), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g717 ( .A(n_416), .B(n_417), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_416), .B(n_707), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_417), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_618), .Y(n_421) );
NOR4xp75_ASAP7_75t_L g422 ( .A(n_423), .B(n_541), .C(n_566), .D(n_593), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_478), .B(n_519), .Y(n_423) );
NOR4xp25_ASAP7_75t_L g424 ( .A(n_425), .B(n_462), .C(n_469), .D(n_473), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_447), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_438), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_429), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_429), .B(n_466), .Y(n_612) );
AND2x2_ASAP7_75t_L g637 ( .A(n_429), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g662 ( .A(n_429), .B(n_457), .Y(n_662) );
AND2x2_ASAP7_75t_L g703 ( .A(n_429), .B(n_471), .Y(n_703) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_SL g475 ( .A(n_430), .B(n_468), .Y(n_475) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_449), .Y(n_477) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_430), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g538 ( .A(n_430), .Y(n_538) );
AND2x2_ASAP7_75t_L g544 ( .A(n_430), .B(n_471), .Y(n_544) );
BUFx2_ASAP7_75t_L g557 ( .A(n_430), .Y(n_557) );
AND2x4_ASAP7_75t_L g588 ( .A(n_430), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g635 ( .A(n_430), .B(n_636), .Y(n_635) );
OR2x6_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g629 ( .A(n_438), .Y(n_629) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g468 ( .A(n_439), .Y(n_468) );
AND2x2_ASAP7_75t_L g471 ( .A(n_439), .B(n_449), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_447), .B(n_647), .Y(n_700) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g537 ( .A(n_448), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_457), .Y(n_448) );
INVx2_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
INVx2_ASAP7_75t_L g528 ( .A(n_449), .Y(n_528) );
AND2x2_ASAP7_75t_L g638 ( .A(n_449), .B(n_468), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .Y(n_450) );
INVx2_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
BUFx3_ASAP7_75t_L g543 ( .A(n_457), .Y(n_543) );
AND2x2_ASAP7_75t_L g570 ( .A(n_457), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x4_ASAP7_75t_L g464 ( .A(n_458), .B(n_459), .Y(n_464) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx2_ASAP7_75t_L g472 ( .A(n_463), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_463), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g641 ( .A(n_463), .B(n_581), .Y(n_641) );
AND2x2_ASAP7_75t_L g665 ( .A(n_463), .B(n_475), .Y(n_665) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g561 ( .A(n_464), .B(n_467), .Y(n_561) );
AND2x2_ASAP7_75t_L g643 ( .A(n_464), .B(n_636), .Y(n_643) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g686 ( .A(n_466), .Y(n_686) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g571 ( .A(n_467), .Y(n_571) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_468), .Y(n_575) );
INVx2_ASAP7_75t_L g583 ( .A(n_468), .Y(n_583) );
INVx1_ASAP7_75t_L g589 ( .A(n_468), .Y(n_589) );
AOI222xp33_ASAP7_75t_SL g519 ( .A1(n_469), .A2(n_520), .B1(n_524), .B2(n_529), .C1(n_536), .C2(n_539), .Y(n_519) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g596 ( .A(n_471), .Y(n_596) );
BUFx2_ASAP7_75t_L g625 ( .A(n_471), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_472), .A2(n_620), .B(n_624), .C(n_632), .Y(n_619) );
OR2x2_ASAP7_75t_L g690 ( .A(n_472), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g698 ( .A(n_472), .B(n_603), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_475), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g673 ( .A(n_475), .B(n_561), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_475), .B(n_653), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_476), .B(n_543), .Y(n_681) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g603 ( .A(n_477), .B(n_575), .Y(n_603) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_498), .Y(n_479) );
INVx1_ASAP7_75t_L g697 ( .A(n_480), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
AND2x2_ASAP7_75t_L g540 ( .A(n_481), .B(n_499), .Y(n_540) );
INVx1_ASAP7_75t_L g617 ( .A(n_481), .Y(n_617) );
OR2x2_ASAP7_75t_L g676 ( .A(n_481), .B(n_499), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_481), .B(n_548), .Y(n_682) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g523 ( .A(n_482), .Y(n_523) );
OR2x2_ASAP7_75t_L g555 ( .A(n_482), .B(n_509), .Y(n_555) );
AND2x2_ASAP7_75t_L g564 ( .A(n_482), .B(n_491), .Y(n_564) );
NAND2x1_ASAP7_75t_L g592 ( .A(n_482), .B(n_499), .Y(n_592) );
AND2x2_ASAP7_75t_L g639 ( .A(n_482), .B(n_534), .Y(n_639) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g522 ( .A(n_491), .Y(n_522) );
INVx1_ASAP7_75t_L g532 ( .A(n_491), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_491), .B(n_535), .Y(n_548) );
INVx2_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
OR2x2_ASAP7_75t_L g649 ( .A(n_491), .B(n_499), .Y(n_649) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
NOR2x1_ASAP7_75t_SL g534 ( .A(n_499), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g552 ( .A(n_499), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g565 ( .A(n_499), .B(n_509), .Y(n_565) );
BUFx2_ASAP7_75t_L g584 ( .A(n_499), .Y(n_584) );
INVx2_ASAP7_75t_SL g611 ( .A(n_499), .Y(n_611) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_507), .Y(n_499) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g521 ( .A(n_509), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g667 ( .A(n_509), .B(n_609), .Y(n_667) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_510) );
AO21x1_ASAP7_75t_SL g535 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_520), .A2(n_544), .B(n_684), .C(n_688), .Y(n_683) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_521), .B(n_599), .Y(n_634) );
BUFx2_ASAP7_75t_L g598 ( .A(n_522), .Y(n_598) );
OR2x2_ASAP7_75t_L g546 ( .A(n_523), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g631 ( .A(n_523), .B(n_565), .Y(n_631) );
AND2x2_ASAP7_75t_L g652 ( .A(n_523), .B(n_608), .Y(n_652) );
INVx2_ASAP7_75t_L g659 ( .A(n_523), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_524), .A2(n_665), .B(n_666), .Y(n_664) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND2x2_ASAP7_75t_L g606 ( .A(n_525), .B(n_588), .Y(n_606) );
OR2x2_ASAP7_75t_L g685 ( .A(n_525), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_526), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_528), .Y(n_559) );
AND2x2_ASAP7_75t_L g636 ( .A(n_528), .B(n_583), .Y(n_636) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g621 ( .A(n_531), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_SL g630 ( .A(n_531), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_531), .B(n_540), .Y(n_663) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g539 ( .A(n_532), .B(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g658 ( .A(n_533), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g608 ( .A(n_534), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g578 ( .A(n_535), .B(n_553), .Y(n_578) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_536), .A2(n_586), .A3(n_588), .B(n_590), .Y(n_585) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_538), .B(n_561), .Y(n_587) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
OR2x2_ASAP7_75t_L g597 ( .A(n_543), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g702 ( .A(n_543), .Y(n_702) );
INVx2_ASAP7_75t_SL g687 ( .A(n_544), .Y(n_687) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g591 ( .A(n_547), .B(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g675 ( .A(n_547), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_548), .B(n_611), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_556), .B1(n_560), .B2(n_562), .Y(n_549) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_550), .A2(n_669), .B(n_670), .Y(n_668) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g609 ( .A(n_553), .Y(n_609) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g623 ( .A(n_555), .B(n_584), .Y(n_623) );
OR2x2_ASAP7_75t_L g648 ( .A(n_555), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_557), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_557), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g647 ( .A(n_557), .Y(n_647) );
INVx2_ASAP7_75t_L g576 ( .A(n_558), .Y(n_576) );
INVx1_ASAP7_75t_L g656 ( .A(n_559), .Y(n_656) );
AND2x2_ASAP7_75t_L g579 ( .A(n_561), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g653 ( .A(n_561), .Y(n_653) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_567), .B(n_585), .Y(n_566) );
OAI321xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .A3(n_577), .B1(n_578), .B2(n_579), .C(n_584), .Y(n_567) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_568), .A2(n_599), .A3(n_694), .B1(n_696), .B2(n_698), .C1(n_699), .C2(n_704), .Y(n_693) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g646 ( .A(n_571), .Y(n_646) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_573), .B(n_653), .Y(n_670) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g678 ( .A(n_576), .Y(n_678) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_578), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI21xp33_ASAP7_75t_SL g677 ( .A1(n_581), .A2(n_587), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx3_ASAP7_75t_L g599 ( .A(n_592), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_613), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B1(n_600), .B2(n_601), .C(n_604), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
AND2x2_ASAP7_75t_L g600 ( .A(n_598), .B(n_599), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B1(n_610), .B2(n_612), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g616 ( .A(n_608), .B(n_617), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_611), .A2(n_700), .B(n_701), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g618 ( .A(n_619), .B(n_650), .C(n_671), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_623), .A2(n_658), .B1(n_685), .B2(n_687), .Y(n_684) );
OAI21xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_630), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_625), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_631), .A2(n_673), .B1(n_674), .B2(n_677), .C(n_679), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_639), .C(n_640), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g669 ( .A(n_635), .Y(n_669) );
INVx1_ASAP7_75t_L g691 ( .A(n_636), .Y(n_691) );
INVx1_ASAP7_75t_SL g689 ( .A(n_637), .Y(n_689) );
AOI31xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .A3(n_644), .B(n_648), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_641), .A2(n_651), .B1(n_653), .B2(n_654), .C(n_753), .Y(n_650) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_668), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g666 ( .A(n_659), .B(n_667), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g695 ( .A(n_667), .Y(n_695) );
BUFx2_ASAP7_75t_SL g704 ( .A(n_667), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_683), .C(n_693), .Y(n_671) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_682), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_692), .Y(n_688) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g714 ( .A(n_705), .Y(n_714) );
CKINVDCx11_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx4_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_727), .Y(n_720) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_726), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_SL g744 ( .A(n_724), .B(n_726), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_724), .A2(n_747), .B(n_750), .Y(n_746) );
BUFx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
BUFx2_ASAP7_75t_L g736 ( .A(n_728), .Y(n_736) );
BUFx3_ASAP7_75t_L g739 ( .A(n_728), .Y(n_739) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_735), .B(n_737), .Y(n_730) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g750 ( .A(n_736), .Y(n_750) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_740), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx9p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
CKINVDCx8_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
endmodule