module fake_aes_543_n_690 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_690);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_690;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g78 ( .A(n_41), .Y(n_78) );
BUFx6f_ASAP7_75t_SL g79 ( .A(n_34), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_19), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_5), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_35), .B(n_31), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_70), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_51), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_74), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_76), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_77), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_50), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_38), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_0), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_71), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_6), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_65), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_14), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_37), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_18), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_46), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_64), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_33), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_63), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_23), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_30), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_62), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_22), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_25), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_32), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
NOR2xp67_ASAP7_75t_L g118 ( .A(n_18), .B(n_17), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_67), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_56), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_45), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_16), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_104), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_119), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_89), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_119), .B(n_1), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_111), .Y(n_133) );
NOR2x1_ASAP7_75t_L g134 ( .A(n_100), .B(n_1), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_85), .B(n_2), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_103), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_87), .B(n_27), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_88), .B(n_28), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g143 ( .A(n_79), .B(n_75), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_81), .B(n_4), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_104), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_85), .B(n_6), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_121), .B(n_7), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_83), .B(n_7), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_93), .B(n_8), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_93), .B(n_8), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_96), .B(n_124), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_83), .B(n_9), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_108), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_101), .B(n_9), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_98), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_97), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_98), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_164), .Y(n_172) );
NAND2xp33_ASAP7_75t_SL g173 ( .A(n_151), .B(n_79), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_164), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
AND2x6_ASAP7_75t_L g176 ( .A(n_128), .B(n_115), .Y(n_176) );
INVx6_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_164), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_130), .B(n_105), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_155), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_164), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_128), .A2(n_113), .B1(n_114), .B2(n_97), .Y(n_186) );
INVx5_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_132), .B(n_82), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_130), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_141), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_133), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_168), .B(n_101), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_132), .B(n_115), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_126), .B(n_86), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_126), .B(n_91), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_168), .B(n_113), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
OR2x6_ASAP7_75t_L g207 ( .A(n_136), .B(n_118), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_136), .B(n_114), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_135), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_131), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_151), .B(n_105), .Y(n_211) );
AO22x2_ASAP7_75t_L g212 ( .A1(n_129), .A2(n_124), .B1(n_82), .B2(n_109), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_154), .B(n_107), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_129), .B(n_86), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_139), .B(n_106), .Y(n_215) );
INVx8_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_139), .B(n_116), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_137), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_142), .B(n_102), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_146), .B(n_125), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_138), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_146), .B(n_99), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_148), .B(n_102), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_148), .B(n_110), .Y(n_227) );
NAND3x1_ASAP7_75t_L g228 ( .A(n_137), .B(n_123), .C(n_122), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_208), .B(n_165), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_199), .B(n_152), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_176), .A2(n_162), .B1(n_140), .B2(n_138), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_221), .B(n_169), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_200), .B(n_152), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_227), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_208), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_226), .B(n_169), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_192), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_219), .A2(n_150), .B1(n_157), .B2(n_160), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_218), .B(n_166), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_170), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_190), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_181), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_226), .B(n_167), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_217), .B(n_167), .Y(n_248) );
OAI221xp5_ASAP7_75t_L g249 ( .A1(n_186), .A2(n_160), .B1(n_150), .B2(n_157), .C(n_166), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_216), .Y(n_251) );
CKINVDCx11_ASAP7_75t_R g252 ( .A(n_193), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_176), .A2(n_196), .B1(n_208), .B2(n_212), .Y(n_253) );
AO22x1_ASAP7_75t_L g254 ( .A1(n_176), .A2(n_140), .B1(n_138), .B2(n_162), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_218), .B(n_161), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_208), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_197), .B(n_156), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_176), .A2(n_162), .B1(n_140), .B2(n_165), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_194), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_172), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_182), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_176), .A2(n_163), .B1(n_162), .B2(n_143), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_184), .B(n_163), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_206), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_205), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_174), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_218), .B(n_161), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_176), .A2(n_162), .B1(n_143), .B2(n_153), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_174), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_206), .Y(n_277) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_190), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_214), .B(n_156), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_190), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_182), .B(n_153), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_205), .A2(n_224), .B(n_222), .C(n_198), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_211), .B(n_162), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_176), .A2(n_196), .B1(n_212), .B2(n_205), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_180), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_183), .B(n_78), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_184), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_211), .B(n_162), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_180), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_205), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_203), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_239), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_289), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_239), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_245), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_229), .A2(n_196), .B1(n_212), .B2(n_219), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_240), .B(n_191), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_244), .B(n_222), .Y(n_301) );
OR2x6_ASAP7_75t_L g302 ( .A(n_272), .B(n_213), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_278), .A2(n_183), .B1(n_196), .B2(n_189), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_229), .B(n_213), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_253), .A2(n_213), .B1(n_212), .B2(n_228), .Y(n_305) );
BUFx4_ASAP7_75t_SL g306 ( .A(n_260), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_281), .B(n_195), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_266), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_252), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_285), .A2(n_228), .B1(n_203), .B2(n_204), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_245), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_272), .B(n_216), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_252), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_229), .A2(n_196), .B1(n_173), .B2(n_224), .Y(n_316) );
CKINVDCx6p67_ASAP7_75t_R g317 ( .A(n_231), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_292), .B(n_195), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_292), .B(n_196), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
AO21x1_ASAP7_75t_L g321 ( .A1(n_241), .A2(n_127), .B(n_145), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_268), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_238), .B(n_196), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_237), .B(n_222), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_263), .B(n_203), .Y(n_325) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_284), .B(n_204), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_257), .B(n_224), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_283), .A2(n_179), .B(n_195), .C(n_207), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_260), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_247), .B(n_195), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g332 ( .A(n_275), .B(n_204), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_267), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_271), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_279), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_267), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_243), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_216), .B(n_187), .Y(n_340) );
BUFx2_ASAP7_75t_SL g341 ( .A(n_251), .Y(n_341) );
AND2x6_ASAP7_75t_L g342 ( .A(n_243), .B(n_134), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_279), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_230), .B(n_215), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
NOR2x1_ASAP7_75t_SL g346 ( .A(n_341), .B(n_251), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_305), .A2(n_194), .B1(n_249), .B2(n_287), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_335), .A2(n_207), .B1(n_235), .B2(n_236), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_294), .Y(n_350) );
INVx8_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_328), .A2(n_274), .B(n_255), .C(n_258), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_299), .A2(n_265), .B1(n_277), .B2(n_259), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_300), .A2(n_207), .B1(n_248), .B2(n_280), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_301), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_207), .B1(n_233), .B2(n_220), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_301), .B(n_277), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_316), .A2(n_234), .B1(n_232), .B2(n_251), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_315), .A2(n_140), .B1(n_79), .B2(n_288), .Y(n_361) );
OAI22xp33_ASAP7_75t_SL g362 ( .A1(n_302), .A2(n_134), .B1(n_120), .B2(n_117), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_316), .A2(n_288), .B1(n_245), .B2(n_250), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_162), .B1(n_140), .B2(n_282), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_315), .A2(n_309), .B1(n_330), .B2(n_295), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_296), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_344), .A2(n_254), .B1(n_92), .B2(n_110), .C(n_210), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_333), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_301), .A2(n_162), .B1(n_140), .B2(n_293), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_301), .B(n_254), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_302), .A2(n_261), .B1(n_250), .B2(n_246), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_317), .A2(n_187), .B1(n_293), .B2(n_263), .Y(n_374) );
AO31x2_ASAP7_75t_L g375 ( .A1(n_321), .A2(n_127), .A3(n_145), .B(n_178), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_307), .B(n_140), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_297), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_369), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_321), .A3(n_322), .B(n_308), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_342), .B1(n_302), .B2(n_311), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_369), .B(n_304), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_369), .A2(n_302), .B(n_332), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_342), .B1(n_303), .B2(n_317), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_376), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_355), .A2(n_342), .B1(n_330), .B2(n_324), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_351), .A2(n_341), .B1(n_342), .B2(n_307), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_358), .B(n_329), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_349), .A2(n_331), .B1(n_318), .B2(n_322), .C(n_334), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_323), .B1(n_342), .B2(n_308), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_362), .A2(n_318), .B(n_324), .C(n_110), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_376), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_345), .B1(n_329), .B2(n_336), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_351), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_351), .A2(n_342), .B1(n_356), .B2(n_358), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_376), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_351), .A2(n_342), .B1(n_334), .B2(n_336), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_319), .B(n_337), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_345), .B1(n_343), .B2(n_337), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_347), .A2(n_313), .B1(n_343), .B2(n_306), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_366), .A2(n_324), .B1(n_327), .B2(n_313), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_347), .A2(n_313), .B1(n_332), .B2(n_324), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_361), .B(n_333), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_350), .B(n_327), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_401), .A2(n_360), .A3(n_378), .B1(n_354), .B2(n_350), .B3(n_127), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_402), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_357), .B1(n_365), .B2(n_354), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_397), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_390), .A2(n_378), .B1(n_366), .B2(n_327), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_393), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
OAI33xp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_145), .A3(n_178), .B1(n_363), .B2(n_377), .B3(n_374), .Y(n_418) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_367), .B(n_372), .Y(n_419) );
OAI33xp33_ASAP7_75t_L g420 ( .A1(n_403), .A2(n_373), .A3(n_185), .B1(n_210), .B2(n_225), .B3(n_14), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_327), .B1(n_92), .B2(n_110), .C(n_364), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_140), .B1(n_326), .B2(n_110), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_382), .B(n_92), .C(n_135), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_404), .A2(n_185), .A3(n_225), .B1(n_12), .B2(n_13), .B3(n_15), .Y(n_425) );
OAI31xp33_ASAP7_75t_SL g426 ( .A1(n_388), .A2(n_346), .A3(n_326), .B(n_12), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_383), .B(n_375), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_389), .B(n_375), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_381), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_391), .A2(n_140), .B1(n_92), .B2(n_313), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_389), .B(n_375), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_395), .B(n_375), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
OAI222xp33_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_368), .B1(n_370), .B2(n_313), .C1(n_371), .C2(n_17), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_381), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_396), .A2(n_339), .B1(n_370), .B2(n_368), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_399), .B(n_135), .C(n_147), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_411), .A2(n_426), .B(n_410), .C(n_422), .Y(n_441) );
OA332x1_ASAP7_75t_L g442 ( .A1(n_425), .A2(n_10), .A3(n_11), .B1(n_13), .B2(n_15), .B3(n_20), .C1(n_21), .C2(n_22), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_409), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_413), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_421), .B(n_395), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_412), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_379), .B1(n_400), .B2(n_405), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_407), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_424), .B(n_135), .C(n_147), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g453 ( .A(n_424), .B(n_379), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_421), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_440), .B(n_379), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_431), .B(n_375), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_420), .A2(n_384), .B1(n_149), .B2(n_147), .C(n_135), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_432), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_415), .B(n_370), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_414), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_435), .A2(n_149), .B(n_147), .C(n_135), .Y(n_462) );
OAI222xp33_ASAP7_75t_L g463 ( .A1(n_427), .A2(n_370), .B1(n_368), .B2(n_21), .C1(n_24), .C2(n_25), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_414), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_440), .A2(n_346), .B1(n_368), .B2(n_339), .Y(n_465) );
AOI33xp33_ASAP7_75t_L g466 ( .A1(n_429), .A2(n_201), .A3(n_188), .B1(n_24), .B2(n_26), .B3(n_11), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_431), .B(n_20), .Y(n_467) );
AOI21xp33_ASAP7_75t_SL g468 ( .A1(n_416), .A2(n_26), .B(n_36), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_427), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_432), .A2(n_314), .A3(n_312), .B(n_310), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_149), .Y(n_473) );
INVx11_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
AOI211xp5_ASAP7_75t_L g476 ( .A1(n_429), .A2(n_149), .B(n_147), .C(n_201), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_434), .A2(n_149), .B(n_147), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_434), .A2(n_149), .B1(n_147), .B2(n_188), .C(n_276), .Y(n_478) );
OAI33xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_149), .A3(n_325), .B1(n_291), .B2(n_286), .B3(n_276), .Y(n_479) );
OAI33xp33_ASAP7_75t_L g480 ( .A1(n_436), .A2(n_242), .A3(n_291), .B1(n_286), .B2(n_273), .B3(n_270), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_433), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_439), .B(n_298), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_433), .B(n_298), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_438), .B(n_298), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_408), .B(n_314), .C(n_312), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_419), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_430), .A2(n_314), .B(n_312), .C(n_310), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_419), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_444), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_445), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_444), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_467), .B(n_454), .Y(n_493) );
NOR2x1_ASAP7_75t_L g494 ( .A(n_453), .B(n_419), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_457), .B(n_430), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_457), .B(n_423), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_459), .B(n_39), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_459), .B(n_42), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_456), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_456), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_471), .B(n_43), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_467), .B(n_298), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_471), .B(n_44), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_484), .B(n_47), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_475), .B(n_48), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_484), .B(n_53), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_470), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_464), .B(n_310), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_314), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_487), .B(n_54), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_441), .A2(n_418), .B1(n_209), .B2(n_175), .C(n_270), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_452), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_487), .B(n_55), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_461), .B(n_312), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_486), .A2(n_310), .B1(n_333), .B2(n_177), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_463), .A2(n_340), .B(n_187), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_462), .A2(n_333), .B1(n_177), .B2(n_187), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_466), .B(n_209), .C(n_175), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_469), .B(n_57), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_446), .B(n_58), .Y(n_522) );
NAND2xp67_ASAP7_75t_L g523 ( .A(n_442), .B(n_59), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_475), .B(n_61), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_449), .A2(n_177), .B1(n_209), .B2(n_175), .C(n_256), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_443), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_443), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_468), .B(n_209), .C(n_175), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_468), .B(n_458), .C(n_480), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_450), .B(n_72), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_447), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_447), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_489), .B(n_73), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_481), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_450), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_465), .B(n_187), .Y(n_537) );
AND4x1_ASAP7_75t_L g538 ( .A(n_476), .B(n_177), .C(n_187), .D(n_175), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_489), .B(n_209), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_455), .B(n_242), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_473), .B(n_262), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_482), .B(n_262), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_483), .B(n_256), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_460), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_474), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_495), .B(n_472), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_495), .B(n_485), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_490), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_490), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_492), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_491), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_513), .B(n_442), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_492), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_493), .B(n_499), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_528), .A2(n_477), .B(n_488), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_499), .B(n_485), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_500), .B(n_478), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_500), .B(n_451), .Y(n_559) );
XOR2x2_ASAP7_75t_L g560 ( .A(n_497), .B(n_474), .Y(n_560) );
AND2x4_ASAP7_75t_SL g561 ( .A(n_497), .B(n_479), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_508), .B(n_273), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_508), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_546), .A2(n_246), .B1(n_250), .B2(n_261), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_523), .A2(n_246), .B(n_250), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_519), .B(n_246), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_519), .B(n_246), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_546), .A2(n_250), .B1(n_261), .B2(n_263), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_531), .B(n_261), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
NAND3xp33_ASAP7_75t_SL g573 ( .A(n_538), .B(n_261), .C(n_263), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_531), .B(n_264), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_546), .B(n_264), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_528), .B(n_264), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_536), .B(n_264), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_546), .B(n_264), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_535), .B(n_293), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_535), .B(n_293), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_498), .A2(n_293), .B1(n_541), .B2(n_501), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_533), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_496), .B(n_532), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_498), .B(n_530), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_545), .B(n_510), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_496), .B(n_539), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_501), .B(n_503), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_518), .A2(n_520), .B(n_503), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_506), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_545), .B(n_523), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_530), .B(n_538), .Y(n_594) );
INVx4_ASAP7_75t_L g595 ( .A(n_506), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_515), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_502), .B(n_534), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_576), .B(n_595), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_591), .A2(n_520), .B(n_518), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_552), .A2(n_494), .B(n_534), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_555), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_549), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_595), .B(n_494), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_553), .A2(n_529), .B(n_521), .C(n_537), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_554), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_586), .B(n_515), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_595), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_589), .B(n_548), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_563), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_550), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_560), .A2(n_506), .B1(n_512), .B2(n_522), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_560), .B(n_506), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_556), .B(n_524), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_568), .B(n_544), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_589), .B(n_539), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_551), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_594), .B(n_524), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_588), .B(n_544), .Y(n_621) );
AOI32xp33_ASAP7_75t_L g622 ( .A1(n_561), .A2(n_505), .A3(n_507), .B1(n_514), .B2(n_511), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_592), .B(n_505), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_578), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_588), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_593), .B(n_509), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_571), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g628 ( .A(n_548), .B(n_542), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_585), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_547), .A2(n_525), .B1(n_511), .B2(n_514), .C(n_507), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_596), .B(n_542), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
AOI21xp5_ASAP7_75t_SL g633 ( .A1(n_587), .A2(n_543), .B(n_540), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_596), .B(n_516), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_572), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_577), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_577), .Y(n_637) );
AOI221x1_ASAP7_75t_SL g638 ( .A1(n_565), .A2(n_517), .B1(n_590), .B2(n_597), .C(n_592), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_558), .B(n_547), .Y(n_639) );
XNOR2x1_ASAP7_75t_L g640 ( .A(n_582), .B(n_578), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_557), .B(n_558), .C(n_559), .D(n_575), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_579), .A2(n_561), .B(n_584), .Y(n_642) );
NAND2xp33_ASAP7_75t_L g643 ( .A(n_584), .B(n_583), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_562), .B(n_567), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_573), .A2(n_569), .B(n_564), .C(n_583), .Y(n_645) );
O2A1O1Ixp5_ASAP7_75t_L g646 ( .A1(n_562), .A2(n_566), .B(n_567), .C(n_580), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_562), .B(n_580), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_581), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_581), .A2(n_574), .B(n_570), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_574), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_570), .B(n_586), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_549), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_553), .A2(n_593), .B(n_309), .C(n_591), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_549), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_653), .A2(n_646), .B(n_600), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_602), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_615), .A2(n_639), .B1(n_616), .B2(n_640), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_616), .A2(n_640), .B1(n_626), .B2(n_641), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_620), .B(n_642), .C(n_606), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_610), .A2(n_628), .B1(n_644), .B2(n_649), .Y(n_660) );
AOI22x1_ASAP7_75t_L g661 ( .A1(n_610), .A2(n_624), .B1(n_638), .B2(n_615), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_626), .A2(n_646), .B1(n_625), .B2(n_611), .C(n_622), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_634), .A2(n_620), .B1(n_601), .B2(n_644), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_637), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_636), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_635), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g667 ( .A1(n_605), .A2(n_651), .B(n_611), .Y(n_667) );
NOR4xp75_ASAP7_75t_L g668 ( .A(n_605), .B(n_599), .C(n_610), .D(n_617), .Y(n_668) );
OAI211xp5_ASAP7_75t_L g669 ( .A1(n_661), .A2(n_614), .B(n_599), .C(n_630), .Y(n_669) );
OA211x2_ASAP7_75t_L g670 ( .A1(n_655), .A2(n_621), .B(n_631), .C(n_645), .Y(n_670) );
NOR3x1_ASAP7_75t_L g671 ( .A(n_660), .B(n_608), .C(n_647), .Y(n_671) );
AND3x2_ASAP7_75t_L g672 ( .A(n_659), .B(n_618), .C(n_623), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_662), .B(n_643), .C(n_629), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_658), .A2(n_643), .B1(n_648), .B2(n_619), .C(n_613), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_658), .A2(n_627), .B(n_632), .Y(n_675) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_657), .A2(n_650), .B(n_618), .C(n_604), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_673), .Y(n_677) );
XNOR2xp5_ASAP7_75t_L g678 ( .A(n_670), .B(n_656), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_674), .A2(n_663), .B1(n_667), .B2(n_623), .Y(n_679) );
NOR2x2_ASAP7_75t_L g680 ( .A(n_671), .B(n_668), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_669), .B(n_663), .C(n_665), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_676), .B1(n_675), .B2(n_672), .Y(n_682) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_678), .A2(n_666), .B1(n_664), .B2(n_623), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_677), .B(n_598), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_683), .A2(n_679), .B(n_680), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_682), .B(n_603), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_685), .B(n_684), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_686), .B(n_609), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_607), .B(n_652), .Y(n_689) );
AOI21xp33_ASAP7_75t_SL g690 ( .A1(n_689), .A2(n_612), .B(n_654), .Y(n_690) );
endmodule