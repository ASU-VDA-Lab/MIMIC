module fake_netlist_6_2133_n_762 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_762);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_762;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_724;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_372;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_139;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_68),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_136),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_62),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_39),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_82),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_95),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_50),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_41),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_119),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_109),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_32),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_84),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_98),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_81),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_101),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_63),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_112),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_79),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_30),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_51),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_46),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_26),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_154),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_0),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_1),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_143),
.B(n_2),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_135),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_22),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_132),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_23),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_2),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_3),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_24),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_3),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_142),
.B(n_25),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_4),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_4),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_5),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_146),
.B(n_5),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_147),
.B(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_190),
.B1(n_189),
.B2(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_167),
.B1(n_186),
.B2(n_184),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_155),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_166),
.B1(n_181),
.B2(n_179),
.Y(n_234)
);

OR2x6_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_6),
.Y(n_235)
);

AO22x2_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_165),
.B1(n_176),
.B2(n_171),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

AO22x2_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_R g240 ( 
.A1(n_209),
.A2(n_192),
.B1(n_217),
.B2(n_195),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_197),
.B1(n_213),
.B2(n_224),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_162),
.B1(n_170),
.B2(n_169),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_187),
.B1(n_168),
.B2(n_163),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_226),
.B1(n_191),
.B2(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_160),
.B1(n_157),
.B2(n_156),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_161),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g248 ( 
.A1(n_201),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_215),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_27),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_13),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_193),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g256 ( 
.A1(n_195),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_R g257 ( 
.A1(n_209),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_258)
);

AO22x2_ASAP7_75t_L g259 ( 
.A1(n_201),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_259)
);

AOI22x1_ASAP7_75t_SL g260 ( 
.A1(n_225),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_201),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_215),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_215),
.Y(n_266)
);

AOI22x1_ASAP7_75t_SL g267 ( 
.A1(n_221),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_202),
.A2(n_204),
.B1(n_214),
.B2(n_227),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_201),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_53),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_219),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_203),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_203),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

BUFx6f_ASAP7_75t_SL g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_202),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_220),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_236),
.B(n_203),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_202),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

NAND2x1p5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_203),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_273),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_206),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_204),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_204),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_220),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_206),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_206),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_259),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_235),
.B(n_214),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_243),
.B(n_206),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_234),
.B(n_220),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_237),
.A2(n_207),
.B(n_221),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_221),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_247),
.B(n_229),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_236),
.B(n_221),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_231),
.B(n_229),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_229),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_258),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_240),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_260),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_233),
.B(n_229),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_238),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_252),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_229),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_218),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_289),
.B(n_280),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_287),
.B(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_292),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_280),
.B(n_229),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_218),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_324),
.Y(n_360)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_304),
.B(n_207),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_317),
.B(n_207),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_326),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_207),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_207),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_207),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_207),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_279),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_295),
.B(n_208),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_318),
.Y(n_379)
);

BUFx4f_ASAP7_75t_SL g380 ( 
.A(n_326),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_302),
.B(n_61),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_293),
.B(n_218),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_295),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_303),
.B(n_208),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_283),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_293),
.B(n_211),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_302),
.B(n_211),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_278),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_313),
.B(n_64),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_318),
.B(n_211),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_294),
.B(n_66),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_211),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_294),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_300),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_322),
.B(n_211),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_315),
.A2(n_325),
.B(n_335),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_316),
.B(n_208),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_298),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_298),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

BUFx4f_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_305),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_305),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_327),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_397),
.B(n_306),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_307),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_343),
.B(n_312),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_319),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_320),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

NAND2x1_ASAP7_75t_L g428 ( 
.A(n_374),
.B(n_323),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_343),
.B(n_297),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_384),
.B(n_329),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_297),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_330),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_374),
.B(n_333),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_333),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_380),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_363),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_291),
.Y(n_442)
);

AND2x2_ASAP7_75t_SL g443 ( 
.A(n_399),
.B(n_334),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_350),
.B(n_331),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_353),
.B(n_334),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_368),
.B(n_291),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

NAND2x1_ASAP7_75t_L g454 ( 
.A(n_374),
.B(n_198),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_388),
.B(n_308),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_388),
.B(n_401),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_67),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_374),
.B(n_196),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_371),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_377),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_354),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_430),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_346),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_385),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_416),
.Y(n_473)
);

BUFx4f_ASAP7_75t_SL g474 ( 
.A(n_464),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_435),
.A2(n_404),
.B1(n_398),
.B2(n_399),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_445),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_410),
.A2(n_398),
.B1(n_367),
.B2(n_405),
.Y(n_484)
);

BUFx8_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_416),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_416),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_430),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_430),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_453),
.Y(n_496)
);

BUFx6f_ASAP7_75t_SL g497 ( 
.A(n_437),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_434),
.B(n_401),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_431),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_464),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_451),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_431),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_400),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_460),
.Y(n_509)
);

BUFx4_ASAP7_75t_SL g510 ( 
.A(n_441),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_395),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_474),
.A2(n_435),
.B1(n_414),
.B2(n_413),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_469),
.A2(n_410),
.B1(n_455),
.B2(n_458),
.Y(n_513)
);

BUFx2_ASAP7_75t_SL g514 ( 
.A(n_479),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_410),
.B1(n_442),
.B2(n_450),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_498),
.A2(n_444),
.B1(n_415),
.B2(n_447),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_503),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_498),
.A2(n_415),
.B1(n_459),
.B2(n_443),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_444),
.B1(n_447),
.B2(n_437),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_444),
.B1(n_443),
.B2(n_457),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_479),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_478),
.A2(n_451),
.B1(n_452),
.B2(n_439),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_472),
.A2(n_511),
.B1(n_505),
.B2(n_452),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_509),
.A2(n_422),
.B1(n_438),
.B2(n_427),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_501),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_424),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_475),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_509),
.A2(n_423),
.B1(n_421),
.B2(n_438),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_507),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_480),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_476),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_481),
.Y(n_543)
);

BUFx2_ASAP7_75t_SL g544 ( 
.A(n_488),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_487),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_485),
.A2(n_457),
.B1(n_285),
.B2(n_441),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_497),
.A2(n_427),
.B1(n_418),
.B2(n_460),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_485),
.A2(n_285),
.B1(n_438),
.B2(n_361),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_490),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_497),
.A2(n_285),
.B1(n_361),
.B2(n_440),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_512),
.A2(n_497),
.B1(n_460),
.B2(n_400),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_547),
.A2(n_477),
.B1(n_400),
.B2(n_361),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_515),
.A2(n_516),
.B1(n_520),
.B2(n_518),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_517),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_546),
.A2(n_550),
.B(n_552),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_522),
.Y(n_558)
);

BUFx8_ASAP7_75t_SL g559 ( 
.A(n_525),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_515),
.A2(n_400),
.B1(n_378),
.B2(n_373),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_518),
.A2(n_521),
.B1(n_513),
.B2(n_533),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_L g562 ( 
.A1(n_526),
.A2(n_418),
.B(n_471),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_519),
.B(n_486),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_539),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_524),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_547),
.A2(n_544),
.B1(n_514),
.B2(n_542),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_534),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_531),
.B(n_423),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_540),
.Y(n_569)
);

OAI22x1_ASAP7_75t_L g570 ( 
.A1(n_530),
.A2(n_421),
.B1(n_504),
.B2(n_407),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_549),
.A2(n_421),
.B1(n_378),
.B2(n_373),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_547),
.A2(n_391),
.B1(n_370),
.B2(n_484),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_530),
.A2(n_536),
.B1(n_535),
.B2(n_528),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_513),
.A2(n_378),
.B1(n_373),
.B2(n_389),
.Y(n_574)
);

BUFx4f_ASAP7_75t_SL g575 ( 
.A(n_538),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_526),
.A2(n_428),
.B1(n_491),
.B2(n_504),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_529),
.A2(n_389),
.B1(n_392),
.B2(n_387),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_536),
.A2(n_467),
.B1(n_376),
.B2(n_362),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_529),
.A2(n_392),
.B1(n_387),
.B2(n_372),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_527),
.A2(n_372),
.B1(n_409),
.B2(n_375),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_527),
.A2(n_428),
.B1(n_491),
.B2(n_495),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_523),
.A2(n_409),
.B1(n_375),
.B2(n_390),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_409),
.B1(n_375),
.B2(n_390),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_537),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_545),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_538),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_541),
.A2(n_394),
.B1(n_369),
.B2(n_357),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_541),
.A2(n_394),
.B1(n_369),
.B2(n_357),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_539),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_541),
.A2(n_491),
.B1(n_500),
.B2(n_371),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_548),
.A2(n_394),
.B1(n_362),
.B2(n_396),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_548),
.A2(n_467),
.B1(n_362),
.B2(n_365),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_548),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_512),
.A2(n_362),
.B1(n_396),
.B2(n_406),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_539),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_547),
.A2(n_365),
.B1(n_492),
.B2(n_473),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_568),
.B(n_483),
.Y(n_601)
);

NOR3xp33_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_408),
.C(n_407),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_579),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_403),
.B1(n_408),
.B2(n_395),
.C(n_205),
.Y(n_604)
);

OAI221xp5_ASAP7_75t_L g605 ( 
.A1(n_553),
.A2(n_342),
.B1(n_386),
.B2(n_402),
.C(n_364),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_555),
.A2(n_396),
.B1(n_365),
.B2(n_354),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_561),
.A2(n_396),
.B1(n_365),
.B2(n_354),
.Y(n_607)
);

HB1xp67_ASAP7_75t_SL g608 ( 
.A(n_558),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_402),
.B1(n_473),
.B2(n_492),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_573),
.A2(n_483),
.B1(n_489),
.B2(n_482),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_556),
.A2(n_473),
.B1(n_492),
.B2(n_499),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_598),
.A2(n_489),
.B1(n_482),
.B2(n_502),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_563),
.B(n_502),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_566),
.B(n_499),
.Y(n_614)
);

OAI221xp5_ASAP7_75t_L g615 ( 
.A1(n_557),
.A2(n_402),
.B1(n_358),
.B2(n_502),
.C(n_506),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_580),
.B(n_205),
.C(n_208),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_581),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_581),
.B(n_506),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_588),
.A2(n_402),
.B1(n_449),
.B2(n_462),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_588),
.A2(n_506),
.B1(n_456),
.B2(n_466),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_596),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_572),
.A2(n_466),
.B1(n_456),
.B2(n_470),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g623 ( 
.A1(n_556),
.A2(n_493),
.B1(n_470),
.B2(n_468),
.Y(n_623)
);

OAI222xp33_ASAP7_75t_L g624 ( 
.A1(n_577),
.A2(n_493),
.B1(n_470),
.B2(n_468),
.C1(n_429),
.C2(n_420),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_558),
.A2(n_383),
.B1(n_382),
.B2(n_371),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_205),
.B1(n_208),
.B2(n_426),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_589),
.B(n_205),
.C(n_208),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_587),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_567),
.B(n_468),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_560),
.A2(n_426),
.B1(n_420),
.B2(n_429),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_571),
.A2(n_493),
.B1(n_461),
.B2(n_351),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_570),
.A2(n_351),
.B1(n_463),
.B2(n_462),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_591),
.A2(n_463),
.B1(n_462),
.B2(n_449),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_578),
.A2(n_351),
.B1(n_463),
.B2(n_462),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_L g635 ( 
.A1(n_582),
.A2(n_351),
.B(n_510),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_69),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_567),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_569),
.Y(n_638)
);

AOI221xp5_ASAP7_75t_L g639 ( 
.A1(n_604),
.A2(n_576),
.B1(n_583),
.B2(n_569),
.C(n_574),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_621),
.B(n_597),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_617),
.B(n_590),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_602),
.B(n_600),
.C(n_584),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_613),
.B(n_575),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_610),
.B(n_602),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_608),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_637),
.B(n_585),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_615),
.B(n_594),
.C(n_595),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_614),
.B(n_592),
.C(n_599),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_624),
.A2(n_593),
.B(n_599),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_601),
.B(n_564),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_564),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_618),
.B(n_564),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_607),
.B(n_579),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_606),
.B(n_559),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_559),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_196),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_611),
.B(n_463),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_212),
.C(n_196),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_603),
.B(n_623),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_620),
.B(n_212),
.C(n_196),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_603),
.B(n_71),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_603),
.B(n_72),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_634),
.A2(n_73),
.B(n_75),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_632),
.B(n_212),
.C(n_462),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_651),
.B(n_622),
.Y(n_665)
);

NOR3xp33_ASAP7_75t_L g666 ( 
.A(n_644),
.B(n_605),
.C(n_616),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_649),
.B(n_609),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_644),
.A2(n_612),
.B1(n_627),
.B2(n_619),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_650),
.B(n_638),
.Y(n_669)
);

NAND4xp75_ASAP7_75t_L g670 ( 
.A(n_657),
.B(n_625),
.C(n_633),
.D(n_83),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_648),
.B(n_631),
.Y(n_671)
);

NAND4xp75_ASAP7_75t_L g672 ( 
.A(n_657),
.B(n_78),
.C(n_80),
.D(n_85),
.Y(n_672)
);

NAND4xp75_ASAP7_75t_L g673 ( 
.A(n_659),
.B(n_87),
.C(n_89),
.D(n_90),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_643),
.B(n_91),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_649),
.B(n_626),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_652),
.B(n_626),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_642),
.B(n_630),
.C(n_212),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_655),
.B(n_92),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_641),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_640),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_649),
.B(n_630),
.Y(n_681)
);

NOR4xp25_ASAP7_75t_L g682 ( 
.A(n_647),
.B(n_93),
.C(n_94),
.D(n_96),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_679),
.B(n_646),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_669),
.Y(n_684)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_680),
.B(n_645),
.Y(n_685)
);

NOR4xp25_ASAP7_75t_L g686 ( 
.A(n_671),
.B(n_663),
.C(n_654),
.D(n_658),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_676),
.B(n_639),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_676),
.B(n_656),
.Y(n_689)
);

NAND4xp75_ASAP7_75t_SL g690 ( 
.A(n_675),
.B(n_662),
.C(n_664),
.D(n_660),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_665),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_667),
.B(n_653),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_685),
.B(n_673),
.Y(n_694)
);

OA22x2_ASAP7_75t_L g695 ( 
.A1(n_691),
.A2(n_671),
.B1(n_681),
.B2(n_675),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_665),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_691),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_687),
.B1(n_693),
.B2(n_689),
.Y(n_699)
);

OAI22x1_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_684),
.B1(n_688),
.B2(n_692),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_697),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_698),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_694),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_703),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_701),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_702),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

OAI322xp33_ASAP7_75t_L g708 ( 
.A1(n_704),
.A2(n_699),
.A3(n_694),
.B1(n_683),
.B2(n_677),
.C1(n_700),
.C2(n_692),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_705),
.A2(n_668),
.B1(n_683),
.B2(n_666),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_705),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_710),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_SL g712 ( 
.A1(n_709),
.A2(n_706),
.B(n_707),
.C(n_674),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_710),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_713),
.B(n_704),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_711),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_712),
.A2(n_704),
.B1(n_706),
.B2(n_707),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_706),
.B1(n_704),
.B2(n_672),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_711),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_711),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_713),
.B(n_704),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_715),
.B(n_704),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_721),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_719),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_706),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_720),
.Y(n_726)
);

NOR2x1_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_690),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_718),
.B(n_661),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_716),
.B(n_99),
.Y(n_729)
);

AND4x1_ASAP7_75t_L g730 ( 
.A(n_727),
.B(n_686),
.C(n_682),
.D(n_681),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_723),
.A2(n_670),
.B1(n_463),
.B2(n_431),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_722),
.B(n_100),
.Y(n_732)
);

OR3x2_ASAP7_75t_L g733 ( 
.A(n_724),
.B(n_103),
.C(n_104),
.Y(n_733)
);

AND4x1_ASAP7_75t_L g734 ( 
.A(n_728),
.B(n_726),
.C(n_725),
.D(n_729),
.Y(n_734)
);

NOR4xp25_ASAP7_75t_L g735 ( 
.A(n_722),
.B(n_105),
.C(n_106),
.D(n_107),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_722),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_722),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_732),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_110),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_737),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_734),
.Y(n_741)
);

OAI211xp5_ASAP7_75t_L g742 ( 
.A1(n_735),
.A2(n_212),
.B(n_198),
.C(n_449),
.Y(n_742)
);

BUFx4f_ASAP7_75t_SL g743 ( 
.A(n_733),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_731),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_730),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_449),
.B1(n_212),
.B2(n_383),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_745),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_741),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_449),
.B1(n_383),
.B2(n_382),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_740),
.A2(n_383),
.B1(n_382),
.B2(n_371),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_738),
.A2(n_383),
.B1(n_382),
.B2(n_371),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_746),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_753),
.A2(n_744),
.B1(n_742),
.B2(n_751),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_SL g757 ( 
.A1(n_752),
.A2(n_739),
.B1(n_750),
.B2(n_382),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_757),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_L g759 ( 
.A1(n_758),
.A2(n_756),
.B1(n_755),
.B2(n_754),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_759),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_754),
.B1(n_454),
.B2(n_116),
.C(n_117),
.Y(n_761)
);

AOI211xp5_ASAP7_75t_L g762 ( 
.A1(n_761),
.A2(n_113),
.B(n_114),
.C(n_118),
.Y(n_762)
);


endmodule