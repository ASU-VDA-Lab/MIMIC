module fake_netlist_1_12327_n_500 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_500);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_500;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_84;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_5), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_24), .Y(n_71) );
INVxp67_ASAP7_75t_L g72 ( .A(n_27), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_38), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_61), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_28), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_16), .Y(n_76) );
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_18), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_35), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_55), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_62), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_69), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_66), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_4), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_26), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_5), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_25), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_56), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_39), .Y(n_98) );
AND2x2_ASAP7_75t_L g99 ( .A(n_23), .B(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_37), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_46), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_70), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_74), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_77), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_104), .B(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_79), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_79), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_93), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_80), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_93), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_96), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_96), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_86), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_87), .B(n_0), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_114), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_127), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_127), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_115), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_107), .B(n_98), .Y(n_132) );
BUFx10_ASAP7_75t_L g133 ( .A(n_117), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
BUFx4f_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx5_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_111), .B(n_76), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_106), .B(n_76), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
INVxp33_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_109), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_127), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_113), .B(n_71), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_113), .A2(n_103), .B1(n_94), .B2(n_100), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
CKINVDCx8_ASAP7_75t_R g150 ( .A(n_110), .Y(n_150) );
AND3x4_ASAP7_75t_L g151 ( .A(n_112), .B(n_86), .C(n_89), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_132), .B(n_121), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_134), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_131), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_136), .A2(n_126), .B(n_116), .C(n_118), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_142), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_134), .B(n_122), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_134), .B(n_116), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_139), .B(n_112), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_139), .B(n_138), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_136), .B(n_89), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_136), .Y(n_167) );
NOR2xp33_ASAP7_75t_R g168 ( .A(n_150), .B(n_126), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_146), .B(n_118), .Y(n_170) );
NOR3xp33_ASAP7_75t_SL g171 ( .A(n_145), .B(n_125), .C(n_97), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_131), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_146), .B(n_126), .Y(n_174) );
NOR3xp33_ASAP7_75t_SL g175 ( .A(n_145), .B(n_88), .C(n_103), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_138), .B(n_126), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_128), .B(n_72), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_136), .B(n_124), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_147), .B(n_99), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_161), .B(n_147), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_154), .B(n_149), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_180), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_176), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_180), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_182), .Y(n_189) );
BUFx2_ASAP7_75t_SL g190 ( .A(n_173), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_138), .B(n_148), .C(n_108), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_161), .B(n_147), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_174), .A2(n_147), .B(n_138), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_156), .Y(n_198) );
AOI222xp33_ASAP7_75t_L g199 ( .A1(n_161), .A2(n_141), .B1(n_82), .B2(n_108), .C1(n_123), .C2(n_124), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_182), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_135), .B(n_129), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_160), .B(n_150), .Y(n_202) );
NOR2xp67_ASAP7_75t_L g203 ( .A(n_156), .B(n_1), .Y(n_203) );
INVx6_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
BUFx4f_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_167), .Y(n_209) );
INVx3_ASAP7_75t_SL g210 ( .A(n_165), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_171), .B(n_123), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_206), .B(n_153), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_188), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_212), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_212), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_212), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_189), .A2(n_175), .B1(n_123), .B2(n_124), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_208), .Y(n_219) );
NAND2xp33_ASAP7_75t_SL g220 ( .A(n_189), .B(n_151), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_197), .B(n_164), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_197), .A2(n_151), .B1(n_152), .B2(n_167), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_200), .A2(n_151), .B1(n_179), .B2(n_177), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_200), .B(n_164), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_186), .B(n_172), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_188), .A2(n_172), .B1(n_181), .B2(n_157), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_186), .B(n_133), .Y(n_228) );
BUFx8_ASAP7_75t_SL g229 ( .A(n_198), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_205), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_205), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_185), .B(n_133), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_133), .B1(n_99), .B2(n_91), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_202), .B(n_91), .Y(n_237) );
OAI21xp33_ASAP7_75t_SL g238 ( .A1(n_237), .A2(n_199), .B(n_203), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_219), .A2(n_191), .B(n_201), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_211), .B(n_207), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_217), .A2(n_178), .B(n_162), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_223), .B(n_192), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_219), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_223), .B(n_185), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_233), .B(n_184), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_237), .A2(n_202), .B1(n_204), .B2(n_193), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
OAI21xp33_ASAP7_75t_SL g249 ( .A1(n_237), .A2(n_199), .B(n_202), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_216), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_237), .A2(n_204), .B1(n_196), .B2(n_209), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_236), .Y(n_252) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_222), .A2(n_190), .B1(n_210), .B2(n_195), .C(n_194), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_221), .B(n_158), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_133), .B1(n_90), .B2(n_92), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_234), .B(n_158), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_249), .A2(n_218), .B1(n_237), .B2(n_222), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_249), .Y(n_261) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_238), .A2(n_224), .B(n_235), .C(n_233), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_246), .Y(n_263) );
OAI21x1_ASAP7_75t_SL g264 ( .A1(n_247), .A2(n_218), .B(n_236), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_238), .B(n_237), .C(n_224), .Y(n_265) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_239), .A2(n_227), .B(n_85), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_239), .A2(n_73), .B(n_105), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_252), .B(n_221), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_247), .A2(n_234), .B1(n_214), .B2(n_228), .C(n_231), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_239), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_244), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
NAND4xp25_ASAP7_75t_L g275 ( .A(n_253), .B(n_214), .C(n_234), .D(n_95), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_254), .Y(n_276) );
INVxp67_ASAP7_75t_R g277 ( .A(n_251), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_256), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g279 ( .A1(n_251), .A2(n_232), .B1(n_230), .B2(n_221), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_272), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_274), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_261), .B(n_248), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_261), .B(n_248), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_278), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_270), .B(n_245), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_266), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_266), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_265), .B(n_253), .C(n_255), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_260), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_278), .Y(n_292) );
AOI211xp5_ASAP7_75t_L g293 ( .A1(n_275), .A2(n_241), .B(n_257), .C(n_230), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_264), .A2(n_258), .B(n_256), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_271), .B(n_258), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_271), .B(n_241), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_262), .A2(n_263), .B1(n_264), .B2(n_259), .C(n_267), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_273), .B(n_254), .Y(n_302) );
OR2x6_ASAP7_75t_L g303 ( .A(n_276), .B(n_258), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_269), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_269), .B(n_240), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_276), .B(n_254), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_259), .B(n_250), .Y(n_308) );
AOI211xp5_ASAP7_75t_SL g309 ( .A1(n_293), .A2(n_277), .B(n_229), .C(n_250), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_291), .B(n_299), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_300), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_291), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_300), .B(n_250), .Y(n_313) );
NAND2xp33_ASAP7_75t_R g314 ( .A(n_296), .B(n_277), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_283), .B(n_268), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_299), .B(n_279), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_300), .B(n_268), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
NOR3xp33_ASAP7_75t_SL g320 ( .A(n_290), .B(n_84), .C(n_101), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_302), .B(n_240), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_304), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_240), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_281), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_306), .B(n_240), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_287), .B(n_240), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_280), .B(n_254), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_297), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_295), .B(n_250), .Y(n_335) );
OAI33xp33_ASAP7_75t_L g336 ( .A1(n_290), .A2(n_102), .A3(n_243), .B1(n_3), .B2(n_4), .B3(n_6), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_280), .B(n_1), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_280), .B(n_243), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_295), .B(n_2), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_282), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_305), .B(n_216), .Y(n_343) );
NAND4xp25_ASAP7_75t_L g344 ( .A(n_301), .B(n_231), .C(n_226), .D(n_135), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_286), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_282), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_305), .B(n_6), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_295), .B(n_7), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_319), .B(n_305), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_345), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_344), .A2(n_301), .B1(n_293), .B2(n_305), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_320), .A2(n_336), .B(n_348), .C(n_337), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_322), .B(n_295), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_342), .B(n_289), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_340), .Y(n_360) );
NAND2x1_ASAP7_75t_L g361 ( .A(n_341), .B(n_289), .Y(n_361) );
OAI322xp33_ASAP7_75t_L g362 ( .A1(n_316), .A2(n_308), .A3(n_288), .B1(n_289), .B2(n_298), .C1(n_296), .C2(n_292), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_333), .B(n_298), .Y(n_363) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_341), .B(n_289), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g365 ( .A1(n_348), .A2(n_288), .B(n_296), .Y(n_365) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_350), .B(n_296), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_315), .A2(n_288), .B1(n_303), .B2(n_307), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_309), .B(n_303), .C(n_307), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_311), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_303), .B1(n_292), .B2(n_286), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_347), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_350), .A2(n_292), .B1(n_231), .B2(n_230), .C1(n_232), .C2(n_225), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_318), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_303), .Y(n_376) );
OAI321xp33_ASAP7_75t_L g377 ( .A1(n_331), .A2(n_303), .A3(n_232), .B1(n_230), .B2(n_215), .C(n_225), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_321), .A2(n_226), .B1(n_140), .B2(n_143), .C(n_129), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_332), .B(n_7), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_327), .B(n_294), .Y(n_382) );
OAI21xp33_ASAP7_75t_SL g383 ( .A1(n_315), .A2(n_294), .B(n_242), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_313), .B(n_294), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_335), .B(n_9), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_311), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_338), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_327), .A2(n_226), .B1(n_140), .B2(n_143), .C(n_130), .Y(n_388) );
AOI21xp33_ASAP7_75t_SL g389 ( .A1(n_314), .A2(n_9), .B(n_10), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_317), .B(n_12), .Y(n_390) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_335), .A2(n_226), .A3(n_13), .B1(n_14), .B2(n_15), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_325), .A2(n_232), .B1(n_230), .B2(n_226), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_325), .A2(n_232), .B1(n_230), .B2(n_217), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_317), .A2(n_130), .B(n_217), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_313), .A2(n_242), .B(n_215), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
OAI21xp33_ASAP7_75t_SL g398 ( .A1(n_349), .A2(n_242), .B(n_225), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_343), .A2(n_232), .B(n_230), .C(n_130), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_318), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
AOI21x1_ASAP7_75t_SL g402 ( .A1(n_390), .A2(n_343), .B(n_313), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_357), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_330), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_366), .A2(n_343), .B1(n_330), .B2(n_329), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_369), .B(n_363), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_354), .A2(n_329), .B1(n_326), .B2(n_232), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_387), .B(n_326), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_373), .B(n_12), .Y(n_415) );
NOR3x1_ASAP7_75t_L g416 ( .A(n_368), .B(n_13), .C(n_14), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_389), .B(n_215), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_356), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_355), .A2(n_15), .B1(n_16), .B2(n_137), .C(n_169), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_364), .A2(n_215), .B1(n_163), .B2(n_169), .Y(n_420) );
AOI32xp33_ASAP7_75t_L g421 ( .A1(n_381), .A2(n_17), .A3(n_19), .B1(n_21), .B2(n_22), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_353), .B(n_29), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
NAND2xp33_ASAP7_75t_SL g424 ( .A(n_361), .B(n_30), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_376), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_386), .B(n_31), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_400), .B(n_32), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_375), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_380), .B(n_34), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_351), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_382), .B(n_36), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_385), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_365), .B(n_40), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_362), .B(n_41), .Y(n_436) );
AOI32xp33_ASAP7_75t_L g437 ( .A1(n_367), .A2(n_43), .A3(n_44), .B1(n_45), .B2(n_47), .Y(n_437) );
AOI211xp5_ASAP7_75t_L g438 ( .A1(n_383), .A2(n_169), .B(n_163), .C(n_158), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_371), .B(n_48), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_384), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_415), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_441), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g446 ( .A(n_434), .B(n_392), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_403), .B(n_377), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
NAND4xp75_ASAP7_75t_L g449 ( .A(n_416), .B(n_398), .C(n_388), .D(n_396), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_418), .B(n_374), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_430), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_436), .A2(n_399), .B1(n_395), .B2(n_393), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_432), .B(n_391), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_411), .B(n_379), .Y(n_454) );
XOR2x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_377), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_440), .B(n_50), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_423), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_427), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_404), .Y(n_462) );
AOI21xp33_ASAP7_75t_SL g463 ( .A1(n_437), .A2(n_52), .B(n_54), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_419), .B(n_178), .C(n_166), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_408), .B(n_57), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_409), .B(n_137), .Y(n_466) );
NOR2xp33_ASAP7_75t_R g467 ( .A(n_446), .B(n_424), .Y(n_467) );
AOI322xp5_ASAP7_75t_L g468 ( .A1(n_444), .A2(n_406), .A3(n_412), .B1(n_422), .B2(n_439), .C1(n_435), .C2(n_414), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_444), .B(n_414), .Y(n_469) );
NOR2xp67_ASAP7_75t_L g470 ( .A(n_463), .B(n_409), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_445), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g472 ( .A(n_449), .B(n_431), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_448), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_450), .B(n_425), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_453), .A2(n_409), .B1(n_421), .B2(n_433), .C(n_405), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_447), .A2(n_438), .B(n_420), .C(n_433), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_455), .A2(n_429), .B1(n_428), .B2(n_402), .Y(n_477) );
NOR2xp33_ASAP7_75t_R g478 ( .A(n_443), .B(n_428), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_466), .A2(n_429), .B(n_137), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_460), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_442), .B(n_58), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_454), .A2(n_59), .B(n_60), .Y(n_482) );
OAI211xp5_ASAP7_75t_L g483 ( .A1(n_452), .A2(n_137), .B(n_166), .C(n_162), .Y(n_483) );
NAND5xp2_ASAP7_75t_L g484 ( .A(n_464), .B(n_63), .C(n_64), .D(n_68), .E(n_137), .Y(n_484) );
NAND4xp75_ASAP7_75t_L g485 ( .A(n_456), .B(n_465), .C(n_459), .D(n_461), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_457), .A2(n_163), .B1(n_169), .B2(n_464), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_462), .B(n_169), .C(n_458), .Y(n_487) );
OAI221xp5_ASAP7_75t_R g488 ( .A1(n_451), .A2(n_446), .B1(n_406), .B2(n_452), .C(n_444), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_467), .A2(n_472), .B1(n_488), .B2(n_478), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_480), .Y(n_490) );
NOR2x1p5_ASAP7_75t_L g491 ( .A(n_485), .B(n_474), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_475), .B(n_482), .C(n_483), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_490), .Y(n_493) );
NOR4xp25_ASAP7_75t_L g494 ( .A(n_489), .B(n_482), .C(n_469), .D(n_476), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_492), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g496 ( .A1(n_495), .A2(n_491), .B1(n_470), .B2(n_471), .C1(n_473), .C2(n_481), .Y(n_496) );
NOR4xp25_ASAP7_75t_SL g497 ( .A(n_494), .B(n_468), .C(n_477), .D(n_484), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_496), .Y(n_498) );
OAI221xp5_ASAP7_75t_R g499 ( .A1(n_498), .A2(n_497), .B1(n_493), .B2(n_487), .C(n_486), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_499), .A2(n_493), .B(n_479), .Y(n_500) );
endmodule