module fake_jpeg_5721_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_24),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_42),
.Y(n_69)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_62),
.B1(n_16),
.B2(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_26),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_12),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_20),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_52),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_28),
.B1(n_23),
.B2(n_26),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_21),
.B1(n_18),
.B2(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_63),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_16),
.B1(n_17),
.B2(n_22),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_21),
.B1(n_20),
.B2(n_13),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_52),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_46),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_64),
.B1(n_65),
.B2(n_58),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_86),
.B1(n_64),
.B2(n_68),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_81),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_51),
.B(n_63),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_63),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_48),
.B1(n_52),
.B2(n_51),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_92),
.B1(n_90),
.B2(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_68),
.B1(n_54),
.B2(n_56),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_98),
.B1(n_102),
.B2(n_83),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_108),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_110),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_80),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_113),
.B1(n_93),
.B2(n_88),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_68),
.B1(n_64),
.B2(n_55),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_117),
.B(n_88),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_30),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_67),
.Y(n_119)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_75),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_126),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_138),
.B1(n_141),
.B2(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_86),
.B1(n_70),
.B2(n_89),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_137),
.B1(n_117),
.B2(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_76),
.B1(n_87),
.B2(n_58),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_73),
.C(n_79),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.C(n_110),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_73),
.C(n_79),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_135),
.Y(n_170)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_61),
.B1(n_77),
.B2(n_65),
.Y(n_137)
);

AO21x2_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_87),
.B(n_71),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_61),
.B(n_30),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_116),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_104),
.B1(n_135),
.B2(n_72),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_111),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_154),
.B1(n_162),
.B2(n_168),
.Y(n_195)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_99),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_155),
.C(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_108),
.B1(n_103),
.B2(n_117),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_171),
.B1(n_141),
.B2(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_117),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_103),
.B1(n_100),
.B2(n_112),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_100),
.B(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_122),
.B(n_143),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_105),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_105),
.C(n_59),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_169),
.C(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_47),
.C(n_44),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_72),
.B1(n_58),
.B2(n_104),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_137),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_183),
.B(n_150),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_187),
.B1(n_30),
.B2(n_61),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_133),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_182),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_178),
.C(n_185),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_125),
.C(n_139),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_153),
.B1(n_152),
.B2(n_157),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_181),
.B1(n_190),
.B2(n_166),
.Y(n_207)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_131),
.B1(n_141),
.B2(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_125),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_120),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_141),
.B1(n_72),
.B2(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_189),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_141),
.B1(n_120),
.B2(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_148),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_127),
.C(n_123),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_142),
.C(n_24),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_163),
.B1(n_171),
.B2(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_209),
.B1(n_216),
.B2(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_154),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_208),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_217),
.B(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_165),
.B1(n_162),
.B2(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_212),
.B1(n_32),
.B2(n_29),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_123),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_142),
.B1(n_30),
.B2(n_33),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_213),
.C(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_24),
.C(n_32),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_215),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_191),
.B1(n_196),
.B2(n_180),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_222),
.B(n_27),
.Y(n_256)
);

AOI21x1_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_173),
.B(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_185),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_177),
.C(n_174),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_237),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_239),
.B1(n_199),
.B2(n_209),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_24),
.C(n_32),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_240),
.C(n_210),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_33),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_29),
.C(n_27),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_244),
.B1(n_255),
.B2(n_226),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_205),
.B1(n_217),
.B2(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_211),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_219),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_206),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_228),
.C(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_210),
.B1(n_27),
.B2(n_19),
.Y(n_255)
);

FAx1_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_225),
.CI(n_236),
.CON(n_257),
.SN(n_257)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_263),
.B1(n_267),
.B2(n_266),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_229),
.B1(n_256),
.B2(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_269),
.C(n_0),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_235),
.B1(n_240),
.B2(n_2),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_9),
.C(n_14),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_9),
.C(n_15),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_0),
.C(n_1),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_276),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_251),
.B1(n_1),
.B2(n_3),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_275),
.A2(n_280),
.B1(n_12),
.B2(n_11),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_13),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_3),
.C(n_4),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_275),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_277),
.B(n_279),
.C(n_10),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_10),
.B1(n_12),
.B2(n_5),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_4),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_10),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_295),
.B(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_284),
.B(n_283),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_298),
.B(n_294),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_287),
.B(n_5),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_299),
.B(n_5),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_4),
.B(n_5),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_6),
.B(n_7),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_7),
.Y(n_307)
);


endmodule