module fake_netlist_5_719_n_2471 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_382, n_554, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2471);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2471;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2339;
wire n_2320;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_602;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_2460;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_2431;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_518),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_552),
.Y(n_579)
);

BUFx5_ASAP7_75t_L g580 ( 
.A(n_0),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_571),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_279),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_235),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_11),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_519),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_20),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_381),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_542),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_357),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_20),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_533),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_167),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_560),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_282),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_271),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_446),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_26),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_413),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_82),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_559),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_219),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_115),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_28),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_108),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_76),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_191),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_466),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_528),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_200),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_243),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_9),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_360),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_12),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_189),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_246),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_298),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_561),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_114),
.Y(n_620)
);

INVxp33_ASAP7_75t_L g621 ( 
.A(n_548),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_489),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_97),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_302),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_25),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_546),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_47),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_225),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_141),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_350),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_328),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_325),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_221),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_212),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_511),
.Y(n_635)
);

CKINVDCx14_ASAP7_75t_R g636 ( 
.A(n_361),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_116),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_113),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_175),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_395),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_442),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_453),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_411),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_452),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_364),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_112),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_123),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_193),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_18),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_398),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_267),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_431),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_445),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_496),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_377),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_129),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_8),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_501),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_508),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_327),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_213),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_412),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_209),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_447),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_507),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_78),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_383),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_309),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_59),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_121),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_275),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_451),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_233),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_294),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_462),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_93),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_540),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_467),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_154),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_543),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_311),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_459),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_448),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_563),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_283),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_279),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_267),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_574),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_539),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_420),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_73),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_99),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_395),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_292),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_427),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_259),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_474),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_30),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_166),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_113),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_303),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_547),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_31),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_425),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_198),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_268),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_75),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_412),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_523),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_328),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_16),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_433),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_306),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_58),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_379),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_550),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_421),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_174),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_162),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_285),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_343),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_488),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_336),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_468),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_541),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_352),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_480),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_142),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_399),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_320),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_103),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_450),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_414),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_229),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_55),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_562),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_347),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_372),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_173),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_193),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_100),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_149),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_354),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_372),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_215),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_505),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_39),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_23),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_117),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_409),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_535),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_208),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_263),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_260),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_510),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_475),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_129),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_403),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_146),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_185),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_529),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_326),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_314),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_190),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_329),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_325),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_206),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_176),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_47),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_225),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_183),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_18),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_498),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_271),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_36),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_469),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_238),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_252),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_429),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_6),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_237),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_257),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_355),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_440),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_33),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_417),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_92),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_492),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_51),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_333),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_22),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_295),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_84),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_282),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_240),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_149),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_219),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_375),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_580),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_580),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_580),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_635),
.Y(n_803)
);

CKINVDCx14_ASAP7_75t_R g804 ( 
.A(n_636),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_580),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_605),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_580),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_580),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_580),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_580),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_642),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_621),
.B(n_1),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_623),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_623),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_613),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_630),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_768),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_768),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_722),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_768),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_614),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_623),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_768),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_600),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_600),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_639),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_581),
.B(n_1),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_660),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_611),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_642),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_611),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_747),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_693),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_693),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_778),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_778),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_773),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_592),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_604),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_747),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_612),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_616),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_710),
.B(n_2),
.Y(n_846)
);

INVxp33_ASAP7_75t_SL g847 ( 
.A(n_582),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_640),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_661),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_615),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_624),
.Y(n_851)
);

INVxp33_ASAP7_75t_SL g852 ( 
.A(n_582),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_639),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_629),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_780),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_632),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_649),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_637),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_617),
.Y(n_859)
);

INVxp33_ASAP7_75t_L g860 ( 
.A(n_650),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_651),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_780),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_670),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_652),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_657),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_667),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_674),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_675),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_677),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_680),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_663),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_682),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_695),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_583),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_700),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_583),
.Y(n_876)
);

INVxp33_ASAP7_75t_L g877 ( 
.A(n_704),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_725),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_723),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_620),
.Y(n_880)
);

INVxp33_ASAP7_75t_SL g881 ( 
.A(n_584),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_707),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_723),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_719),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_720),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_625),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_724),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_729),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_701),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_734),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_627),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_741),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_663),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_668),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_628),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_754),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_584),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_761),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_763),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_725),
.B(n_2),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_874),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_830),
.A2(n_766),
.B1(n_589),
.B2(n_586),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_818),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_812),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_812),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_818),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_811),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_819),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_803),
.B(n_789),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_811),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_823),
.B(n_591),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_800),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_804),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_812),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_812),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_832),
.B(n_593),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_819),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_821),
.Y(n_920)
);

OAI22x1_ASAP7_75t_R g921 ( 
.A1(n_806),
.A2(n_794),
.B1(n_716),
.B2(n_586),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_820),
.A2(n_587),
.B1(n_594),
.B2(n_590),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_821),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_816),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_879),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_879),
.Y(n_928)
);

BUFx8_ASAP7_75t_SL g929 ( 
.A(n_806),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_824),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_816),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_834),
.B(n_697),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_800),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_813),
.B(n_665),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_801),
.A2(n_619),
.B(n_596),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_883),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_825),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_817),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_883),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_883),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_883),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_839),
.A2(n_587),
.B1(n_594),
.B2(n_590),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_843),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_843),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_823),
.B(n_654),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_825),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_802),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_805),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_853),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_829),
.A2(n_788),
.B1(n_790),
.B2(n_786),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_814),
.B(n_673),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_853),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_807),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_878),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_855),
.B(n_697),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_878),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_815),
.B(n_678),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_871),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_808),
.B(n_683),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_862),
.B(n_706),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_862),
.B(n_706),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_871),
.Y(n_962)
);

OAI22x1_ASAP7_75t_R g963 ( 
.A1(n_817),
.A2(n_598),
.B1(n_599),
.B2(n_595),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_831),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_905),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_905),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_929),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_909),
.B(n_894),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_938),
.B(n_822),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_915),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_915),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_905),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_964),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_R g974 ( 
.A(n_934),
.B(n_822),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_960),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_912),
.B(n_850),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_947),
.A2(n_810),
.B(n_809),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_964),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_925),
.B(n_679),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_911),
.B(n_850),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_909),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_931),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_909),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_912),
.B(n_859),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_914),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_943),
.B(n_859),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_944),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_944),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_921),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_944),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_922),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_943),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_921),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_959),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_948),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_905),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_960),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_905),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_963),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_963),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_948),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_933),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_953),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_R g1005 ( 
.A(n_932),
.B(n_880),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_961),
.B(n_880),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_942),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_953),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_953),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_902),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_904),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_918),
.Y(n_1012)
);

AND3x2_ASAP7_75t_L g1013 ( 
.A(n_961),
.B(n_901),
.C(n_840),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_950),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_904),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_950),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_933),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_903),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_932),
.B(n_886),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_955),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_951),
.B(n_957),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_933),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_955),
.B(n_886),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_919),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_908),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_908),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_951),
.B(n_891),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_959),
.B(n_891),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_R g1029 ( 
.A(n_935),
.B(n_895),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_935),
.A2(n_878),
.B(n_713),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_959),
.B(n_847),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_910),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_951),
.B(n_848),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_959),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_939),
.B(n_895),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_910),
.A2(n_728),
.B(n_696),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_919),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_935),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_L g1039 ( 
.A(n_949),
.B(n_723),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_920),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_939),
.B(n_849),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_951),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_923),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_957),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_935),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_957),
.A2(n_847),
.B1(n_881),
.B2(n_852),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_924),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_968),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_977),
.Y(n_1049)
);

NOR2x1p5_ASAP7_75t_L g1050 ( 
.A(n_1033),
.B(n_595),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_965),
.Y(n_1051)
);

XOR2xp5_ASAP7_75t_L g1052 ( 
.A(n_967),
.B(n_849),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_977),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_995),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_977),
.Y(n_1055)
);

AND2x6_ASAP7_75t_L g1056 ( 
.A(n_995),
.B(n_723),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_968),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_983),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_975),
.B(n_726),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_967),
.B(n_863),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1019),
.B(n_852),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_1021),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_985),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_976),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1021),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_1021),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1003),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_981),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_973),
.B(n_913),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1003),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_978),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_987),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1017),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1042),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_990),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_984),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1017),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1011),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1015),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1022),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_990),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1034),
.B(n_726),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1034),
.B(n_726),
.Y(n_1084)
);

INVx8_ASAP7_75t_L g1085 ( 
.A(n_970),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1038),
.A2(n_739),
.B1(n_740),
.B2(n_727),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_965),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1022),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_969),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_998),
.B(n_913),
.Y(n_1090)
);

AND3x1_ASAP7_75t_L g1091 ( 
.A(n_979),
.B(n_1046),
.C(n_1023),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1031),
.B(n_726),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1024),
.Y(n_1093)
);

INVxp33_ASAP7_75t_SL g1094 ( 
.A(n_974),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1006),
.B(n_881),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_988),
.B(n_913),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1024),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_965),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_971),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1025),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1026),
.B(n_913),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_L g1102 ( 
.A(n_1038),
.B(n_578),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1028),
.B(n_726),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_1027),
.B(n_752),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1032),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1040),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1037),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1043),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1037),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1005),
.B(n_846),
.C(n_898),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_992),
.B(n_945),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1047),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1047),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1020),
.B(n_876),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1041),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_994),
.A2(n_930),
.B(n_923),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_996),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1002),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1045),
.A2(n_739),
.B1(n_740),
.B2(n_727),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_SL g1121 ( 
.A(n_971),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1045),
.B(n_945),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1013),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1008),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_980),
.B(n_876),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1029),
.A2(n_945),
.B1(n_618),
.B2(n_622),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1044),
.A2(n_1020),
.B1(n_986),
.B2(n_1016),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

AND3x2_ASAP7_75t_L g1129 ( 
.A(n_993),
.B(n_857),
.C(n_781),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1009),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_966),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1044),
.B(n_945),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_970),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1030),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1036),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1010),
.B(n_757),
.Y(n_1136)
);

AND3x2_ASAP7_75t_L g1137 ( 
.A(n_971),
.B(n_781),
.C(n_770),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1036),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_982),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_966),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1036),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_966),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1035),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1030),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_982),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_966),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_972),
.B(n_937),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_972),
.B(n_937),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_972),
.B(n_946),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_972),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1007),
.B(n_646),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1014),
.B(n_1016),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1007),
.B(n_658),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_997),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1039),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_997),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_991),
.B(n_777),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_997),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1014),
.B(n_702),
.Y(n_1159)
);

INVxp33_ASAP7_75t_L g1160 ( 
.A(n_1018),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1039),
.Y(n_1161)
);

AOI22x1_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_833),
.B1(n_836),
.B2(n_835),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_999),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_999),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_999),
.B(n_787),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1018),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_999),
.Y(n_1167)
);

CKINVDCx6p67_ASAP7_75t_R g1168 ( 
.A(n_989),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_989),
.B(n_579),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1000),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1000),
.B(n_841),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1001),
.B(n_626),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1001),
.A2(n_749),
.B1(n_860),
.B2(n_858),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1012),
.B(n_877),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1174),
.B(n_863),
.Y(n_1175)
);

BUFx5_ASAP7_75t_L g1176 ( 
.A(n_1144),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1085),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1062),
.B(n_927),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1086),
.B(n_930),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1048),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1057),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1086),
.B(n_1120),
.Y(n_1182)
);

AO221x1_ASAP7_75t_L g1183 ( 
.A1(n_1127),
.A2(n_784),
.B1(n_791),
.B2(n_782),
.C(n_764),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1057),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1120),
.B(n_946),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1076),
.B(n_585),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1122),
.B(n_588),
.C(n_585),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1062),
.Y(n_1188)
);

INVxp33_ASAP7_75t_L g1189 ( 
.A(n_1114),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1062),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1095),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1095),
.B(n_889),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1094),
.B(n_588),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1049),
.B(n_924),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1107),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1151),
.B(n_597),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_SL g1197 ( 
.A(n_1076),
.B(n_1082),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_1085),
.B(n_837),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1079),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1060),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1080),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1066),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_L g1203 ( 
.A(n_1151),
.B(n_838),
.C(n_842),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1107),
.Y(n_1204)
);

AND2x2_ASAP7_75t_SL g1205 ( 
.A(n_1091),
.B(n_793),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1153),
.B(n_1065),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1153),
.B(n_1159),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1100),
.B(n_949),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1109),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1105),
.B(n_949),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1077),
.B(n_597),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1159),
.B(n_1061),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1106),
.B(n_958),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1112),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1066),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1118),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1049),
.B(n_958),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1059),
.B(n_608),
.C(n_601),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1061),
.B(n_601),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1060),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1090),
.B(n_1111),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1118),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1085),
.B(n_1099),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1115),
.B(n_608),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1066),
.B(n_1067),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1066),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1067),
.B(n_609),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1067),
.B(n_927),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1125),
.B(n_649),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1067),
.B(n_609),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1119),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1054),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1059),
.B(n_958),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1054),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1125),
.B(n_649),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1054),
.B(n_785),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1072),
.B(n_789),
.C(n_785),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1054),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1132),
.B(n_958),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1063),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1143),
.B(n_631),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1101),
.B(n_962),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1069),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1096),
.B(n_962),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1096),
.B(n_962),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1063),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1119),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1058),
.B(n_641),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1058),
.B(n_633),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1064),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1130),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_L g1253 ( 
.A(n_1173),
.B(n_845),
.C(n_844),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1087),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1073),
.B(n_643),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1133),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_L g1258 ( 
.A(n_1173),
.B(n_854),
.C(n_851),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1073),
.B(n_645),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1117),
.B(n_952),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1124),
.B(n_952),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1075),
.Y(n_1262)
);

NOR2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1099),
.B(n_598),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1097),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1126),
.B(n_653),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1110),
.B(n_655),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1136),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1157),
.B(n_634),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1139),
.B(n_1123),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1053),
.B(n_659),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1157),
.B(n_1069),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1139),
.B(n_1051),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_SL g1273 ( 
.A(n_1051),
.B(n_796),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1089),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1050),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1152),
.B(n_638),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1166),
.B(n_1136),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1171),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1093),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1087),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1102),
.A2(n_676),
.B1(n_681),
.B2(n_666),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1160),
.B(n_644),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1053),
.B(n_684),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1113),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1160),
.B(n_686),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1068),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1051),
.B(n_685),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1169),
.B(n_647),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1055),
.B(n_689),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1051),
.B(n_690),
.Y(n_1290)
);

INVxp33_ASAP7_75t_L g1291 ( 
.A(n_1052),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1055),
.B(n_939),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_1171),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1071),
.Y(n_1294)
);

NOR2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1168),
.B(n_599),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1113),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1074),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1135),
.A2(n_1141),
.B(n_1138),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1169),
.B(n_648),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1121),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1074),
.B(n_939),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1078),
.B(n_940),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1172),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1078),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1081),
.B(n_940),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1081),
.B(n_940),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1083),
.B(n_656),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1088),
.B(n_940),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1088),
.B(n_927),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1083),
.B(n_662),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1104),
.B(n_691),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1084),
.B(n_664),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1116),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1104),
.B(n_698),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1147),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1129),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1104),
.B(n_703),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1154),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1154),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1121),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_SL g1321 ( 
.A(n_1104),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1084),
.B(n_856),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1148),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1158),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1158),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

INVx8_ASAP7_75t_L g1327 ( 
.A(n_1104),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1134),
.A2(n_1103),
.B(n_1092),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1170),
.B(n_1092),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1087),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1103),
.B(n_705),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1167),
.B(n_669),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1087),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1155),
.B(n_671),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1070),
.B(n_686),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1161),
.B(n_672),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1070),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1128),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1131),
.B(n_717),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1128),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1129),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1131),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1131),
.B(n_718),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1131),
.B(n_733),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1146),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1140),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1165),
.B(n_756),
.C(n_737),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1140),
.B(n_762),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1146),
.Y(n_1349)
);

AO22x2_ASAP7_75t_L g1350 ( 
.A1(n_1182),
.A2(n_798),
.B1(n_797),
.B2(n_1165),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1207),
.B(n_1142),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1212),
.B(n_1056),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1199),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1222),
.B(n_1056),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1200),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1201),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1337),
.B(n_1137),
.Y(n_1357)
);

OAI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1268),
.A2(n_606),
.B1(n_607),
.B2(n_603),
.C(n_602),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1188),
.B(n_1098),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1244),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1214),
.Y(n_1361)
);

AO22x2_ASAP7_75t_L g1362 ( 
.A1(n_1182),
.A2(n_1137),
.B1(n_864),
.B2(n_865),
.Y(n_1362)
);

AO22x2_ASAP7_75t_L g1363 ( 
.A1(n_1230),
.A2(n_866),
.B1(n_867),
.B2(n_861),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1217),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1191),
.B(n_1140),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1223),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1232),
.Y(n_1367)
);

AO22x2_ASAP7_75t_L g1368 ( 
.A1(n_1236),
.A2(n_869),
.B1(n_870),
.B2(n_868),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1248),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1252),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1192),
.B(n_872),
.Y(n_1371)
);

AO22x2_ASAP7_75t_L g1372 ( 
.A1(n_1267),
.A2(n_875),
.B1(n_882),
.B2(n_873),
.Y(n_1372)
);

AO22x2_ASAP7_75t_L g1373 ( 
.A1(n_1219),
.A2(n_885),
.B1(n_887),
.B2(n_884),
.Y(n_1373)
);

AO22x2_ASAP7_75t_L g1374 ( 
.A1(n_1219),
.A2(n_890),
.B1(n_892),
.B2(n_888),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1241),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1247),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1175),
.B(n_897),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1180),
.Y(n_1378)
);

OAI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1196),
.A2(n_606),
.B1(n_607),
.B2(n_603),
.C(n_602),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1220),
.A2(n_786),
.B1(n_788),
.B2(n_783),
.C(n_610),
.Y(n_1380)
);

AO22x2_ASAP7_75t_L g1381 ( 
.A1(n_1206),
.A2(n_900),
.B1(n_899),
.B2(n_735),
.Y(n_1381)
);

AO22x2_ASAP7_75t_L g1382 ( 
.A1(n_1277),
.A2(n_735),
.B1(n_686),
.B2(n_826),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1215),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1271),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1304),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1276),
.B(n_735),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1255),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1262),
.B(n_1150),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1303),
.A2(n_1056),
.B1(n_774),
.B2(n_1150),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1187),
.A2(n_827),
.B1(n_828),
.B2(n_826),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1195),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1204),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1177),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1251),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1285),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1329),
.A2(n_1164),
.B1(n_1156),
.B2(n_1163),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1288),
.A2(n_790),
.B1(n_792),
.B2(n_783),
.C(n_610),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1188),
.B(n_1156),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1188),
.B(n_1163),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1299),
.A2(n_1056),
.B1(n_1164),
.B2(n_1140),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1316),
.Y(n_1401)
);

BUFx8_ASAP7_75t_L g1402 ( 
.A(n_1341),
.Y(n_1402)
);

NAND2x1p5_ASAP7_75t_L g1403 ( 
.A(n_1190),
.B(n_1162),
.Y(n_1403)
);

AO22x2_ASAP7_75t_L g1404 ( 
.A1(n_1187),
.A2(n_828),
.B1(n_893),
.B2(n_827),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1209),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1315),
.B(n_1056),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1323),
.B(n_687),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1326),
.B(n_688),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1189),
.B(n_692),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1278),
.A2(n_799),
.B1(n_795),
.B2(n_792),
.C(n_708),
.Y(n_1410)
);

AND2x6_ASAP7_75t_L g1411 ( 
.A(n_1190),
.B(n_893),
.Y(n_1411)
);

OAI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1293),
.A2(n_799),
.B1(n_795),
.B2(n_709),
.C(n_711),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1257),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1286),
.Y(n_1414)
);

AO22x2_ASAP7_75t_L g1415 ( 
.A1(n_1266),
.A2(n_896),
.B1(n_4),
.B2(n_0),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1282),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1225),
.B(n_694),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

AO22x2_ASAP7_75t_L g1419 ( 
.A1(n_1183),
.A2(n_896),
.B1(n_5),
.B2(n_3),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1202),
.B(n_954),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1334),
.B(n_699),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1336),
.B(n_712),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1224),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1297),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1193),
.B(n_714),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1260),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1205),
.B(n_715),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1181),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1261),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1233),
.Y(n_1430)
);

AO22x2_ASAP7_75t_L g1431 ( 
.A1(n_1253),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1274),
.Y(n_1432)
);

AO22x2_ASAP7_75t_L g1433 ( 
.A1(n_1258),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1264),
.Y(n_1434)
);

AO22x2_ASAP7_75t_L g1435 ( 
.A1(n_1272),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1279),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1284),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1203),
.A2(n_731),
.B1(n_732),
.B2(n_730),
.C(n_721),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1242),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1296),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1184),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1238),
.A2(n_1335),
.B1(n_1185),
.B2(n_1179),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1318),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1319),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1238),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1324),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1325),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1208),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1307),
.A2(n_738),
.B1(n_742),
.B2(n_736),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1210),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1345),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1310),
.A2(n_745),
.B1(n_746),
.B2(n_744),
.C(n_743),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_L g1453 ( 
.A(n_1250),
.B(n_415),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1313),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1213),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1301),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1312),
.B(n_894),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1179),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1302),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1302),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1224),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1269),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1197),
.B(n_954),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1305),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1269),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_L g1466 ( 
.A(n_1202),
.B(n_748),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1216),
.B(n_954),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1224),
.B(n_906),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1216),
.B(n_954),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1269),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1305),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1275),
.B(n_416),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1332),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1198),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1308),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1211),
.A2(n_753),
.B1(n_755),
.B2(n_751),
.C(n_750),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_SL g1478 ( 
.A(n_1198),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1197),
.B(n_954),
.Y(n_1479)
);

AO22x2_ASAP7_75t_L g1480 ( 
.A1(n_1185),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1292),
.Y(n_1481)
);

BUFx8_ASAP7_75t_L g1482 ( 
.A(n_1321),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1292),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1245),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1198),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1233),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1246),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1216),
.B(n_954),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1227),
.B(n_418),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1338),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1340),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1221),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1349),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1228),
.A2(n_760),
.B1(n_765),
.B2(n_759),
.C(n_758),
.Y(n_1494)
);

BUFx8_ASAP7_75t_L g1495 ( 
.A(n_1321),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1265),
.A2(n_771),
.B1(n_772),
.B2(n_769),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1339),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1239),
.B(n_775),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1227),
.B(n_906),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_L g1500 ( 
.A(n_1227),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1320),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1320),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1235),
.Y(n_1503)
);

OR2x6_ASAP7_75t_SL g1504 ( 
.A(n_1300),
.B(n_776),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1194),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1235),
.B(n_956),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1226),
.B(n_419),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1231),
.A2(n_779),
.B1(n_19),
.B2(n_16),
.C(n_17),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1254),
.B(n_956),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1218),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1218),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1240),
.B(n_19),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1298),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1237),
.A2(n_956),
.B1(n_907),
.B2(n_916),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1186),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1309),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1254),
.B(n_1346),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1254),
.Y(n_1518)
);

AO22x2_ASAP7_75t_L g1519 ( 
.A1(n_1347),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1291),
.B(n_27),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1263),
.B(n_906),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1249),
.B(n_27),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1351),
.A2(n_1243),
.B(n_1327),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1417),
.A2(n_1322),
.B1(n_1281),
.B2(n_1256),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1489),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1353),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1478),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1516),
.A2(n_1327),
.B(n_1314),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1471),
.A2(n_1328),
.B(n_1234),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1384),
.B(n_1339),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1354),
.A2(n_1479),
.B(n_1463),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1505),
.A2(n_1314),
.B(n_1311),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1356),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1371),
.B(n_1343),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1497),
.B(n_1343),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1426),
.B(n_1270),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1425),
.A2(n_1347),
.B1(n_1348),
.B2(n_1344),
.Y(n_1538)
);

OAI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1352),
.A2(n_1289),
.B(n_1283),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_L g1540 ( 
.A(n_1439),
.B(n_1259),
.C(n_1317),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1361),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1454),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1378),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1386),
.B(n_1295),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1522),
.A2(n_1331),
.B1(n_1287),
.B2(n_1290),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1429),
.B(n_1331),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1383),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1385),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1364),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1510),
.A2(n_1229),
.B(n_1178),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1430),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1377),
.B(n_1328),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1474),
.B(n_1416),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1387),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1511),
.A2(n_1229),
.B(n_1178),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1360),
.B(n_1342),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1396),
.A2(n_1342),
.B(n_1333),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1457),
.B(n_1280),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1481),
.A2(n_1346),
.B(n_1342),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1407),
.B(n_1280),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1408),
.B(n_1330),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1483),
.A2(n_1453),
.B(n_1406),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1442),
.A2(n_1450),
.B(n_1448),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1400),
.A2(n_1346),
.B1(n_1330),
.B2(n_1176),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1455),
.A2(n_1176),
.B(n_941),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_R g1568 ( 
.A(n_1502),
.B(n_1273),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1423),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1484),
.B(n_28),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1413),
.B(n_29),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1395),
.B(n_1427),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1366),
.A2(n_1369),
.B1(n_1370),
.B2(n_1367),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1512),
.A2(n_941),
.B(n_423),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1489),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1375),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1432),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1397),
.A2(n_32),
.B(n_29),
.C(n_30),
.Y(n_1578)
);

OAI321xp33_ASAP7_75t_L g1579 ( 
.A1(n_1515),
.A2(n_34),
.A3(n_36),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_1579)
);

AO22x1_ASAP7_75t_L g1580 ( 
.A1(n_1402),
.A2(n_1473),
.B1(n_1401),
.B2(n_1357),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1487),
.B(n_34),
.Y(n_1581)
);

BUFx4f_ASAP7_75t_L g1582 ( 
.A(n_1423),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1380),
.A2(n_907),
.B(n_916),
.C(n_906),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1363),
.B(n_35),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1363),
.B(n_37),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1368),
.B(n_37),
.Y(n_1586)
);

O2A1O1Ixp5_ASAP7_75t_L g1587 ( 
.A1(n_1365),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1358),
.A2(n_41),
.B(n_38),
.C(n_40),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1503),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1368),
.B(n_41),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1409),
.B(n_1492),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1456),
.B(n_42),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1379),
.B(n_42),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1376),
.Y(n_1594)
);

BUFx8_ASAP7_75t_L g1595 ( 
.A(n_1475),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_L g1596 ( 
.A(n_1498),
.B(n_422),
.Y(n_1596)
);

BUFx4f_ASAP7_75t_L g1597 ( 
.A(n_1475),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1459),
.B(n_43),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1393),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1460),
.A2(n_1472),
.B(n_1464),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1394),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1476),
.A2(n_917),
.B(n_916),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1414),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1452),
.B(n_43),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1513),
.A2(n_928),
.B(n_926),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1389),
.A2(n_426),
.B(n_424),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1424),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1402),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1388),
.B(n_926),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1470),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1441),
.A2(n_430),
.B(n_428),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1508),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1434),
.B(n_1388),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1372),
.B(n_44),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1372),
.B(n_45),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1507),
.B(n_46),
.Y(n_1616)
);

INVx11_ASAP7_75t_L g1617 ( 
.A(n_1482),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1436),
.A2(n_1437),
.B1(n_1440),
.B2(n_1428),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1391),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1392),
.A2(n_434),
.B(n_432),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1438),
.B(n_48),
.C(n_49),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1507),
.B(n_1373),
.Y(n_1622)
);

BUFx4f_ASAP7_75t_L g1623 ( 
.A(n_1357),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1415),
.A2(n_936),
.B1(n_50),
.B2(n_48),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1412),
.B(n_49),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1405),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1461),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1499),
.A2(n_936),
.B(n_436),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1499),
.A2(n_1398),
.B(n_1359),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1373),
.B(n_50),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1418),
.A2(n_437),
.B(n_435),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1443),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1449),
.B(n_936),
.C(n_52),
.Y(n_1633)
);

AOI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1350),
.A2(n_1404),
.B(n_1390),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1494),
.A2(n_1477),
.B(n_1410),
.C(n_1520),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1485),
.Y(n_1636)
);

BUFx4f_ASAP7_75t_L g1637 ( 
.A(n_1411),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1399),
.A2(n_439),
.B(n_438),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1415),
.A2(n_1431),
.B1(n_1433),
.B2(n_1374),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1374),
.B(n_53),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1444),
.A2(n_443),
.B(n_441),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1446),
.A2(n_449),
.B(n_444),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1473),
.B(n_54),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1451),
.B(n_54),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1466),
.A2(n_1496),
.B(n_1521),
.C(n_1490),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1447),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1355),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1390),
.B(n_55),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1468),
.A2(n_455),
.B(n_454),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1486),
.B(n_456),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1517),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1431),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1404),
.B(n_1381),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1509),
.A2(n_458),
.B(n_457),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1381),
.B(n_56),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1491),
.A2(n_461),
.B(n_460),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1411),
.B(n_57),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1518),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1521),
.B(n_577),
.Y(n_1659)
);

NAND2xp33_ASAP7_75t_L g1660 ( 
.A(n_1411),
.B(n_463),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1403),
.A2(n_1493),
.B(n_1514),
.Y(n_1661)
);

BUFx8_ASAP7_75t_L g1662 ( 
.A(n_1501),
.Y(n_1662)
);

NOR2xp67_ASAP7_75t_L g1663 ( 
.A(n_1482),
.B(n_576),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1420),
.A2(n_465),
.B(n_464),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1362),
.B(n_59),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1419),
.A2(n_575),
.B(n_471),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1495),
.B(n_470),
.Y(n_1667)
);

BUFx8_ASAP7_75t_L g1668 ( 
.A(n_1495),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1506),
.A2(n_1469),
.B(n_1467),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1382),
.B(n_60),
.Y(n_1670)
);

NAND2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1488),
.B(n_472),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1435),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1382),
.B(n_60),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1435),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1433),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1519),
.B(n_473),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1504),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1419),
.B(n_64),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1445),
.B(n_64),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1554),
.B(n_1445),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1604),
.A2(n_1519),
.B1(n_1480),
.B2(n_1458),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1635),
.A2(n_1480),
.B(n_67),
.C(n_65),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1555),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1591),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1526),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1523),
.A2(n_573),
.B(n_478),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1647),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1675),
.A2(n_69),
.B(n_66),
.C(n_68),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1534),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1577),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1533),
.A2(n_479),
.B(n_476),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1541),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1543),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1565),
.A2(n_1574),
.B(n_1539),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1527),
.B(n_482),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1535),
.B(n_68),
.Y(n_1697)
);

O2A1O1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1593),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1577),
.B(n_483),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_SL g1700 ( 
.A1(n_1625),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1531),
.B(n_72),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1524),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1624),
.A2(n_1639),
.B1(n_1676),
.B2(n_1652),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1572),
.B(n_74),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1637),
.B(n_1633),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1529),
.A2(n_485),
.B(n_484),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_76),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1546),
.B(n_77),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1550),
.A2(n_572),
.B(n_487),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1537),
.B(n_77),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1547),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1556),
.A2(n_490),
.B(n_486),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1540),
.B(n_78),
.Y(n_1713)
);

NOR2x1_ASAP7_75t_L g1714 ( 
.A(n_1633),
.B(n_491),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1548),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1525),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1562),
.B(n_79),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1525),
.B(n_80),
.Y(n_1718)
);

BUFx12f_ASAP7_75t_L g1719 ( 
.A(n_1668),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1599),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1575),
.Y(n_1721)
);

NOR2xp67_ASAP7_75t_SL g1722 ( 
.A(n_1579),
.B(n_81),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1549),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1544),
.B(n_1557),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1524),
.B(n_81),
.Y(n_1725)
);

O2A1O1Ixp5_ASAP7_75t_L g1726 ( 
.A1(n_1606),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1564),
.A2(n_570),
.B(n_493),
.Y(n_1727)
);

AOI33xp33_ASAP7_75t_L g1728 ( 
.A1(n_1652),
.A2(n_1677),
.A3(n_1624),
.B1(n_1639),
.B2(n_1588),
.B3(n_1578),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1557),
.B(n_83),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1621),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_SL g1731 ( 
.A1(n_1678),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1619),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1600),
.A2(n_569),
.B(n_494),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1637),
.B(n_88),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1575),
.B(n_89),
.Y(n_1735)
);

O2A1O1Ixp5_ASAP7_75t_L g1736 ( 
.A1(n_1666),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1532),
.A2(n_568),
.B(n_495),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1527),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1676),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1610),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1662),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1676),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1645),
.B(n_95),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1563),
.B(n_96),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1570),
.B(n_97),
.Y(n_1745)
);

NAND2xp33_ASAP7_75t_L g1746 ( 
.A(n_1527),
.B(n_98),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1597),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1612),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1627),
.B(n_101),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1632),
.Y(n_1750)
);

BUFx12f_ASAP7_75t_L g1751 ( 
.A(n_1668),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1643),
.B(n_497),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1660),
.A2(n_566),
.B(n_499),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1673),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1672),
.A2(n_105),
.B1(n_102),
.B2(n_104),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1636),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1626),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1597),
.Y(n_1758)
);

OAI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1655),
.A2(n_104),
.B(n_105),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1616),
.B(n_500),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1567),
.A2(n_565),
.B(n_503),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1569),
.B(n_502),
.Y(n_1762)
);

OAI22x1_ASAP7_75t_L g1763 ( 
.A1(n_1672),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_SL g1764 ( 
.A1(n_1656),
.A2(n_1631),
.B(n_1641),
.C(n_1620),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1545),
.A2(n_109),
.B(n_106),
.C(n_107),
.Y(n_1765)
);

BUFx4f_ASAP7_75t_L g1766 ( 
.A(n_1569),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1605),
.A2(n_564),
.B(n_506),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1582),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1679),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1651),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1545),
.B(n_110),
.Y(n_1771)
);

OAI21xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1642),
.A2(n_509),
.B(n_504),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1589),
.Y(n_1773)
);

BUFx4f_ASAP7_75t_L g1774 ( 
.A(n_1569),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1581),
.B(n_111),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1622),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1659),
.B(n_116),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1538),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1552),
.B(n_118),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1674),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1661),
.A2(n_513),
.B(n_512),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1659),
.B(n_120),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1658),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1566),
.A2(n_1611),
.B(n_1602),
.Y(n_1784)
);

OR2x6_ASAP7_75t_L g1785 ( 
.A(n_1629),
.B(n_514),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1653),
.B(n_122),
.C(n_123),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1584),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1623),
.B(n_124),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1582),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1585),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1790)
);

INVx4_ASAP7_75t_L g1791 ( 
.A(n_1623),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1596),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1613),
.B(n_515),
.Y(n_1793)
);

O2A1O1Ixp33_ASAP7_75t_SL g1794 ( 
.A1(n_1583),
.A2(n_131),
.B(n_128),
.C(n_130),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1646),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_SL g1796 ( 
.A1(n_1664),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1796)
);

NAND2x2_ASAP7_75t_L g1797 ( 
.A(n_1586),
.B(n_1590),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1592),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1559),
.A2(n_517),
.B(n_516),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1651),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1662),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1658),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1598),
.A2(n_1615),
.B1(n_1614),
.B2(n_1580),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1576),
.B(n_134),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1595),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1594),
.B(n_135),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1601),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1542),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_SL g1809 ( 
.A(n_1630),
.B(n_136),
.C(n_137),
.Y(n_1809)
);

BUFx4f_ASAP7_75t_L g1810 ( 
.A(n_1608),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1560),
.B(n_138),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1640),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1595),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1573),
.Y(n_1814)
);

NAND2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1558),
.B(n_520),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1651),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1603),
.B(n_139),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1607),
.B(n_140),
.Y(n_1818)
);

A2O1A1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1561),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1665),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1648),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1644),
.B(n_521),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1568),
.B(n_147),
.C(n_148),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1618),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1530),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1571),
.B(n_147),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1634),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1617),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1698),
.B(n_1657),
.C(n_1587),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1690),
.B(n_1667),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1687),
.Y(n_1831)
);

AO21x2_ASAP7_75t_L g1832 ( 
.A1(n_1695),
.A2(n_1628),
.B(n_1649),
.Y(n_1832)
);

AO22x2_ASAP7_75t_L g1833 ( 
.A1(n_1703),
.A2(n_1609),
.B1(n_1638),
.B2(n_1654),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1705),
.B(n_1803),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1827),
.Y(n_1835)
);

OR2x6_ASAP7_75t_L g1836 ( 
.A(n_1791),
.B(n_1650),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1764),
.A2(n_1669),
.B(n_1671),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1783),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1784),
.A2(n_1663),
.B(n_1551),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1705),
.B(n_1528),
.Y(n_1840)
);

OAI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1728),
.A2(n_1759),
.B(n_1702),
.Y(n_1841)
);

O2A1O1Ixp33_ASAP7_75t_L g1842 ( 
.A1(n_1765),
.A2(n_1528),
.B(n_151),
.C(n_148),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1791),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1825),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1680),
.B(n_1551),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1683),
.B(n_1691),
.Y(n_1846)
);

OR2x6_ASAP7_75t_L g1847 ( 
.A(n_1785),
.B(n_1719),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1785),
.B(n_522),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1756),
.Y(n_1849)
);

AO31x2_ASAP7_75t_L g1850 ( 
.A1(n_1703),
.A2(n_525),
.A3(n_526),
.B(n_524),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1707),
.B(n_527),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1724),
.B(n_530),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1695),
.A2(n_532),
.B(n_531),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1777),
.B(n_534),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1766),
.Y(n_1855)
);

OAI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1706),
.A2(n_537),
.B(n_536),
.Y(n_1856)
);

AOI21x1_ASAP7_75t_L g1857 ( 
.A1(n_1743),
.A2(n_544),
.B(n_538),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1747),
.Y(n_1858)
);

OAI22x1_ASAP7_75t_L g1859 ( 
.A1(n_1684),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1753),
.A2(n_549),
.B(n_545),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1802),
.B(n_150),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1730),
.B(n_152),
.C(n_153),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1735),
.B(n_1704),
.Y(n_1863)
);

CKINVDCx6p67_ASAP7_75t_R g1864 ( 
.A(n_1751),
.Y(n_1864)
);

BUFx2_ASAP7_75t_R g1865 ( 
.A(n_1741),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1806),
.B(n_551),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1814),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1708),
.B(n_153),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1750),
.B(n_1773),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1693),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1726),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1692),
.A2(n_554),
.B(n_553),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1778),
.A2(n_1682),
.B(n_1713),
.C(n_1725),
.Y(n_1873)
);

BUFx4f_ASAP7_75t_L g1874 ( 
.A(n_1747),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1785),
.B(n_155),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1760),
.B(n_1822),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1716),
.B(n_555),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1729),
.B(n_556),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1694),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1779),
.B(n_156),
.Y(n_1880)
);

OAI21x1_ASAP7_75t_L g1881 ( 
.A1(n_1686),
.A2(n_558),
.B(n_557),
.Y(n_1881)
);

INVx5_ASAP7_75t_L g1882 ( 
.A(n_1800),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1782),
.B(n_157),
.Y(n_1883)
);

A2O1A1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1748),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_1884)
);

BUFx4f_ASAP7_75t_L g1885 ( 
.A(n_1747),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1720),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1781),
.A2(n_160),
.B(n_161),
.Y(n_1887)
);

INVx4_ASAP7_75t_SL g1888 ( 
.A(n_1758),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1800),
.Y(n_1889)
);

AOI221x1_ASAP7_75t_L g1890 ( 
.A1(n_1739),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.C(n_164),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_SL g1891 ( 
.A(n_1801),
.B(n_163),
.Y(n_1891)
);

OAI21x1_ASAP7_75t_L g1892 ( 
.A1(n_1709),
.A2(n_164),
.B(n_165),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1811),
.B(n_1809),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1766),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1772),
.A2(n_168),
.B(n_169),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1710),
.B(n_414),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1758),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1727),
.A2(n_168),
.B(n_169),
.Y(n_1898)
);

NOR2xp67_ASAP7_75t_SL g1899 ( 
.A(n_1805),
.B(n_170),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1688),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1712),
.A2(n_172),
.B(n_173),
.Y(n_1901)
);

INVx4_ASAP7_75t_L g1902 ( 
.A(n_1758),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1711),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1810),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1714),
.A2(n_174),
.B(n_175),
.Y(n_1905)
);

AOI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1771),
.A2(n_176),
.B(n_177),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1715),
.Y(n_1907)
);

OA21x2_ASAP7_75t_L g1908 ( 
.A1(n_1736),
.A2(n_177),
.B(n_178),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1742),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_1909)
);

NOR3xp33_ASAP7_75t_L g1910 ( 
.A(n_1739),
.B(n_179),
.C(n_180),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1737),
.A2(n_181),
.B(n_182),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1723),
.Y(n_1912)
);

AO22x2_ASAP7_75t_L g1913 ( 
.A1(n_1780),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1799),
.A2(n_1733),
.B(n_1796),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1794),
.A2(n_184),
.B(n_185),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_R g1916 ( 
.A(n_1828),
.B(n_184),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1767),
.A2(n_186),
.B(n_187),
.Y(n_1917)
);

INVx5_ASAP7_75t_L g1918 ( 
.A(n_1800),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1824),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1740),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1744),
.B(n_186),
.Y(n_1921)
);

OR2x6_ASAP7_75t_L g1922 ( 
.A(n_1813),
.B(n_187),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1697),
.B(n_188),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1732),
.Y(n_1924)
);

OAI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1761),
.A2(n_188),
.B(n_189),
.Y(n_1925)
);

OAI22x1_ASAP7_75t_L g1926 ( 
.A1(n_1792),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1793),
.B(n_1752),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1810),
.Y(n_1928)
);

INVxp67_ASAP7_75t_SL g1929 ( 
.A(n_1685),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1716),
.B(n_192),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1681),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1831),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1882),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1870),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1870),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1879),
.B(n_1757),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1882),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1838),
.B(n_1795),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1846),
.B(n_1689),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1867),
.Y(n_1940)
);

NAND2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1839),
.B(n_1722),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1869),
.B(n_1808),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1882),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1914),
.A2(n_1815),
.B(n_1721),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1876),
.A2(n_1754),
.B(n_1820),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1871),
.A2(n_1819),
.B(n_1775),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1830),
.A2(n_1786),
.B1(n_1798),
.B2(n_1797),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1887),
.A2(n_1835),
.B(n_1892),
.Y(n_1948)
);

NAND3xp33_ASAP7_75t_L g1949 ( 
.A(n_1905),
.B(n_1769),
.C(n_1812),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1834),
.A2(n_1823),
.B1(n_1790),
.B2(n_1787),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1847),
.Y(n_1951)
);

OAI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1837),
.A2(n_1718),
.B(n_1807),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1867),
.Y(n_1953)
);

BUFx12f_ASAP7_75t_L g1954 ( 
.A(n_1928),
.Y(n_1954)
);

INVxp33_ASAP7_75t_L g1955 ( 
.A(n_1849),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1841),
.A2(n_1746),
.B1(n_1776),
.B2(n_1821),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1843),
.B(n_1745),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1903),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1856),
.A2(n_1818),
.B(n_1817),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1903),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1907),
.B(n_1763),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1910),
.A2(n_1755),
.B1(n_1701),
.B2(n_1734),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1927),
.A2(n_1788),
.B1(n_1717),
.B2(n_1755),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1881),
.A2(n_1816),
.B(n_1770),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1912),
.B(n_1749),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1901),
.A2(n_1816),
.B(n_1770),
.Y(n_1966)
);

OAI21x1_ASAP7_75t_L g1967 ( 
.A1(n_1925),
.A2(n_1804),
.B(n_1826),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1922),
.A2(n_1699),
.B1(n_1789),
.B2(n_1768),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1847),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1918),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1865),
.B(n_1738),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1859),
.A2(n_1731),
.B1(n_1700),
.B2(n_196),
.C(n_197),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1924),
.Y(n_1973)
);

A2O1A1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1873),
.A2(n_1774),
.B(n_1762),
.C(n_1696),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_SL g1975 ( 
.A1(n_1913),
.A2(n_1762),
.B1(n_1774),
.B2(n_1738),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1853),
.A2(n_194),
.B(n_195),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1924),
.Y(n_1977)
);

OA21x2_ASAP7_75t_L g1978 ( 
.A1(n_1895),
.A2(n_197),
.B(n_198),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1919),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1844),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_SL g1981 ( 
.A(n_1848),
.B(n_199),
.Y(n_1981)
);

NOR3xp33_ASAP7_75t_L g1982 ( 
.A(n_1862),
.B(n_199),
.C(n_200),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1898),
.A2(n_201),
.B(n_202),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1909),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1844),
.A2(n_203),
.B(n_204),
.Y(n_1985)
);

AO21x2_ASAP7_75t_L g1986 ( 
.A1(n_1915),
.A2(n_204),
.B(n_205),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1918),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1919),
.A2(n_205),
.B(n_206),
.Y(n_1988)
);

OA21x2_ASAP7_75t_L g1989 ( 
.A1(n_1911),
.A2(n_207),
.B(n_208),
.Y(n_1989)
);

AO21x2_ASAP7_75t_L g1990 ( 
.A1(n_1832),
.A2(n_207),
.B(n_209),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1929),
.Y(n_1991)
);

INVx4_ASAP7_75t_L g1992 ( 
.A(n_1848),
.Y(n_1992)
);

NAND2x1p5_ASAP7_75t_L g1993 ( 
.A(n_1875),
.B(n_210),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1864),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1935),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1935),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1944),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1991),
.B(n_1850),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1932),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1944),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1949),
.A2(n_1917),
.B(n_1842),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1982),
.A2(n_1829),
.B1(n_1913),
.B2(n_1893),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1940),
.Y(n_2003)
);

BUFx2_ASAP7_75t_R g2004 ( 
.A(n_1932),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1950),
.A2(n_1926),
.B1(n_1931),
.B2(n_1883),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1945),
.A2(n_1854),
.B1(n_1840),
.B2(n_1833),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1953),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1956),
.A2(n_1896),
.B1(n_1868),
.B2(n_1921),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1963),
.A2(n_1890),
.B1(n_1891),
.B2(n_1922),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1960),
.B(n_1850),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1991),
.Y(n_2011)
);

CKINVDCx20_ASAP7_75t_R g2012 ( 
.A(n_1994),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1973),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1934),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1958),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1952),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_SL g2017 ( 
.A1(n_1992),
.A2(n_1947),
.B1(n_1955),
.B2(n_1951),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1980),
.B(n_1850),
.Y(n_2018)
);

CKINVDCx6p67_ASAP7_75t_R g2019 ( 
.A(n_1954),
.Y(n_2019)
);

BUFx2_ASAP7_75t_R g2020 ( 
.A(n_1933),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1983),
.A2(n_1923),
.B1(n_1899),
.B2(n_1880),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_1951),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1977),
.B(n_1863),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1979),
.Y(n_2024)
);

OR2x6_ASAP7_75t_L g2025 ( 
.A(n_1992),
.B(n_1833),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1962),
.A2(n_1920),
.B1(n_1908),
.B2(n_1861),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1992),
.A2(n_1852),
.B1(n_1872),
.B2(n_1860),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1936),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1984),
.A2(n_1908),
.B1(n_1930),
.B2(n_1851),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1936),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1948),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_1951),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1986),
.A2(n_1930),
.B1(n_1916),
.B2(n_1866),
.Y(n_2033)
);

CKINVDCx6p67_ASAP7_75t_R g2034 ( 
.A(n_2019),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_2001),
.A2(n_1986),
.B1(n_1946),
.B2(n_1975),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1996),
.Y(n_2036)
);

OAI21xp33_ASAP7_75t_L g2037 ( 
.A1(n_2002),
.A2(n_1884),
.B(n_1900),
.Y(n_2037)
);

INVxp67_ASAP7_75t_SL g2038 ( 
.A(n_2003),
.Y(n_2038)
);

BUFx12f_ASAP7_75t_L g2039 ( 
.A(n_1999),
.Y(n_2039)
);

BUFx4f_ASAP7_75t_SL g2040 ( 
.A(n_2012),
.Y(n_2040)
);

OAI22x1_ASAP7_75t_L g2041 ( 
.A1(n_2005),
.A2(n_1993),
.B1(n_1961),
.B2(n_1886),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_SL g2042 ( 
.A1(n_2001),
.A2(n_1981),
.B1(n_1986),
.B2(n_1993),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_2009),
.A2(n_1946),
.B1(n_1969),
.B2(n_1951),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_2009),
.A2(n_1946),
.B1(n_1969),
.B2(n_1951),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_SL g2046 ( 
.A1(n_2017),
.A2(n_1981),
.B1(n_1993),
.B2(n_1978),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2028),
.B(n_1955),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1995),
.Y(n_2048)
);

AOI222xp33_ASAP7_75t_L g2049 ( 
.A1(n_2021),
.A2(n_1968),
.B1(n_1961),
.B2(n_1976),
.C1(n_1974),
.C2(n_1957),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2006),
.A2(n_1969),
.B1(n_1990),
.B2(n_1978),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2005),
.A2(n_1969),
.B1(n_1941),
.B2(n_1845),
.Y(n_2051)
);

CKINVDCx16_ASAP7_75t_R g2052 ( 
.A(n_2017),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_SL g2053 ( 
.A1(n_2025),
.A2(n_1978),
.B1(n_1989),
.B2(n_1990),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_2026),
.A2(n_1969),
.B1(n_1990),
.B2(n_1976),
.Y(n_2054)
);

OAI21xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2021),
.A2(n_1941),
.B(n_1878),
.Y(n_2055)
);

AOI222xp33_ASAP7_75t_L g2056 ( 
.A1(n_2008),
.A2(n_1965),
.B1(n_1967),
.B2(n_1939),
.C1(n_1988),
.C2(n_1942),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_2026),
.A2(n_1989),
.B1(n_1941),
.B2(n_1967),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_SL g2058 ( 
.A1(n_2025),
.A2(n_1989),
.B1(n_1971),
.B2(n_1988),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_2033),
.A2(n_1959),
.B1(n_1836),
.B2(n_1843),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_R g2060 ( 
.A(n_2039),
.B(n_1994),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_2039),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_R g2062 ( 
.A(n_2040),
.B(n_2019),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_2047),
.B(n_2032),
.Y(n_2063)
);

NAND2xp33_ASAP7_75t_R g2064 ( 
.A(n_2052),
.B(n_2022),
.Y(n_2064)
);

NAND2xp33_ASAP7_75t_R g2065 ( 
.A(n_2052),
.B(n_2022),
.Y(n_2065)
);

NAND2xp33_ASAP7_75t_R g2066 ( 
.A(n_2047),
.B(n_2004),
.Y(n_2066)
);

XNOR2xp5_ASAP7_75t_L g2067 ( 
.A(n_2041),
.B(n_1904),
.Y(n_2067)
);

XNOR2xp5_ASAP7_75t_L g2068 ( 
.A(n_2041),
.B(n_2008),
.Y(n_2068)
);

XNOR2xp5_ASAP7_75t_L g2069 ( 
.A(n_2051),
.B(n_2023),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2038),
.B(n_2003),
.Y(n_2070)
);

INVxp67_ASAP7_75t_L g2071 ( 
.A(n_2056),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2034),
.B(n_2023),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2063),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_2061),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2070),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2070),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2064),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2072),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2075),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2074),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2075),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2076),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2078),
.B(n_2068),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_2074),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2077),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2073),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2074),
.B(n_2071),
.Y(n_2087)
);

AND2x6_ASAP7_75t_L g2088 ( 
.A(n_2074),
.B(n_1858),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2081),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_2084),
.B(n_2071),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2079),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2085),
.B(n_2069),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2087),
.B(n_2063),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2082),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2080),
.B(n_2034),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2086),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2087),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2084),
.B(n_2060),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2083),
.B(n_2023),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2088),
.B(n_2044),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_2098),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2090),
.B(n_2088),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2089),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2097),
.B(n_2067),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2093),
.Y(n_2105)
);

NOR2x1p5_ASAP7_75t_SL g2106 ( 
.A(n_2100),
.B(n_2031),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2096),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2092),
.A2(n_2037),
.B(n_2045),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2095),
.B(n_2062),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2109),
.B(n_2090),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2101),
.A2(n_2090),
.B1(n_2037),
.B2(n_2099),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2102),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2105),
.B(n_2099),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2112),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2110),
.B(n_2102),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2111),
.B(n_2103),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2113),
.B(n_2091),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2115),
.B(n_2108),
.Y(n_2118)
);

CKINVDCx20_ASAP7_75t_R g2119 ( 
.A(n_2116),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2114),
.B(n_2108),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2117),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2117),
.B(n_2107),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2114),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2119),
.Y(n_2124)
);

OAI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_2118),
.A2(n_2104),
.B1(n_2094),
.B2(n_2004),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2120),
.A2(n_2088),
.B1(n_2065),
.B2(n_2066),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2123),
.B(n_2019),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2122),
.B(n_1938),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2121),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2122),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2122),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2119),
.A2(n_2046),
.B1(n_2042),
.B2(n_2020),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2122),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_2125),
.A2(n_2106),
.B(n_2049),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2124),
.Y(n_2135)
);

CKINVDCx14_ASAP7_75t_R g2136 ( 
.A(n_2127),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2129),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2130),
.B(n_2088),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2131),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_L g2140 ( 
.A(n_2133),
.B(n_1972),
.C(n_2058),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2128),
.Y(n_2141)
);

AOI21xp33_ASAP7_75t_L g2142 ( 
.A1(n_2132),
.A2(n_1954),
.B(n_210),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2126),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2124),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2124),
.B(n_2055),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2125),
.A2(n_1885),
.B(n_1874),
.Y(n_2146)
);

OAI21xp33_ASAP7_75t_L g2147 ( 
.A1(n_2135),
.A2(n_2020),
.B(n_2033),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2144),
.Y(n_2148)
);

AOI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2142),
.A2(n_2050),
.B1(n_2035),
.B2(n_2057),
.C(n_2054),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_2146),
.A2(n_1885),
.B(n_1874),
.Y(n_2150)
);

AOI211xp5_ASAP7_75t_L g2151 ( 
.A1(n_2143),
.A2(n_1858),
.B(n_1897),
.C(n_1894),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2137),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2138),
.Y(n_2153)
);

OAI211xp5_ASAP7_75t_L g2154 ( 
.A1(n_2136),
.A2(n_2053),
.B(n_1902),
.C(n_1855),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2145),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_2134),
.A2(n_2059),
.B1(n_2029),
.B2(n_1858),
.C(n_2027),
.Y(n_2156)
);

OAI322xp33_ASAP7_75t_L g2157 ( 
.A1(n_2139),
.A2(n_1902),
.A3(n_1998),
.B1(n_213),
.B2(n_214),
.C1(n_215),
.C2(n_216),
.Y(n_2157)
);

OAI21xp33_ASAP7_75t_L g2158 ( 
.A1(n_2140),
.A2(n_2032),
.B(n_1965),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2141),
.B(n_211),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_L g2160 ( 
.A(n_2135),
.B(n_1877),
.C(n_1918),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_SL g2161 ( 
.A(n_2135),
.Y(n_2161)
);

OAI211xp5_ASAP7_75t_L g2162 ( 
.A1(n_2148),
.A2(n_214),
.B(n_211),
.C(n_212),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2147),
.A2(n_2158),
.B1(n_2161),
.B2(n_2155),
.Y(n_2163)
);

O2A1O1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_2157),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_2153),
.A2(n_1888),
.B1(n_2032),
.B2(n_2025),
.Y(n_2165)
);

NOR3xp33_ASAP7_75t_L g2166 ( 
.A(n_2152),
.B(n_1906),
.C(n_1959),
.Y(n_2166)
);

OAI322xp33_ASAP7_75t_L g2167 ( 
.A1(n_2159),
.A2(n_217),
.A3(n_218),
.B1(n_220),
.B2(n_221),
.C1(n_222),
.C2(n_223),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2151),
.B(n_2160),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2150),
.A2(n_1985),
.B(n_1877),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2154),
.B(n_220),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2149),
.A2(n_1888),
.B1(n_2025),
.B2(n_1987),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_SL g2172 ( 
.A1(n_2156),
.A2(n_1937),
.B(n_1933),
.Y(n_2172)
);

AOI211x1_ASAP7_75t_L g2173 ( 
.A1(n_2158),
.A2(n_1857),
.B(n_1998),
.C(n_2048),
.Y(n_2173)
);

OAI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2148),
.A2(n_1985),
.B(n_1952),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2159),
.B(n_222),
.Y(n_2175)
);

OAI221xp5_ASAP7_75t_SL g2176 ( 
.A1(n_2163),
.A2(n_2029),
.B1(n_2025),
.B2(n_1937),
.C(n_1943),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2175),
.B(n_223),
.Y(n_2177)
);

NAND4xp25_ASAP7_75t_L g2178 ( 
.A(n_2164),
.B(n_227),
.C(n_224),
.D(n_226),
.Y(n_2178)
);

OAI211xp5_ASAP7_75t_L g2179 ( 
.A1(n_2170),
.A2(n_227),
.B(n_224),
.C(n_226),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2172),
.A2(n_2168),
.B(n_2162),
.Y(n_2180)
);

OAI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2165),
.A2(n_1970),
.B1(n_1943),
.B2(n_1987),
.Y(n_2181)
);

AOI222xp33_ASAP7_75t_L g2182 ( 
.A1(n_2169),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.C1(n_231),
.C2(n_232),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2166),
.A2(n_1997),
.B1(n_2000),
.B2(n_2025),
.Y(n_2183)
);

NOR3xp33_ASAP7_75t_L g2184 ( 
.A(n_2167),
.B(n_2171),
.C(n_2174),
.Y(n_2184)
);

NOR4xp25_ASAP7_75t_SL g2185 ( 
.A(n_2173),
.B(n_231),
.C(n_228),
.D(n_230),
.Y(n_2185)
);

NOR3xp33_ASAP7_75t_L g2186 ( 
.A(n_2163),
.B(n_232),
.C(n_233),
.Y(n_2186)
);

NAND4xp25_ASAP7_75t_L g2187 ( 
.A(n_2163),
.B(n_236),
.C(n_234),
.D(n_235),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2175),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2164),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.C(n_238),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_L g2190 ( 
.A(n_2163),
.B(n_239),
.C(n_240),
.Y(n_2190)
);

OAI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2163),
.A2(n_1836),
.B1(n_1970),
.B2(n_1889),
.C(n_2011),
.Y(n_2191)
);

AOI221xp5_ASAP7_75t_L g2192 ( 
.A1(n_2164),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.C(n_243),
.Y(n_2192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2193 ( 
.A1(n_2170),
.A2(n_241),
.B(n_242),
.C(n_244),
.D(n_245),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2164),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.C(n_247),
.Y(n_2194)
);

NAND3xp33_ASAP7_75t_SL g2195 ( 
.A(n_2164),
.B(n_247),
.C(n_248),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2162),
.B(n_248),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_L g2197 ( 
.A(n_2163),
.B(n_249),
.C(n_250),
.Y(n_2197)
);

OAI222xp33_ASAP7_75t_L g2198 ( 
.A1(n_2191),
.A2(n_1889),
.B1(n_2043),
.B2(n_2036),
.C1(n_2011),
.C2(n_2048),
.Y(n_2198)
);

AO21x1_ASAP7_75t_L g2199 ( 
.A1(n_2180),
.A2(n_249),
.B(n_250),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2196),
.Y(n_2200)
);

AOI322xp5_ASAP7_75t_L g2201 ( 
.A1(n_2195),
.A2(n_2007),
.A3(n_2043),
.B1(n_2036),
.B2(n_2010),
.C1(n_2018),
.C2(n_2024),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2193),
.A2(n_1966),
.B(n_1964),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2187),
.B(n_251),
.Y(n_2203)
);

NAND3xp33_ASAP7_75t_SL g2204 ( 
.A(n_2189),
.B(n_2194),
.C(n_2192),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_SL g2205 ( 
.A1(n_2179),
.A2(n_251),
.B(n_252),
.Y(n_2205)
);

OAI321xp33_ASAP7_75t_L g2206 ( 
.A1(n_2178),
.A2(n_2181),
.A3(n_2188),
.B1(n_2176),
.B2(n_2183),
.C(n_2177),
.Y(n_2206)
);

AOI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_2186),
.A2(n_2197),
.B1(n_2190),
.B2(n_2184),
.C(n_2185),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_2182),
.B(n_253),
.C(n_254),
.Y(n_2208)
);

AOI221xp5_ASAP7_75t_L g2209 ( 
.A1(n_2181),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.C(n_256),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2181),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.C(n_258),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2180),
.A2(n_258),
.B(n_259),
.Y(n_2211)
);

INVx1_ASAP7_75t_SL g2212 ( 
.A(n_2196),
.Y(n_2212)
);

OAI211xp5_ASAP7_75t_SL g2213 ( 
.A1(n_2180),
.A2(n_260),
.B(n_261),
.C(n_262),
.Y(n_2213)
);

OAI211xp5_ASAP7_75t_SL g2214 ( 
.A1(n_2180),
.A2(n_261),
.B(n_262),
.C(n_264),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2186),
.A2(n_2000),
.B1(n_1997),
.B2(n_2007),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2189),
.B(n_264),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2189),
.B(n_265),
.Y(n_2217)
);

NOR3x1_ASAP7_75t_L g2218 ( 
.A(n_2187),
.B(n_265),
.C(n_266),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2186),
.A2(n_1997),
.B1(n_2000),
.B2(n_2016),
.Y(n_2219)
);

NAND4xp25_ASAP7_75t_L g2220 ( 
.A(n_2189),
.B(n_266),
.C(n_268),
.D(n_269),
.Y(n_2220)
);

AOI211xp5_ASAP7_75t_L g2221 ( 
.A1(n_2179),
.A2(n_269),
.B(n_270),
.C(n_272),
.Y(n_2221)
);

O2A1O1Ixp33_ASAP7_75t_L g2222 ( 
.A1(n_2193),
.A2(n_270),
.B(n_272),
.C(n_273),
.Y(n_2222)
);

AOI211x1_ASAP7_75t_L g2223 ( 
.A1(n_2180),
.A2(n_273),
.B(n_274),
.C(n_275),
.Y(n_2223)
);

AOI322xp5_ASAP7_75t_L g2224 ( 
.A1(n_2195),
.A2(n_2010),
.A3(n_2018),
.B1(n_2024),
.B2(n_2031),
.C1(n_2013),
.C2(n_2015),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2186),
.A2(n_1997),
.B1(n_2000),
.B2(n_2016),
.Y(n_2225)
);

AOI321xp33_ASAP7_75t_L g2226 ( 
.A1(n_2184),
.A2(n_274),
.A3(n_276),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2226)
);

AOI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2181),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2186),
.A2(n_1997),
.B1(n_2000),
.B2(n_2016),
.Y(n_2228)
);

AOI222xp33_ASAP7_75t_L g2229 ( 
.A1(n_2195),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.C1(n_285),
.C2(n_286),
.Y(n_2229)
);

AOI211xp5_ASAP7_75t_L g2230 ( 
.A1(n_2179),
.A2(n_281),
.B(n_284),
.C(n_286),
.Y(n_2230)
);

OAI21xp33_ASAP7_75t_L g2231 ( 
.A1(n_2178),
.A2(n_2000),
.B(n_1997),
.Y(n_2231)
);

NAND5xp2_ASAP7_75t_L g2232 ( 
.A(n_2180),
.B(n_287),
.C(n_288),
.D(n_289),
.E(n_290),
.Y(n_2232)
);

NOR2x1_ASAP7_75t_L g2233 ( 
.A(n_2187),
.B(n_287),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2180),
.A2(n_288),
.B(n_289),
.Y(n_2234)
);

AO22x1_ASAP7_75t_L g2235 ( 
.A1(n_2218),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2226),
.B(n_2199),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2232),
.B(n_291),
.Y(n_2237)
);

NOR2xp67_ASAP7_75t_SL g2238 ( 
.A(n_2211),
.B(n_293),
.Y(n_2238)
);

OAI21xp5_ASAP7_75t_SL g2239 ( 
.A1(n_2205),
.A2(n_2222),
.B(n_2229),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2223),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_L g2241 ( 
.A(n_2221),
.B(n_293),
.C(n_294),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2230),
.B(n_295),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2233),
.Y(n_2243)
);

CKINVDCx16_ASAP7_75t_R g2244 ( 
.A(n_2203),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2234),
.B(n_296),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_L g2246 ( 
.A(n_2209),
.B(n_296),
.C(n_297),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_2213),
.B(n_297),
.Y(n_2247)
);

AOI22x1_ASAP7_75t_L g2248 ( 
.A1(n_2212),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2216),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2217),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2214),
.B(n_299),
.Y(n_2251)
);

NOR4xp25_ASAP7_75t_L g2252 ( 
.A(n_2206),
.B(n_300),
.C(n_301),
.D(n_302),
.Y(n_2252)
);

NOR3xp33_ASAP7_75t_L g2253 ( 
.A(n_2204),
.B(n_301),
.C(n_303),
.Y(n_2253)
);

NAND4xp75_ASAP7_75t_L g2254 ( 
.A(n_2210),
.B(n_304),
.C(n_305),
.D(n_306),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2207),
.B(n_304),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_2220),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2231),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2208),
.B(n_2227),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2200),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2215),
.A2(n_1997),
.B1(n_2000),
.B2(n_2016),
.Y(n_2260)
);

NOR2x1_ASAP7_75t_L g2261 ( 
.A(n_2202),
.B(n_305),
.Y(n_2261)
);

AOI21xp5_ASAP7_75t_L g2262 ( 
.A1(n_2198),
.A2(n_307),
.B(n_308),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2224),
.B(n_2016),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2201),
.B(n_307),
.Y(n_2264)
);

NOR3xp33_ASAP7_75t_L g2265 ( 
.A(n_2219),
.B(n_308),
.C(n_310),
.Y(n_2265)
);

AND4x1_ASAP7_75t_L g2266 ( 
.A(n_2225),
.B(n_310),
.C(n_311),
.D(n_312),
.Y(n_2266)
);

NAND4xp75_ASAP7_75t_L g2267 ( 
.A(n_2255),
.B(n_2228),
.C(n_313),
.D(n_314),
.Y(n_2267)
);

NOR2xp67_ASAP7_75t_L g2268 ( 
.A(n_2241),
.B(n_312),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_L g2269 ( 
.A(n_2244),
.B(n_313),
.C(n_315),
.Y(n_2269)
);

NAND3x1_ASAP7_75t_L g2270 ( 
.A(n_2253),
.B(n_315),
.C(n_316),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2237),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2235),
.Y(n_2272)
);

NOR2x1_ASAP7_75t_L g2273 ( 
.A(n_2243),
.B(n_2245),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2236),
.B(n_316),
.Y(n_2274)
);

NOR2x1_ASAP7_75t_L g2275 ( 
.A(n_2240),
.B(n_317),
.Y(n_2275)
);

NOR3xp33_ASAP7_75t_L g2276 ( 
.A(n_2259),
.B(n_2242),
.C(n_2239),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2238),
.Y(n_2277)
);

NAND2x1p5_ASAP7_75t_L g2278 ( 
.A(n_2266),
.B(n_2248),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2247),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2251),
.Y(n_2280)
);

NOR2x1_ASAP7_75t_L g2281 ( 
.A(n_2239),
.B(n_317),
.Y(n_2281)
);

NOR3xp33_ASAP7_75t_L g2282 ( 
.A(n_2258),
.B(n_318),
.C(n_319),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2256),
.A2(n_2016),
.B1(n_2031),
.B2(n_2018),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2261),
.B(n_2257),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2264),
.Y(n_2285)
);

NOR2x1_ASAP7_75t_L g2286 ( 
.A(n_2254),
.B(n_2246),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2252),
.B(n_318),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2249),
.B(n_319),
.Y(n_2288)
);

NOR2x1p5_ASAP7_75t_L g2289 ( 
.A(n_2250),
.B(n_320),
.Y(n_2289)
);

NOR3x2_ASAP7_75t_L g2290 ( 
.A(n_2265),
.B(n_321),
.C(n_322),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2262),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2263),
.B(n_2260),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2243),
.B(n_321),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_2243),
.B(n_322),
.Y(n_2294)
);

OAI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2252),
.A2(n_323),
.B1(n_324),
.B2(n_326),
.C(n_327),
.Y(n_2295)
);

NAND3x2_ASAP7_75t_L g2296 ( 
.A(n_2237),
.B(n_323),
.C(n_324),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2237),
.Y(n_2297)
);

NOR3x2_ASAP7_75t_L g2298 ( 
.A(n_2254),
.B(n_329),
.C(n_330),
.Y(n_2298)
);

NAND4xp75_ASAP7_75t_L g2299 ( 
.A(n_2255),
.B(n_330),
.C(n_331),
.D(n_332),
.Y(n_2299)
);

NOR2xp67_ASAP7_75t_L g2300 ( 
.A(n_2241),
.B(n_331),
.Y(n_2300)
);

NAND3xp33_ASAP7_75t_L g2301 ( 
.A(n_2253),
.B(n_332),
.C(n_333),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2248),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2237),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2238),
.B(n_334),
.Y(n_2304)
);

AOI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2247),
.A2(n_2016),
.B1(n_2010),
.B2(n_2013),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2248),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_L g2307 ( 
.A(n_2253),
.B(n_334),
.C(n_335),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_L g2308 ( 
.A(n_2253),
.B(n_335),
.C(n_337),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2237),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_L g2310 ( 
.A(n_2255),
.B(n_337),
.C(n_338),
.D(n_339),
.Y(n_2310)
);

OAI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2252),
.A2(n_1966),
.B(n_1964),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2237),
.B(n_338),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2255),
.B(n_339),
.C(n_340),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2293),
.Y(n_2314)
);

INVx1_ASAP7_75t_SL g2315 ( 
.A(n_2298),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2294),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2310),
.B(n_340),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2288),
.Y(n_2318)
);

BUFx12f_ASAP7_75t_L g2319 ( 
.A(n_2304),
.Y(n_2319)
);

NAND3x1_ASAP7_75t_L g2320 ( 
.A(n_2281),
.B(n_341),
.C(n_342),
.Y(n_2320)
);

OA22x2_ASAP7_75t_L g2321 ( 
.A1(n_2272),
.A2(n_2305),
.B1(n_2287),
.B2(n_2277),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2289),
.B(n_341),
.Y(n_2322)
);

OAI211xp5_ASAP7_75t_L g2323 ( 
.A1(n_2296),
.A2(n_342),
.B(n_343),
.C(n_344),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2284),
.B(n_344),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2274),
.B(n_2028),
.Y(n_2325)
);

NOR2x1_ASAP7_75t_L g2326 ( 
.A(n_2275),
.B(n_345),
.Y(n_2326)
);

NOR4xp25_ASAP7_75t_L g2327 ( 
.A(n_2291),
.B(n_345),
.C(n_346),
.D(n_347),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_2270),
.Y(n_2328)
);

NAND4xp75_ASAP7_75t_L g2329 ( 
.A(n_2273),
.B(n_2286),
.C(n_2268),
.D(n_2300),
.Y(n_2329)
);

NOR2xp67_ASAP7_75t_L g2330 ( 
.A(n_2295),
.B(n_346),
.Y(n_2330)
);

NAND5xp2_ASAP7_75t_L g2331 ( 
.A(n_2276),
.B(n_348),
.C(n_349),
.D(n_350),
.E(n_351),
.Y(n_2331)
);

AOI211xp5_ASAP7_75t_L g2332 ( 
.A1(n_2301),
.A2(n_348),
.B(n_349),
.C(n_351),
.Y(n_2332)
);

INVxp33_ASAP7_75t_L g2333 ( 
.A(n_2278),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2269),
.B(n_352),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2284),
.B(n_353),
.Y(n_2335)
);

NOR3xp33_ASAP7_75t_L g2336 ( 
.A(n_2312),
.B(n_353),
.C(n_354),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2293),
.Y(n_2337)
);

NOR2x1_ASAP7_75t_L g2338 ( 
.A(n_2299),
.B(n_355),
.Y(n_2338)
);

NOR3xp33_ASAP7_75t_L g2339 ( 
.A(n_2271),
.B(n_356),
.C(n_357),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2282),
.B(n_356),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2307),
.A2(n_2013),
.B1(n_2014),
.B2(n_2015),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2290),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2313),
.B(n_358),
.Y(n_2343)
);

AND2x2_ASAP7_75t_SL g2344 ( 
.A(n_2302),
.B(n_358),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_2308),
.Y(n_2345)
);

NOR3xp33_ASAP7_75t_L g2346 ( 
.A(n_2297),
.B(n_359),
.C(n_360),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2306),
.B(n_2028),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2303),
.B(n_359),
.Y(n_2348)
);

NAND5xp2_ASAP7_75t_L g2349 ( 
.A(n_2309),
.B(n_361),
.C(n_362),
.D(n_363),
.E(n_364),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2279),
.B(n_362),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2285),
.B(n_2030),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2267),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2280),
.B(n_2030),
.Y(n_2353)
);

NOR2x1_ASAP7_75t_L g2354 ( 
.A(n_2292),
.B(n_365),
.Y(n_2354)
);

AOI221xp5_ASAP7_75t_L g2355 ( 
.A1(n_2292),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.C(n_368),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2283),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2344),
.B(n_2311),
.Y(n_2357)
);

XOR2xp5_ASAP7_75t_L g2358 ( 
.A(n_2333),
.B(n_366),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_SL g2359 ( 
.A(n_2328),
.B(n_367),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2327),
.B(n_368),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2322),
.B(n_369),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_R g2362 ( 
.A(n_2319),
.B(n_369),
.Y(n_2362)
);

NAND2xp33_ASAP7_75t_SL g2363 ( 
.A(n_2316),
.B(n_370),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_R g2364 ( 
.A(n_2337),
.B(n_370),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_R g2365 ( 
.A(n_2337),
.B(n_371),
.Y(n_2365)
);

NAND2xp33_ASAP7_75t_SL g2366 ( 
.A(n_2318),
.B(n_371),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2322),
.B(n_373),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2314),
.B(n_373),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_R g2369 ( 
.A(n_2342),
.B(n_374),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2339),
.B(n_374),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2346),
.B(n_375),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_R g2372 ( 
.A(n_2317),
.B(n_376),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_R g2373 ( 
.A(n_2350),
.B(n_376),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2332),
.B(n_377),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2326),
.B(n_2336),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2354),
.B(n_378),
.Y(n_2376)
);

XNOR2xp5_ASAP7_75t_L g2377 ( 
.A(n_2320),
.B(n_378),
.Y(n_2377)
);

NOR3xp33_ASAP7_75t_SL g2378 ( 
.A(n_2329),
.B(n_379),
.C(n_380),
.Y(n_2378)
);

NAND3xp33_ASAP7_75t_L g2379 ( 
.A(n_2338),
.B(n_2334),
.C(n_2323),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2324),
.B(n_380),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2335),
.B(n_381),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2348),
.B(n_382),
.Y(n_2382)
);

XNOR2xp5_ASAP7_75t_L g2383 ( 
.A(n_2352),
.B(n_382),
.Y(n_2383)
);

NAND3xp33_ASAP7_75t_L g2384 ( 
.A(n_2340),
.B(n_383),
.C(n_384),
.Y(n_2384)
);

NAND2xp33_ASAP7_75t_SL g2385 ( 
.A(n_2343),
.B(n_2356),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2347),
.B(n_384),
.Y(n_2386)
);

NAND3xp33_ASAP7_75t_L g2387 ( 
.A(n_2355),
.B(n_385),
.C(n_386),
.Y(n_2387)
);

NOR3xp33_ASAP7_75t_SL g2388 ( 
.A(n_2331),
.B(n_385),
.C(n_386),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2330),
.B(n_387),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2315),
.B(n_387),
.Y(n_2390)
);

XNOR2xp5_ASAP7_75t_L g2391 ( 
.A(n_2321),
.B(n_2351),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_R g2392 ( 
.A(n_2345),
.B(n_388),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2358),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2383),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2377),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2361),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2376),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2382),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2380),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2381),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2368),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2389),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2390),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2362),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2378),
.B(n_2353),
.Y(n_2405)
);

BUFx12f_ASAP7_75t_L g2406 ( 
.A(n_2391),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_2364),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2379),
.B(n_2325),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2384),
.Y(n_2409)
);

INVx5_ASAP7_75t_L g2410 ( 
.A(n_2359),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2370),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_2388),
.B(n_2349),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2371),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2404),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2405),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2412),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2410),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2410),
.Y(n_2418)
);

XNOR2xp5_ASAP7_75t_L g2419 ( 
.A(n_2393),
.B(n_2360),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2410),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2406),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2408),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2401),
.Y(n_2423)
);

OAI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2407),
.A2(n_2387),
.B1(n_2375),
.B2(n_2357),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2403),
.Y(n_2425)
);

INVxp67_ASAP7_75t_L g2426 ( 
.A(n_2395),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2398),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2394),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2396),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_2409),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2402),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2397),
.A2(n_2374),
.B1(n_2341),
.B2(n_2372),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2399),
.Y(n_2433)
);

OAI22x1_ASAP7_75t_L g2434 ( 
.A1(n_2421),
.A2(n_2400),
.B1(n_2413),
.B2(n_2411),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2417),
.A2(n_2367),
.B(n_2385),
.Y(n_2435)
);

XNOR2xp5_ASAP7_75t_L g2436 ( 
.A(n_2419),
.B(n_2363),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2418),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_L g2438 ( 
.A1(n_2422),
.A2(n_2373),
.B1(n_2369),
.B2(n_2366),
.Y(n_2438)
);

AND2x4_ASAP7_75t_L g2439 ( 
.A(n_2425),
.B(n_2392),
.Y(n_2439)
);

AND2x2_ASAP7_75t_SL g2440 ( 
.A(n_2431),
.B(n_2386),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2414),
.B(n_2365),
.Y(n_2441)
);

OAI21xp5_ASAP7_75t_L g2442 ( 
.A1(n_2426),
.A2(n_388),
.B(n_389),
.Y(n_2442)
);

XNOR2x1_ASAP7_75t_L g2443 ( 
.A(n_2428),
.B(n_389),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2423),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_SL g2445 ( 
.A(n_2416),
.B(n_390),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_2420),
.Y(n_2446)
);

OAI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2435),
.A2(n_2437),
.B(n_2436),
.Y(n_2447)
);

AO22x2_ASAP7_75t_L g2448 ( 
.A1(n_2443),
.A2(n_2432),
.B1(n_2424),
.B2(n_2430),
.Y(n_2448)
);

CKINVDCx20_ASAP7_75t_R g2449 ( 
.A(n_2438),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2446),
.Y(n_2450)
);

INVx1_ASAP7_75t_SL g2451 ( 
.A(n_2440),
.Y(n_2451)
);

CKINVDCx20_ASAP7_75t_R g2452 ( 
.A(n_2449),
.Y(n_2452)
);

OAI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2450),
.A2(n_2429),
.B1(n_2415),
.B2(n_2427),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2451),
.B(n_2445),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_2447),
.A2(n_2439),
.B1(n_2433),
.B2(n_2441),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2452),
.B(n_2442),
.Y(n_2456)
);

OAI22xp33_ASAP7_75t_L g2457 ( 
.A1(n_2454),
.A2(n_2434),
.B1(n_2444),
.B2(n_2448),
.Y(n_2457)
);

AOI221xp5_ASAP7_75t_L g2458 ( 
.A1(n_2453),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.C(n_394),
.Y(n_2458)
);

OAI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2457),
.A2(n_2455),
.B(n_2456),
.Y(n_2459)
);

OAI322xp33_ASAP7_75t_L g2460 ( 
.A1(n_2458),
.A2(n_393),
.A3(n_394),
.B1(n_396),
.B2(n_397),
.C1(n_398),
.C2(n_399),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_L g2461 ( 
.A(n_2456),
.B(n_396),
.Y(n_2461)
);

OAI21x1_ASAP7_75t_L g2462 ( 
.A1(n_2458),
.A2(n_397),
.B(n_400),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2459),
.A2(n_2462),
.B(n_2461),
.Y(n_2463)
);

NAND3xp33_ASAP7_75t_L g2464 ( 
.A(n_2460),
.B(n_400),
.C(n_401),
.Y(n_2464)
);

NAND3xp33_ASAP7_75t_L g2465 ( 
.A(n_2459),
.B(n_401),
.C(n_402),
.Y(n_2465)
);

XNOR2x1_ASAP7_75t_L g2466 ( 
.A(n_2463),
.B(n_402),
.Y(n_2466)
);

AO221x2_ASAP7_75t_L g2467 ( 
.A1(n_2464),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.C(n_406),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2467),
.Y(n_2468)
);

AOI221x1_ASAP7_75t_L g2469 ( 
.A1(n_2468),
.A2(n_2465),
.B1(n_2466),
.B2(n_406),
.C(n_407),
.Y(n_2469)
);

AOI221xp5_ASAP7_75t_L g2470 ( 
.A1(n_2469),
.A2(n_404),
.B1(n_405),
.B2(n_407),
.C(n_408),
.Y(n_2470)
);

AOI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2470),
.A2(n_408),
.B(n_409),
.C(n_410),
.Y(n_2471)
);


endmodule