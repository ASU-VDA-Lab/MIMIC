module fake_jpeg_27011_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx13_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_21),
.Y(n_28)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_11),
.B1(n_21),
.B2(n_23),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_20),
.B(n_16),
.C(n_12),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_10),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_20),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_21),
.B(n_10),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_18),
.B1(n_24),
.B2(n_38),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_6),
.Y(n_53)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_23),
.B(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_49),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_30),
.B1(n_36),
.B2(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_54),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_40),
.B(n_3),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_22),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_43),
.B(n_45),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_59),
.C(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.C(n_22),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_46),
.B(n_47),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_46),
.B1(n_3),
.B2(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_63),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_54),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_5),
.B(n_22),
.C(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_22),
.C(n_18),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_22),
.C(n_1),
.Y(n_70)
);

AOI21x1_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_2),
.Y(n_75)
);


endmodule