module fake_jpeg_2500_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_36),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_14),
.B(n_33),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_44),
.B(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_40),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_37),
.C(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_72),
.C(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_20),
.Y(n_84)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_44),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_39),
.B(n_2),
.C(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_58),
.B(n_42),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_7),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_11),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_72),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_70),
.C(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_71),
.B(n_12),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_16),
.Y(n_106)
);

XOR2x2_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_13),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_112),
.B(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_110),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_91),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_98),
.B1(n_92),
.B2(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_28),
.C(n_29),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_30),
.B(n_31),
.Y(n_112)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_106),
.C(n_116),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_113),
.C(n_111),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_119),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_105),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_124),
.B(n_109),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_115),
.Y(n_129)
);


endmodule