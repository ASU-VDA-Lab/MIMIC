module fake_aes_7978_n_33 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_18;
wire n_32;
wire n_17;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_7), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_12), .B(n_1), .Y(n_18) );
INVxp33_ASAP7_75t_L g19 ( .A(n_9), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_3), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_2), .Y(n_22) );
BUFx4f_ASAP7_75t_L g23 ( .A(n_13), .Y(n_23) );
NOR4xp25_ASAP7_75t_L g24 ( .A(n_20), .B(n_0), .C(n_2), .D(n_4), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_16), .A2(n_5), .B(n_6), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_17), .A2(n_8), .B(n_10), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
OAI21xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_19), .B(n_22), .Y(n_30) );
AOI222xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_18), .B1(n_21), .B2(n_23), .C1(n_24), .C2(n_28), .Y(n_31) );
OAI21x1_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_11), .B(n_15), .Y(n_32) );
AO21x2_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_23), .B(n_21), .Y(n_33) );
endmodule