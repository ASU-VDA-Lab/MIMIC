module real_aes_14556_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_869;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_633;
wire n_482;
wire n_520;
wire n_926;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g694 ( .A(n_0), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_1), .A2(n_547), .B(n_927), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_2), .Y(n_583) );
INVx1_ASAP7_75t_L g140 ( .A(n_3), .Y(n_140) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_3), .A2(n_49), .B(n_142), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_4), .B(n_253), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_5), .B(n_249), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_6), .B(n_208), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_7), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g674 ( .A(n_8), .B(n_236), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_9), .A2(n_92), .B1(n_559), .B2(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_9), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_10), .B(n_267), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_11), .B(n_156), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_12), .B(n_181), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_13), .Y(n_137) );
BUFx3_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
INVx1_ASAP7_75t_L g175 ( .A(n_14), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_15), .B(n_235), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_16), .A2(n_189), .B(n_190), .C(n_192), .Y(n_188) );
BUFx10_ASAP7_75t_L g122 ( .A(n_17), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_18), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_19), .A2(n_124), .B(n_540), .Y(n_123) );
AOI31xp33_ASAP7_75t_L g540 ( .A1(n_19), .A2(n_541), .A3(n_542), .B(n_547), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_20), .B(n_267), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_21), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_22), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_23), .B(n_255), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_24), .A2(n_172), .B(n_176), .C(n_179), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_25), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_26), .B(n_277), .C(n_707), .Y(n_709) );
AND2x2_ASAP7_75t_L g245 ( .A(n_27), .B(n_244), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_28), .B(n_208), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_29), .B(n_235), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_30), .A2(n_74), .B1(n_159), .B2(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g148 ( .A(n_31), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_32), .A2(n_104), .B1(n_118), .B2(n_931), .Y(n_103) );
INVx1_ASAP7_75t_L g212 ( .A(n_33), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_34), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_35), .B(n_159), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_36), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
AND3x2_ASAP7_75t_L g930 ( .A(n_37), .B(n_112), .C(n_554), .Y(n_930) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_38), .B(n_173), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_39), .B(n_189), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_40), .B(n_235), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_41), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_42), .B(n_197), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_43), .Y(n_191) );
AND2x4_ASAP7_75t_L g147 ( .A(n_44), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_45), .B(n_235), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_46), .B(n_244), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_47), .B(n_235), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_48), .A2(n_86), .B1(n_156), .B2(n_159), .Y(n_155) );
INVx1_ASAP7_75t_L g139 ( .A(n_49), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_50), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_51), .A2(n_669), .B(n_693), .C(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g142 ( .A(n_52), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_53), .B(n_235), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_54), .A2(n_557), .B1(n_558), .B2(n_561), .Y(n_556) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_54), .Y(n_561) );
AND2x4_ASAP7_75t_L g109 ( .A(n_55), .B(n_110), .Y(n_109) );
OAI22xp33_ASAP7_75t_L g126 ( .A1(n_56), .A2(n_99), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_56), .Y(n_128) );
INVx3_ASAP7_75t_L g635 ( .A(n_57), .Y(n_635) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_58), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_58), .B(n_76), .Y(n_539) );
AND2x2_ASAP7_75t_L g319 ( .A(n_59), .B(n_236), .Y(n_319) );
INVx1_ASAP7_75t_L g110 ( .A(n_60), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_61), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_62), .B(n_611), .Y(n_616) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_63), .B(n_189), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_64), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g647 ( .A(n_65), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_66), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_67), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g113 ( .A(n_68), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_69), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_70), .B(n_156), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_71), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_72), .B(n_277), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_73), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_75), .B(n_173), .Y(n_318) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_77), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_78), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_79), .B(n_267), .Y(n_278) );
NAND2xp33_ASAP7_75t_SL g205 ( .A(n_80), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_81), .B(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g687 ( .A(n_82), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_83), .B(n_200), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_84), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_85), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
BUFx3_ASAP7_75t_L g181 ( .A(n_87), .Y(n_181) );
INVx1_ASAP7_75t_L g203 ( .A(n_87), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_88), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_89), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_90), .B(n_156), .Y(n_581) );
INVx1_ASAP7_75t_L g633 ( .A(n_91), .Y(n_633) );
INVx1_ASAP7_75t_L g560 ( .A(n_92), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_93), .B(n_265), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_94), .B(n_236), .Y(n_601) );
NAND2xp33_ASAP7_75t_L g226 ( .A(n_95), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_96), .B(n_615), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_97), .Y(n_629) );
INVx1_ASAP7_75t_L g625 ( .A(n_98), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_99), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_100), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_101), .B(n_197), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_102), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g931 ( .A(n_104), .Y(n_931) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_114), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .C(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_111), .B(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g567 ( .A(n_111), .Y(n_567) );
AND2x2_ASAP7_75t_L g553 ( .A(n_112), .B(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g537 ( .A(n_113), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_550), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g552 ( .A(n_121), .B(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_122), .B(n_930), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_533), .Y(n_124) );
INVx1_ASAP7_75t_L g541 ( .A(n_125), .Y(n_541) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
AOI22x1_ASAP7_75t_L g562 ( .A1(n_129), .A2(n_563), .B1(n_568), .B2(n_922), .Y(n_562) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_437), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_346), .C(n_410), .Y(n_130) );
OAI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_238), .B1(n_285), .B2(n_296), .C(n_301), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_166), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g358 ( .A(n_134), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_134), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g446 ( .A(n_134), .B(n_193), .Y(n_446) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g293 ( .A(n_135), .Y(n_293) );
INVx1_ASAP7_75t_L g325 ( .A(n_135), .Y(n_325) );
AND2x2_ASAP7_75t_L g344 ( .A(n_135), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g371 ( .A(n_135), .B(n_361), .Y(n_371) );
INVxp67_ASAP7_75t_L g386 ( .A(n_135), .Y(n_386) );
AND2x2_ASAP7_75t_L g409 ( .A(n_135), .B(n_220), .Y(n_409) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_135), .Y(n_436) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_143), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_138), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_141), .Y(n_138) );
AOI21x1_ASAP7_75t_L g154 ( .A1(n_139), .A2(n_140), .B(n_141), .Y(n_154) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B1(n_161), .B2(n_163), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .C(n_153), .Y(n_144) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_145), .B(n_153), .C(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g673 ( .A(n_145), .Y(n_673) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_146), .A2(n_186), .B(n_691), .Y(n_696) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx6f_ASAP7_75t_SL g218 ( .A(n_147), .Y(n_218) );
INVx1_ASAP7_75t_L g309 ( .A(n_147), .Y(n_309) );
INVx3_ASAP7_75t_L g627 ( .A(n_147), .Y(n_627) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_150), .B(n_627), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_150), .B(n_627), .C(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx3_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_153), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g636 ( .A(n_153), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
INVx2_ASAP7_75t_L g255 ( .A(n_157), .Y(n_255) );
INVx2_ASAP7_75t_L g585 ( .A(n_157), .Y(n_585) );
INVx3_ASAP7_75t_L g661 ( .A(n_157), .Y(n_661) );
INVx3_ASAP7_75t_L g686 ( .A(n_157), .Y(n_686) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_158), .Y(n_160) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_159), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
INVx1_ASAP7_75t_L g277 ( .A(n_160), .Y(n_277) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_162), .A2(n_280), .B(n_281), .C(n_282), .Y(n_279) );
INVx2_ASAP7_75t_L g313 ( .A(n_162), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_162), .A2(n_595), .B(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g200 ( .A(n_165), .Y(n_200) );
INVx2_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
INVx2_ASAP7_75t_L g317 ( .A(n_165), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_166), .A2(n_415), .B(n_419), .Y(n_414) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_193), .Y(n_166) );
AND2x2_ASAP7_75t_L g516 ( .A(n_167), .B(n_409), .Y(n_516) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g289 ( .A(n_169), .Y(n_289) );
INVx1_ASAP7_75t_L g327 ( .A(n_169), .Y(n_327) );
AND2x2_ASAP7_75t_L g355 ( .A(n_169), .B(n_292), .Y(n_355) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_169), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_170), .B(n_187), .Y(n_169) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_170), .B(n_187), .Y(n_345) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_182), .B(n_185), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_172), .A2(n_611), .B1(n_632), .B2(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_173), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g600 ( .A(n_173), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_173), .B(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx3_ASAP7_75t_L g178 ( .A(n_174), .Y(n_178) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx2_ASAP7_75t_L g189 ( .A(n_178), .Y(n_189) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
INVx2_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_178), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_230), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_180), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g209 ( .A(n_181), .Y(n_209) );
INVx1_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
AOI211x1_ASAP7_75t_L g246 ( .A1(n_181), .A2(n_245), .B(n_247), .C(n_251), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_181), .B(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_181), .B(n_627), .C(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g187 ( .A(n_182), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g618 ( .A(n_183), .Y(n_618) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g283 ( .A(n_184), .Y(n_283) );
INVx1_ASAP7_75t_L g587 ( .A(n_184), .Y(n_587) );
INVxp67_ASAP7_75t_L g672 ( .A(n_186), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_192), .A2(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g671 ( .A(n_192), .Y(n_671) );
AND2x2_ASAP7_75t_L g343 ( .A(n_193), .B(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g532 ( .A(n_193), .Y(n_532) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_219), .Y(n_193) );
INVx2_ASAP7_75t_L g292 ( .A(n_194), .Y(n_292) );
AND2x2_ASAP7_75t_L g326 ( .A(n_194), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g337 ( .A(n_194), .Y(n_337) );
OR2x2_ASAP7_75t_L g375 ( .A(n_194), .B(n_345), .Y(n_375) );
AND2x2_ASAP7_75t_L g387 ( .A(n_194), .B(n_345), .Y(n_387) );
AND2x2_ASAP7_75t_L g457 ( .A(n_194), .B(n_220), .Y(n_457) );
AO31x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_204), .A3(n_210), .B(n_215), .Y(n_194) );
AO21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B(n_201), .Y(n_195) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g206 ( .A(n_198), .Y(n_206) );
INVx1_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
INVx2_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
INVx2_ASAP7_75t_L g281 ( .A(n_200), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_201), .A2(n_252), .B(n_254), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_201), .A2(n_264), .B(n_266), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_201), .A2(n_276), .B(n_278), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_201), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_201), .A2(n_598), .B(n_599), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_201), .A2(n_649), .B(n_650), .Y(n_648) );
BUFx10_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g707 ( .A(n_202), .Y(n_707) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx3_ASAP7_75t_L g665 ( .A(n_203), .Y(n_665) );
AO21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_209), .Y(n_204) );
INVx2_ASAP7_75t_L g267 ( .A(n_206), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_209), .A2(n_261), .B(n_262), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_L g582 ( .A1(n_209), .A2(n_583), .B(n_584), .C(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_211), .A2(n_216), .B(n_218), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVxp33_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx2_ASAP7_75t_L g217 ( .A(n_214), .Y(n_217) );
INVx1_ASAP7_75t_L g237 ( .A(n_214), .Y(n_237) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_214), .Y(n_244) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx3_ASAP7_75t_L g221 ( .A(n_217), .Y(n_221) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_218), .A2(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_218), .A2(n_243), .B(n_245), .Y(n_242) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_218), .A2(n_260), .B(n_263), .Y(n_259) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_218), .A2(n_594), .B(n_597), .Y(n_593) );
OAI21x1_ASAP7_75t_L g641 ( .A1(n_218), .A2(n_642), .B(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g295 ( .A(n_220), .Y(n_295) );
INVx1_ASAP7_75t_L g361 ( .A(n_220), .Y(n_361) );
AND2x2_ASAP7_75t_L g383 ( .A(n_220), .B(n_293), .Y(n_383) );
AND2x2_ASAP7_75t_L g466 ( .A(n_220), .B(n_360), .Y(n_466) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_234), .Y(n_220) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_221), .A2(n_578), .B(n_588), .Y(n_577) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_221), .A2(n_641), .B(n_651), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_226), .B(n_228), .Y(n_223) );
INVx2_ASAP7_75t_L g611 ( .A(n_225), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_225), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g615 ( .A(n_227), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_228), .A2(n_316), .B(n_318), .Y(n_315) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_235), .Y(n_700) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_256), .Y(n_238) );
AND2x2_ASAP7_75t_L g389 ( .A(n_239), .B(n_380), .Y(n_389) );
OR2x2_ASAP7_75t_L g405 ( .A(n_239), .B(n_340), .Y(n_405) );
INVx2_ASAP7_75t_L g417 ( .A(n_239), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_239), .B(n_353), .Y(n_420) );
AND2x2_ASAP7_75t_L g517 ( .A(n_239), .B(n_432), .Y(n_517) );
BUFx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g297 ( .A(n_240), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g427 ( .A(n_240), .B(n_332), .Y(n_427) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g320 ( .A(n_241), .B(n_258), .Y(n_320) );
INVx2_ASAP7_75t_L g351 ( .A(n_241), .Y(n_351) );
BUFx2_ASAP7_75t_L g378 ( .A(n_241), .Y(n_378) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_241), .Y(n_395) );
INVx1_ASAP7_75t_L g402 ( .A(n_241), .Y(n_402) );
AND2x2_ASAP7_75t_L g461 ( .A(n_241), .B(n_404), .Y(n_461) );
INVx1_ASAP7_75t_L g522 ( .A(n_241), .Y(n_522) );
OR2x6_ASAP7_75t_L g241 ( .A(n_242), .B(n_246), .Y(n_241) );
INVxp67_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_244), .Y(n_269) );
NOR2xp67_ASAP7_75t_SL g308 ( .A(n_244), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g745 ( .A(n_244), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_250), .Y(n_247) );
INVx2_ASAP7_75t_L g669 ( .A(n_253), .Y(n_669) );
INVxp67_ASAP7_75t_L g643 ( .A(n_255), .Y(n_643) );
INVxp67_ASAP7_75t_L g667 ( .A(n_255), .Y(n_667) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_271), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_257), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g331 ( .A(n_258), .B(n_332), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_268), .B(n_270), .Y(n_258) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_259), .A2(n_268), .B(n_270), .Y(n_300) );
INVx2_ASAP7_75t_L g663 ( .A(n_265), .Y(n_663) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_268), .A2(n_274), .B(n_284), .Y(n_273) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_268), .A2(n_593), .B(n_601), .Y(n_592) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_268), .A2(n_658), .B(n_730), .Y(n_729) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_268), .A2(n_593), .B(n_601), .Y(n_735) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2x1_ASAP7_75t_SL g617 ( .A(n_269), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g487 ( .A(n_271), .Y(n_487) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g404 ( .A(n_272), .Y(n_404) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
INVx1_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_283), .Y(n_274) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_285), .A2(n_411), .B(n_414), .C(n_421), .Y(n_410) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
AND2x2_ASAP7_75t_L g453 ( .A(n_289), .B(n_383), .Y(n_453) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
AND2x2_ASAP7_75t_L g363 ( .A(n_291), .B(n_359), .Y(n_363) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g424 ( .A(n_292), .Y(n_424) );
INVx2_ASAP7_75t_L g397 ( .A(n_294), .Y(n_397) );
BUFx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_295), .Y(n_499) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g353 ( .A(n_298), .B(n_330), .Y(n_353) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g366 ( .A(n_299), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g380 ( .A(n_299), .B(n_306), .Y(n_380) );
AND2x2_ASAP7_75t_L g503 ( .A(n_299), .B(n_330), .Y(n_503) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g341 ( .A(n_300), .B(n_306), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_321), .B1(n_328), .B2(n_333), .C(n_338), .Y(n_301) );
AOI222xp33_ASAP7_75t_L g495 ( .A1(n_302), .A2(n_433), .B1(n_496), .B2(n_501), .C1(n_504), .C2(n_505), .Y(n_495) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2x1_ASAP7_75t_L g303 ( .A(n_304), .B(n_320), .Y(n_303) );
INVx4_ASAP7_75t_R g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_305), .B(n_396), .Y(n_413) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_306), .B(n_330), .Y(n_340) );
AND2x4_ASAP7_75t_L g401 ( .A(n_306), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_314), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_308), .A2(n_315), .B(n_319), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_313), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_313), .A2(n_614), .B(n_616), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_317), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g356 ( .A(n_320), .Y(n_356) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_323), .B(n_509), .C(n_512), .Y(n_508) );
OR2x2_ASAP7_75t_L g524 ( .A(n_323), .B(n_512), .Y(n_524) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_324), .A2(n_394), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g458 ( .A(n_325), .B(n_345), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_326), .B(n_409), .Y(n_429) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
OR2x2_ASAP7_75t_L g472 ( .A(n_329), .B(n_341), .Y(n_472) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g450 ( .A(n_331), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_331), .B(n_377), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_331), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_331), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_331), .B(n_487), .Y(n_515) );
AND2x4_ASAP7_75t_SL g350 ( .A(n_332), .B(n_351), .Y(n_350) );
NOR2x1p5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_337), .B(n_499), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_342), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx4_ASAP7_75t_L g432 ( .A(n_341), .Y(n_432) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_341), .B(n_521), .Y(n_529) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g464 ( .A(n_344), .B(n_457), .Y(n_464) );
INVx2_ASAP7_75t_L g360 ( .A(n_345), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_390), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_368), .C(n_381), .Y(n_347) );
OAI322xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .A3(n_354), .B1(n_356), .B2(n_357), .C1(n_362), .C2(n_364), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g488 ( .A(n_350), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_352), .A2(n_463), .B1(n_465), .B2(n_467), .Y(n_462) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_353), .B(n_401), .Y(n_506) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_355), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g451 ( .A(n_355), .B(n_409), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_355), .B(n_386), .Y(n_527) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g483 ( .A(n_358), .B(n_424), .Y(n_483) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_364), .A2(n_401), .A3(n_422), .B1(n_425), .B2(n_428), .C1(n_430), .C2(n_433), .Y(n_421) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp33_ASAP7_75t_L g426 ( .A(n_365), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
OR2x2_ASAP7_75t_L g441 ( .A(n_366), .B(n_427), .Y(n_441) );
BUFx2_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_376), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_369), .A2(n_399), .B1(n_405), .B2(n_406), .Y(n_398) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g491 ( .A(n_371), .Y(n_491) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g394 ( .A(n_375), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g434 ( .A(n_375), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g474 ( .A(n_375), .B(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g490 ( .A(n_375), .B(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_378), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g449 ( .A(n_378), .Y(n_449) );
OR2x2_ASAP7_75t_L g467 ( .A(n_379), .B(n_403), .Y(n_467) );
OR2x2_ASAP7_75t_L g493 ( .A(n_379), .B(n_487), .Y(n_493) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_388), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_383), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx2_ASAP7_75t_L g512 ( .A(n_387), .Y(n_512) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_397), .B(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_401), .B(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g521 ( .A(n_404), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_406), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_409), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_411), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_417), .B(n_432), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g531 ( .A(n_435), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR3xp33_ASAP7_75t_SL g437 ( .A(n_438), .B(n_479), .C(n_507), .Y(n_437) );
NAND3xp33_ASAP7_75t_SL g438 ( .A(n_439), .B(n_452), .C(n_468), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_447), .B2(n_451), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_446), .A2(n_514), .B1(n_516), .B2(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_456), .B2(n_459), .C(n_462), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g500 ( .A(n_458), .Y(n_500) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp33_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g528 ( .A(n_467), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_473), .B2(n_476), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI211xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_484), .C(n_495), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_483), .A2(n_485), .B1(n_489), .B2(n_492), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g511 ( .A(n_487), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_498), .Y(n_504) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .C(n_518), .D(n_525), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_528), .B1(n_529), .B2(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx12f_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g546 ( .A(n_536), .Y(n_546) );
NOR2x1p5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_539), .Y(n_554) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_SL g548 ( .A(n_546), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_555), .B(n_926), .Y(n_550) );
BUFx8_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_562), .B1(n_924), .B2(n_925), .Y(n_555) );
INVx1_ASAP7_75t_L g924 ( .A(n_556), .Y(n_924) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g925 ( .A(n_562), .Y(n_925) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx8_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
CKINVDCx10_ASAP7_75t_R g923 ( .A(n_565), .Y(n_923) );
BUFx6f_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_848), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_783), .C(n_809), .Y(n_569) );
NAND4xp25_ASAP7_75t_SL g570 ( .A(n_571), .B(n_652), .C(n_739), .D(n_763), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_589), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g911 ( .A(n_573), .Y(n_911) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_574), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g654 ( .A(n_575), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g816 ( .A(n_575), .B(n_725), .Y(n_816) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g722 ( .A(n_576), .B(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g731 ( .A(n_576), .Y(n_731) );
AND2x2_ASAP7_75t_L g840 ( .A(n_576), .B(n_729), .Y(n_840) );
INVx2_ASAP7_75t_L g887 ( .A(n_576), .Y(n_887) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_587), .Y(n_578) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI21x1_ASAP7_75t_L g701 ( .A1(n_587), .A2(n_702), .B(n_705), .Y(n_701) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_602), .Y(n_589) );
OR2x2_ASAP7_75t_L g856 ( .A(n_590), .B(n_681), .Y(n_856) );
AND2x2_ASAP7_75t_L g868 ( .A(n_590), .B(n_869), .Y(n_868) );
BUFx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g753 ( .A(n_591), .Y(n_753) );
AND2x2_ASAP7_75t_L g807 ( .A(n_591), .B(n_736), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_591), .B(n_825), .Y(n_824) );
AND2x4_ASAP7_75t_L g910 ( .A(n_591), .B(n_792), .Y(n_910) );
AND2x2_ASAP7_75t_L g917 ( .A(n_591), .B(n_604), .Y(n_917) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_592), .Y(n_904) );
INVxp67_ASAP7_75t_L g708 ( .A(n_600), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g850 ( .A1(n_602), .A2(n_796), .B(n_851), .C(n_852), .Y(n_850) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_619), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_603), .B(n_821), .Y(n_832) );
OR2x2_ASAP7_75t_L g847 ( .A(n_603), .B(n_824), .Y(n_847) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_603), .Y(n_859) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g795 ( .A(n_604), .Y(n_795) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g680 ( .A(n_605), .Y(n_680) );
BUFx2_ASAP7_75t_L g713 ( .A(n_605), .Y(n_713) );
OR2x2_ASAP7_75t_L g737 ( .A(n_605), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g742 ( .A(n_605), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g842 ( .A(n_605), .B(n_762), .Y(n_842) );
INVx1_ASAP7_75t_L g899 ( .A(n_605), .Y(n_899) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OAI21x1_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_613), .B(n_617), .Y(n_608) );
AND2x2_ASAP7_75t_L g714 ( .A(n_619), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g808 ( .A(n_619), .B(n_801), .Y(n_808) );
AND2x2_ASAP7_75t_L g839 ( .A(n_619), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g873 ( .A(n_619), .Y(n_873) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_638), .Y(n_619) );
INVx1_ASAP7_75t_L g723 ( .A(n_620), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_620), .B(n_885), .Y(n_884) );
AO21x1_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_636), .Y(n_620) );
AO21x2_ASAP7_75t_L g727 ( .A1(n_621), .A2(n_622), .B(n_636), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_631), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_628), .B2(n_630), .Y(n_623) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx3_ASAP7_75t_L g677 ( .A(n_639), .Y(n_677) );
AND2x2_ASAP7_75t_L g750 ( .A(n_639), .B(n_727), .Y(n_750) );
INVx1_ASAP7_75t_L g759 ( .A(n_639), .Y(n_759) );
INVx1_ASAP7_75t_L g765 ( .A(n_639), .Y(n_765) );
AND2x2_ASAP7_75t_L g777 ( .A(n_639), .B(n_726), .Y(n_777) );
AND2x2_ASAP7_75t_L g812 ( .A(n_639), .B(n_729), .Y(n_812) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_639), .Y(n_831) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_645), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_678), .B1(n_711), .B2(n_714), .C(n_718), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_675), .Y(n_653) );
AND2x2_ASAP7_75t_L g764 ( .A(n_654), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g781 ( .A(n_656), .B(n_731), .Y(n_781) );
OR2x2_ASAP7_75t_L g798 ( .A(n_656), .B(n_677), .Y(n_798) );
AO31x2_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_672), .A3(n_673), .B(n_674), .Y(n_656) );
AO31x2_ASAP7_75t_L g717 ( .A1(n_657), .A2(n_672), .A3(n_673), .B(n_674), .Y(n_717) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22x1_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_665), .B1(n_666), .B2(n_671), .Y(n_658) );
OAI22x1_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g695 ( .A(n_665), .Y(n_695) );
AOI21x1_ASAP7_75t_L g702 ( .A1(n_665), .A2(n_703), .B(n_704), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_666) );
AOI21x1_ASAP7_75t_SL g684 ( .A1(n_671), .A2(n_685), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g730 ( .A(n_674), .Y(n_730) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g846 ( .A(n_676), .B(n_828), .Y(n_846) );
NOR2xp67_ASAP7_75t_L g886 ( .A(n_676), .B(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_679), .A2(n_776), .B1(n_778), .B2(n_782), .Y(n_775) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_680), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g767 ( .A(n_680), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_680), .B(n_771), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_680), .B(n_804), .Y(n_803) );
NOR2xp67_ASAP7_75t_R g870 ( .A(n_680), .B(n_871), .Y(n_870) );
OR2x2_ASAP7_75t_L g712 ( .A(n_681), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g752 ( .A(n_681), .B(n_753), .Y(n_752) );
OR2x6_ASAP7_75t_L g681 ( .A(n_682), .B(n_697), .Y(n_681) );
INVx2_ASAP7_75t_L g792 ( .A(n_682), .Y(n_792) );
OR2x2_ASAP7_75t_SL g822 ( .A(n_682), .B(n_743), .Y(n_822) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g736 ( .A(n_683), .Y(n_736) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_690), .B(n_696), .Y(n_683) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_L g770 ( .A(n_697), .B(n_735), .Y(n_770) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_698), .Y(n_738) );
INVx2_ASAP7_75t_L g762 ( .A(n_698), .Y(n_762) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_710), .Y(n_699) );
OA21x2_ASAP7_75t_L g743 ( .A1(n_701), .A2(n_710), .B(n_744), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B(n_709), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g900 ( .A1(n_711), .A2(n_901), .B(n_905), .Y(n_900) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g845 ( .A(n_713), .B(n_807), .Y(n_845) );
OR2x2_ASAP7_75t_L g875 ( .A(n_713), .B(n_761), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_713), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g747 ( .A(n_716), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g757 ( .A(n_716), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g851 ( .A(n_716), .Y(n_851) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g721 ( .A(n_717), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_724), .B(n_732), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g754 ( .A1(n_719), .A2(n_755), .B1(n_757), .B2(n_760), .Y(n_754) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
AND2x2_ASAP7_75t_L g749 ( .A(n_721), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_721), .B(n_777), .Y(n_776) );
OR2x6_ASAP7_75t_L g786 ( .A(n_721), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g801 ( .A(n_721), .Y(n_801) );
INVx1_ASAP7_75t_L g787 ( .A(n_722), .Y(n_787) );
INVx1_ASAP7_75t_L g828 ( .A(n_722), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
INVx1_ASAP7_75t_L g862 ( .A(n_725), .Y(n_862) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_726), .B(n_731), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_726), .B(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g837 ( .A(n_726), .Y(n_837) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_728), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g836 ( .A(n_728), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g874 ( .A(n_728), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_728), .B(n_750), .Y(n_876) );
AND2x2_ASAP7_75t_L g913 ( .A(n_728), .B(n_914), .Y(n_913) );
AND2x4_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g885 ( .A(n_729), .Y(n_885) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_734), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g864 ( .A(n_734), .B(n_795), .Y(n_864) );
INVx1_ASAP7_75t_L g880 ( .A(n_734), .Y(n_880) );
AOI322xp5_ASAP7_75t_L g912 ( .A1(n_734), .A2(n_913), .A3(n_915), .B1(n_917), .B2(n_918), .C1(n_920), .C2(n_921), .Y(n_912) );
AND2x4_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AND2x4_ASAP7_75t_L g791 ( .A(n_735), .B(n_792), .Y(n_791) );
AND2x4_ASAP7_75t_L g841 ( .A(n_735), .B(n_842), .Y(n_841) );
OR2x2_ASAP7_75t_L g853 ( .A(n_735), .B(n_822), .Y(n_853) );
AND2x2_ASAP7_75t_L g756 ( .A(n_736), .B(n_743), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_736), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_736), .Y(n_771) );
INVx1_ASAP7_75t_L g805 ( .A(n_736), .Y(n_805) );
INVx2_ASAP7_75t_L g916 ( .A(n_737), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_746), .B1(n_749), .B2(n_751), .C(n_754), .Y(n_739) );
OR2x2_ASAP7_75t_L g902 ( .A(n_741), .B(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g806 ( .A(n_742), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g909 ( .A(n_742), .B(n_910), .Y(n_909) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g797 ( .A(n_748), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g813 ( .A(n_748), .Y(n_813) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_750), .Y(n_774) );
AND2x2_ASAP7_75t_L g905 ( .A(n_750), .B(n_840), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_751), .A2(n_788), .B1(n_908), .B2(n_909), .Y(n_907) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g760 ( .A(n_753), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g818 ( .A(n_755), .Y(n_818) );
INVxp67_ASAP7_75t_SL g914 ( .A(n_758), .Y(n_914) );
INVx2_ASAP7_75t_L g768 ( .A(n_761), .Y(n_768) );
INVx1_ASAP7_75t_L g825 ( .A(n_762), .Y(n_825) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_762), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B1(n_769), .B2(n_772), .C(n_775), .Y(n_763) );
INVx2_ASAP7_75t_L g780 ( .A(n_765), .Y(n_780) );
AND2x4_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_767), .B(n_791), .Y(n_790) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_768), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_769), .B(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
AND2x2_ASAP7_75t_L g804 ( .A(n_770), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g878 ( .A(n_774), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_777), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_777), .B(n_801), .Y(n_919) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_779), .B(n_862), .Y(n_861) );
NOR2x1p5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g788 ( .A(n_780), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_784), .B(n_799), .Y(n_783) );
AOI32xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_788), .A3(n_789), .B1(n_793), .B2(n_796), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g920 ( .A(n_786), .Y(n_920) );
INVxp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g895 ( .A(n_792), .Y(n_895) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_SL g817 ( .A(n_798), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B1(n_806), .B2(n_808), .Y(n_799) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g871 ( .A(n_805), .Y(n_871) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_807), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_807), .B(n_842), .Y(n_879) );
INVx1_ASAP7_75t_L g896 ( .A(n_808), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_833), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_814), .B1(n_815), .B2(n_818), .C(n_819), .Y(n_810) );
AND2x4_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g827 ( .A(n_812), .Y(n_827) );
AND2x4_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_826), .B1(n_829), .B2(n_832), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_823), .Y(n_820) );
AND2x2_ASAP7_75t_L g921 ( .A(n_821), .B(n_917), .Y(n_921) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g897 ( .A(n_822), .B(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OR2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
OR2x2_ASAP7_75t_L g889 ( .A(n_830), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_841), .B(n_843), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_838), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_835), .A2(n_844), .B1(n_846), .B2(n_847), .Y(n_843) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_SL g865 ( .A(n_846), .Y(n_865) );
NOR3xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_888), .C(n_906), .Y(n_848) );
NAND3xp33_ASAP7_75t_SL g849 ( .A(n_850), .B(n_854), .C(n_863), .Y(n_849) );
INVx3_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OAI31xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_857), .A3(n_858), .B(n_860), .Y(n_854) );
INVx2_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g908 ( .A(n_862), .Y(n_908) );
AOI211xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B(n_866), .C(n_877), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_872), .B1(n_875), .B2(n_876), .Y(n_866) );
NOR2xp33_ASAP7_75t_SL g867 ( .A(n_868), .B(n_870), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_868), .B(n_893), .Y(n_892) );
OR2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_877) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_886), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_883), .B(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g891 ( .A(n_887), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_892), .B1(n_896), .B2(n_897), .C(n_900), .Y(n_888) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_911), .B(n_912), .Y(n_906) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_SL g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
endmodule