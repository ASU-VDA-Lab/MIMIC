module real_jpeg_3216_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_216;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_2),
.A2(n_28),
.B1(n_51),
.B2(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_38),
.B1(n_51),
.B2(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_30),
.C(n_34),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_3),
.B(n_32),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_51),
.C(n_63),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_3),
.B(n_102),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_44),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_45),
.C(n_47),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_3),
.B(n_66),
.Y(n_243)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_59),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_59),
.Y(n_130)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_115),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_114),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_79),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_16),
.B(n_79),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_69),
.B2(n_72),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_126),
.C(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_20),
.A2(n_21),
.B1(n_126),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_20),
.A2(n_21),
.B1(n_91),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_21),
.B(n_91),
.C(n_163),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_23),
.A2(n_70),
.B(n_71),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_25),
.B(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_34),
.B(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_69),
.C(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_68),
.B1(n_74),
.B2(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_54),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_89),
.B(n_106),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_43),
.A2(n_49),
.B1(n_108),
.B2(n_133),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_43),
.A2(n_49),
.B1(n_108),
.B2(n_133),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_49),
.B(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_54),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_47),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

AOI22x1_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_51),
.B(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_66),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_65),
.B(n_78),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_77),
.B(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_72),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_69),
.A2(n_72),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_69),
.A2(n_72),
.B1(n_153),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_72),
.B(n_146),
.C(n_153),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_72),
.B(n_126),
.C(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.C(n_94),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_87),
.B(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_91),
.B(n_187),
.C(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_91),
.A2(n_171),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_109),
.B(n_110),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_96),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_105),
.B1(n_109),
.B2(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_99),
.B(n_150),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_101),
.A2(n_102),
.B1(n_150),
.B2(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_130),
.B(n_149),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_103),
.A2(n_149),
.B(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_134),
.B(n_267),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_117),
.B(n_119),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_126),
.A2(n_142),
.B1(n_179),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_126),
.A2(n_142),
.B1(n_151),
.B2(n_152),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_126),
.B(n_151),
.C(n_250),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_128),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_131),
.A2(n_132),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_131),
.A2(n_132),
.B1(n_216),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_211),
.C(n_216),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_132),
.B(n_168),
.C(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_157),
.B(n_266),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_154),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_138),
.B(n_154),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_145),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_139),
.B(n_143),
.Y(n_264)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_145),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_147),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_151),
.A2(n_152),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_261),
.B(n_265),
.Y(n_157)
);

OAI211xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_190),
.B(n_204),
.C(n_260),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_180),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_172),
.B2(n_173),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_175),
.C(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_167),
.A2(n_168),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_168),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_231),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_186),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_188),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_205),
.C(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_193),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_196),
.C(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_222),
.B(n_259),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_210),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_253),
.B(n_258),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_247),
.B(n_252),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_239),
.B(n_246),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_233),
.B(n_238),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_230),
.B(n_232),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_245),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);


endmodule