module fake_jpeg_13587_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_38),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_36),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_0),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_1),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_101),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_57),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_68),
.B1(n_75),
.B2(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_68),
.B1(n_72),
.B2(n_65),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_52),
.B(n_58),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_54),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_57),
.B(n_58),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_114),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_74),
.B1(n_64),
.B2(n_66),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_120),
.B1(n_5),
.B2(n_6),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_61),
.B1(n_56),
.B2(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_53),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_53),
.C(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_76),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_8),
.C(n_11),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_1),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_3),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_67),
.C(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_133),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_141),
.B(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_4),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_31),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_145),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_5),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_116),
.B(n_124),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_144),
.B(n_12),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_6),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_8),
.B(n_10),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_33),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_49),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_13),
.C(n_14),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_153),
.B1(n_162),
.B2(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_142),
.B1(n_144),
.B2(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_13),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_163),
.B(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_16),
.B1(n_22),
.B2(n_24),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_28),
.B(n_32),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_43),
.B(n_44),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_136),
.C(n_137),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_163),
.B1(n_159),
.B2(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_135),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_173),
.B1(n_155),
.B2(n_157),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_161),
.B1(n_168),
.B2(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_178),
.C(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_172),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_177),
.B1(n_180),
.B2(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_145),
.Y(n_186)
);


endmodule