module real_jpeg_32157_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_29),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_5),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_9),
.B(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_9),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_59),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_35),
.B(n_58),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_30),
.B(n_34),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_42),
.C(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_98),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_84),
.B1(n_96),
.B2(n_97),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_76),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);


endmodule