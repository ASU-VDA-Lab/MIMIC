module real_aes_13060_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
HB1xp67_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_1), .A2(n_16), .B(n_17), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_2), .B(n_10), .Y(n_9) );
INVx2_ASAP7_75t_L g23 ( .A(n_2), .Y(n_23) );
INVx1_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_5), .B(n_8), .Y(n_17) );
A2O1A1O1Ixp25_ASAP7_75t_SL g6 ( .A1(n_7), .A2(n_9), .B(n_11), .C(n_18), .D(n_19), .Y(n_6) );
AOI21xp33_ASAP7_75t_L g12 ( .A1(n_7), .A2(n_13), .B(n_15), .Y(n_12) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
INVx1_ASAP7_75t_L g25 ( .A(n_10), .Y(n_25) );
INVx1_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
BUFx2_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
NOR3xp33_ASAP7_75t_L g20 ( .A(n_14), .B(n_21), .C(n_22), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_18), .B(n_25), .Y(n_24) );
AND2x2_ASAP7_75t_L g19 ( .A(n_20), .B(n_24), .Y(n_19) );
BUFx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
endmodule