module fake_jpeg_677_n_120 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_21),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_8),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_20),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_40),
.B1(n_30),
.B2(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_70),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_57),
.B1(n_56),
.B2(n_14),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_17),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_50),
.B(n_56),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_73),
.B1(n_46),
.B2(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_52),
.B(n_46),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.C(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_74),
.B1(n_61),
.B2(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_57),
.B1(n_52),
.B2(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_69),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_73),
.B1(n_66),
.B2(n_64),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_93),
.B1(n_85),
.B2(n_3),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_82),
.B1(n_83),
.B2(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_63),
.C(n_82),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_80),
.C(n_81),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_84),
.C(n_85),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_86),
.B(n_3),
.Y(n_103)
);

AO221x1_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_2),
.B1(n_6),
.B2(n_9),
.C(n_10),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_100),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_12),
.B(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_107),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_114),
.A2(n_115),
.B1(n_107),
.B2(n_98),
.Y(n_116)
);

NOR2xp67_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_111),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_2),
.B(n_9),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_10),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_12),
.Y(n_120)
);


endmodule