module fake_jpeg_14008_n_566 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_566);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_566;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_63),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

CKINVDCx9p33_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_0),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_29),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_50),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_23),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_107),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_29),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_36),
.Y(n_144)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_47),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_24),
.B1(n_49),
.B2(n_48),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_112),
.A2(n_119),
.B1(n_146),
.B2(n_38),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_65),
.A2(n_39),
.B1(n_33),
.B2(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_125),
.A2(n_165),
.B1(n_88),
.B2(n_66),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_128),
.B(n_133),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_86),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_171),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_70),
.A2(n_39),
.B1(n_49),
.B2(n_47),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_31),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_31),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_43),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_156),
.B(n_166),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_55),
.A2(n_43),
.B1(n_23),
.B2(n_36),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_52),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_73),
.B(n_52),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_108),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_179),
.B(n_180),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_41),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_181),
.Y(n_256)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_183),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_184),
.Y(n_270)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_86),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_187),
.Y(n_276)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_73),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_189),
.Y(n_269)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_40),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_191),
.B(n_192),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_41),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_112),
.A2(n_104),
.B1(n_77),
.B2(n_101),
.Y(n_200)
);

AO22x2_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_89),
.B1(n_100),
.B2(n_84),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_132),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_45),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_206),
.Y(n_241)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_135),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_131),
.B(n_45),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_208),
.B(n_214),
.Y(n_277)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_212),
.B(n_215),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_146),
.A2(n_119),
.B1(n_121),
.B2(n_117),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_226),
.B1(n_155),
.B2(n_139),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_1),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_216),
.B(n_217),
.Y(n_280)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_47),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_219),
.B(n_221),
.Y(n_286)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_220),
.Y(n_258)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_225),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_111),
.B(n_114),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_234),
.B1(n_235),
.B2(n_130),
.Y(n_261)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_149),
.A2(n_164),
.B1(n_82),
.B2(n_103),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_161),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_230),
.B(n_2),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_232),
.B1(n_116),
.B2(n_87),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_58),
.B1(n_64),
.B2(n_81),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_38),
.Y(n_245)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_157),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_116),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_237),
.A2(n_242),
.B1(n_248),
.B2(n_264),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_244),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_168),
.B1(n_159),
.B2(n_164),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_245),
.B(n_15),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_168),
.B1(n_159),
.B2(n_149),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_246),
.A2(n_261),
.B1(n_284),
.B2(n_287),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_123),
.B1(n_114),
.B2(n_155),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_174),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_254),
.B(n_282),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_150),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_257),
.B(n_190),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_47),
.B1(n_38),
.B2(n_3),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_178),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_278),
.A2(n_8),
.B(n_9),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_175),
.B(n_3),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_213),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_226),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_287)
);

OAI22x1_ASAP7_75t_L g288 ( 
.A1(n_200),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_288)
);

OAI22x1_ASAP7_75t_SL g289 ( 
.A1(n_178),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_196),
.A2(n_188),
.B1(n_198),
.B2(n_186),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_254),
.B(n_189),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_298),
.B(n_304),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_187),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_340),
.C(n_268),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_223),
.B(n_177),
.C(n_215),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_R g355 ( 
.A(n_300),
.B(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_261),
.A2(n_234),
.B1(n_195),
.B2(n_217),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_302),
.A2(n_311),
.B1(n_329),
.B2(n_331),
.Y(n_361)
);

NAND2x1_ASAP7_75t_SL g303 ( 
.A(n_245),
.B(n_203),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_326),
.B(n_278),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_240),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_204),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_307),
.Y(n_351)
);

A2O1A1O1Ixp25_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_220),
.B(n_230),
.C(n_194),
.D(n_183),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_228),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_221),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_309),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_253),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_182),
.B1(n_222),
.B2(n_199),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_313),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_216),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_314),
.B(n_316),
.Y(n_369)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_256),
.B(n_211),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_286),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_323),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_269),
.B(n_176),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_291),
.B(n_10),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_332),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_328),
.A2(n_283),
.B1(n_17),
.B2(n_18),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_239),
.B1(n_257),
.B2(n_287),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_256),
.B(n_235),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_239),
.A2(n_257),
.B1(n_288),
.B2(n_265),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_18),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_239),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_334),
.A2(n_259),
.B1(n_281),
.B2(n_255),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_337),
.Y(n_374)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_265),
.B(n_11),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_326),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_276),
.A2(n_11),
.B(n_13),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_243),
.B(n_275),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_11),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_283),
.B(n_275),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_346),
.B(n_378),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_279),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_373),
.C(n_297),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_359),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_333),
.A2(n_239),
.B1(n_257),
.B2(n_264),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_362),
.B1(n_363),
.B2(n_370),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_280),
.B(n_271),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_333),
.A2(n_267),
.B1(n_258),
.B2(n_266),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_292),
.A2(n_267),
.B1(n_258),
.B2(n_266),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_303),
.A2(n_274),
.B(n_243),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_339),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_305),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_382),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_293),
.A2(n_262),
.B1(n_274),
.B2(n_250),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_371),
.A2(n_377),
.B(n_321),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_299),
.B(n_249),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_249),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_380),
.A2(n_384),
.B1(n_327),
.B2(n_341),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_295),
.A2(n_262),
.B1(n_259),
.B2(n_281),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_311),
.B1(n_302),
.B2(n_310),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_307),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_309),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_406),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_387),
.A2(n_391),
.B1(n_392),
.B2(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_395),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_374),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_390),
.B(n_407),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_329),
.B1(n_362),
.B2(n_310),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_343),
.A2(n_296),
.B1(n_331),
.B2(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_325),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_396),
.A2(n_414),
.B(n_385),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_397),
.A2(n_403),
.B1(n_404),
.B2(n_410),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_346),
.C(n_378),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_361),
.A2(n_294),
.B1(n_304),
.B2(n_296),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_345),
.B1(n_343),
.B2(n_347),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_340),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_419),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_344),
.B(n_353),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_375),
.A2(n_313),
.B(n_306),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_409),
.B(n_418),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_345),
.A2(n_294),
.B1(n_296),
.B2(n_332),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_321),
.C(n_301),
.Y(n_411)
);

AOI22x1_ASAP7_75t_L g412 ( 
.A1(n_355),
.A2(n_338),
.B1(n_300),
.B2(n_315),
.Y(n_412)
);

AOI22x1_ASAP7_75t_L g447 ( 
.A1(n_412),
.A2(n_415),
.B1(n_381),
.B2(n_382),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_356),
.A2(n_314),
.B1(n_324),
.B2(n_336),
.Y(n_413)
);

OA22x2_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_322),
.B1(n_318),
.B2(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_417),
.Y(n_424)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_364),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_421),
.Y(n_429)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_401),
.B(n_351),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_449),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_391),
.A2(n_356),
.B1(n_371),
.B2(n_380),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_423),
.B(n_386),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_359),
.B1(n_363),
.B2(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_387),
.A2(n_364),
.B1(n_367),
.B2(n_369),
.Y(n_434)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_377),
.B1(n_376),
.B2(n_370),
.Y(n_436)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_437),
.A2(n_398),
.B(n_414),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

NAND2x1_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_440),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_400),
.B(n_350),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_441),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_413),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_442),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_411),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_389),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_354),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_451),
.C(n_419),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_374),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_386),
.A2(n_367),
.B1(n_377),
.B2(n_379),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_410),
.A2(n_379),
.B1(n_350),
.B2(n_342),
.Y(n_453)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_319),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_396),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_461),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_462),
.A2(n_477),
.B(n_328),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_433),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_463),
.B(n_470),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_427),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_449),
.C(n_426),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_471),
.C(n_476),
.Y(n_483)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_405),
.C(n_398),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_474),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_446),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_481),
.B1(n_448),
.B2(n_444),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_412),
.C(n_414),
.Y(n_476)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_431),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_484),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_457),
.A2(n_425),
.B1(n_428),
.B2(n_436),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_485),
.A2(n_486),
.B1(n_491),
.B2(n_493),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_457),
.A2(n_425),
.B1(n_392),
.B2(n_453),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_445),
.C(n_451),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_468),
.C(n_471),
.Y(n_513)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_488),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_470),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_476),
.B(n_450),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_501),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_456),
.A2(n_432),
.B1(n_447),
.B2(n_423),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_456),
.A2(n_447),
.B1(n_437),
.B2(n_412),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_440),
.B(n_445),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_494),
.A2(n_454),
.B(n_466),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_448),
.B1(n_415),
.B2(n_422),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_495),
.A2(n_499),
.B1(n_474),
.B2(n_473),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_415),
.B1(n_342),
.B2(n_349),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_498),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_466),
.A2(n_415),
.B1(n_342),
.B2(n_439),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_503),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_L g503 ( 
.A1(n_461),
.A2(n_439),
.B(n_317),
.Y(n_503)
);

O2A1O1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_500),
.A2(n_460),
.B(n_467),
.C(n_477),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_479),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_509),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_514),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_492),
.A2(n_460),
.B(n_454),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_522),
.B(n_502),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_515),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_487),
.C(n_483),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_516),
.C(n_513),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_485),
.A2(n_491),
.B1(n_486),
.B2(n_493),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_519),
.A2(n_499),
.B1(n_496),
.B2(n_489),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_495),
.A2(n_462),
.B1(n_458),
.B2(n_481),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_18),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_492),
.A2(n_475),
.B(n_472),
.C(n_459),
.Y(n_522)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_524),
.B(n_526),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_518),
.A2(n_483),
.B(n_494),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_490),
.C(n_472),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_527),
.B(n_528),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_500),
.C(n_497),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_507),
.A2(n_496),
.B(n_497),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_510),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_536),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_512),
.A2(n_482),
.B(n_459),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_533),
.A2(n_534),
.B1(n_535),
.B2(n_506),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_482),
.B(n_17),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_520),
.A2(n_16),
.B(n_18),
.Y(n_535)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_514),
.C(n_517),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_542),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_528),
.A2(n_519),
.B1(n_517),
.B2(n_508),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_537),
.B(n_515),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_543),
.A2(n_525),
.B(n_534),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_533),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_548),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_547),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_510),
.C(n_520),
.Y(n_548)
);

FAx1_ASAP7_75t_SL g550 ( 
.A(n_548),
.B(n_531),
.CI(n_522),
.CON(n_550),
.SN(n_550)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_544),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_546),
.A2(n_531),
.B(n_505),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_552),
.A2(n_532),
.B(n_545),
.Y(n_558)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_553),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_540),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_558),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_559),
.B(n_538),
.Y(n_561)
);

AOI321xp33_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_557),
.A3(n_551),
.B1(n_549),
.B2(n_545),
.C(n_554),
.Y(n_562)
);

NAND4xp25_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_560),
.C(n_552),
.D(n_550),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_563),
.B(n_556),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_541),
.B(n_527),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_565),
.A2(n_542),
.B(n_535),
.Y(n_566)
);


endmodule