module real_jpeg_33239_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_288;
wire n_221;
wire n_249;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_295;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_0),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_0),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_1),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_1),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_1),
.B(n_278),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_3),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_5),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_7),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_7),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_8),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_11),
.B(n_95),
.Y(n_94)
);

NAND2x1_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_113),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_11),
.B(n_219),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_11),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_11),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_120),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_33),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_15),
.B(n_91),
.Y(n_90)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_15),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_15),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_15),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_33),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_16),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_16),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_189),
.B1(n_297),
.B2(n_298),
.Y(n_18)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_19),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_187),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_128),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_23),
.B(n_128),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_72),
.C(n_107),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_24),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_45),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_25),
.B(n_46),
.C(n_56),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.C(n_40),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_26),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_196)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_30),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_30),
.Y(n_204)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_35),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_35),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_44),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_56),
.Y(n_45)
);

OA21x2_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_55),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_148),
.B1(n_149),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_57),
.B(n_67),
.C(n_71),
.Y(n_167)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_65),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_69),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_72),
.B(n_108),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_86),
.C(n_98),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_73),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_80),
.C(n_85),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_86),
.B(n_98),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.C(n_94),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_87),
.B(n_94),
.Y(n_244)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_90),
.B(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_123),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_124),
.C(n_126),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_120),
.B(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_119),
.B(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_154),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_147),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_185),
.B2(n_186),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_168),
.B2(n_169),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_212),
.B(n_296),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_210),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_192),
.B(n_210),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_208),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_193),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_195),
.B(n_208),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.C(n_201),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_197),
.Y(n_238)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_291),
.B(n_295),
.Y(n_212)
);

OAI21x1_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_246),
.B(n_290),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_235),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_235),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_228),
.C(n_234),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_216),
.A2(n_217),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_241),
.C(n_242),
.Y(n_240)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_229),
.B1(n_234),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_233),
.Y(n_266)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_234),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_245),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_240),
.C(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_283),
.B(n_289),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_267),
.B(n_282),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_249),
.B(n_257),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_254),
.Y(n_275)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_276),
.B(n_281),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);


endmodule