module fake_jpeg_8446_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_1),
.Y(n_14)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_14),
.C(n_13),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_8),
.B1(n_15),
.B2(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_6),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_19),
.C(n_17),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_7),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.C(n_7),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_17),
.B(n_24),
.Y(n_29)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_7),
.B(n_15),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_7),
.A3(n_11),
.B1(n_10),
.B2(n_9),
.C1(n_5),
.C2(n_4),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_10),
.C(n_11),
.Y(n_34)
);

AO21x1_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_10),
.Y(n_35)
);

XNOR2x1_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);


endmodule