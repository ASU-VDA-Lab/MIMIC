module fake_jpeg_26144_n_176 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_12),
.B1(n_20),
.B2(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_40),
.B1(n_16),
.B2(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_32),
.C(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_30),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_24),
.B1(n_33),
.B2(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_64),
.B1(n_67),
.B2(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_13),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_15),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_41),
.B1(n_54),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_47),
.B1(n_31),
.B2(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_24),
.B1(n_39),
.B2(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_26),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_28),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_57),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_45),
.B(n_18),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_21),
.CI(n_11),
.CON(n_90),
.SN(n_90)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_74),
.A2(n_93),
.B(n_0),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_81),
.B1(n_86),
.B2(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_15),
.A3(n_14),
.B1(n_13),
.B2(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_52),
.B1(n_33),
.B2(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_18),
.Y(n_82)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_88),
.Y(n_99)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_26),
.B1(n_21),
.B2(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_10),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_72),
.B1(n_58),
.B2(n_65),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_86),
.A3(n_71),
.B1(n_92),
.B2(n_94),
.C1(n_77),
.C2(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_64),
.C(n_68),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_4),
.C(n_5),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_107),
.B1(n_6),
.B2(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_90),
.B1(n_5),
.B2(n_6),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_14),
.B1(n_13),
.B2(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_1),
.B(n_3),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_113),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_3),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_80),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_111),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_79),
.A3(n_90),
.B1(n_82),
.B2(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_135)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_113),
.C(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_107),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_100),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_95),
.C(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_95),
.CI(n_99),
.CON(n_141),
.SN(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_139),
.C(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_136),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_123),
.C(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_149),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_126),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_97),
.C(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_150),
.A2(n_133),
.B(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_104),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_148),
.C(n_143),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_164),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_147),
.B1(n_112),
.B2(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_105),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_141),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_137),
.B(n_140),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_159),
.B(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_163),
.B(n_105),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_168),
.C(n_166),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_9),
.B(n_174),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_9),
.Y(n_176)
);


endmodule