module fake_jpeg_5154_n_282 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_43),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_35),
.B(n_10),
.C(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_49),
.B(n_53),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_59),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_20),
.B1(n_26),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_70),
.B1(n_76),
.B2(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_20),
.B1(n_26),
.B2(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_60),
.A2(n_71),
.B1(n_84),
.B2(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_75),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_32),
.B1(n_17),
.B2(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_32),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_14),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_88),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_38),
.A2(n_14),
.B1(n_28),
.B2(n_16),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_38),
.A2(n_28),
.B1(n_16),
.B2(n_45),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_39),
.A2(n_23),
.B1(n_22),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_97),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_10),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_15),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_15),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_8),
.B(n_9),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_15),
.B1(n_1),
.B2(n_3),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_108),
.B1(n_124),
.B2(n_96),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_5),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_51),
.B1(n_89),
.B2(n_65),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_127),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_76),
.B(n_68),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_147),
.C(n_73),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_129),
.B(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_50),
.Y(n_133)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_85),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_137),
.B1(n_153),
.B2(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_120),
.B1(n_99),
.B2(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_52),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_49),
.B(n_74),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_149),
.B(n_101),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_97),
.B1(n_90),
.B2(n_51),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_146),
.B1(n_151),
.B2(n_105),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_49),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_53),
.C(n_81),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_86),
.B(n_81),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_83),
.B(n_87),
.C(n_59),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_98),
.B1(n_107),
.B2(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_62),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_158),
.Y(n_161)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_62),
.Y(n_158)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_184),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_73),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_173),
.B(n_139),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_174),
.B1(n_157),
.B2(n_100),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_176),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_162),
.B1(n_173),
.B2(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_73),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_112),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_181),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_180),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_188),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_137),
.B(n_139),
.C(n_135),
.D(n_141),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_102),
.C(n_123),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_198),
.B(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_180),
.B1(n_184),
.B2(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_192),
.B1(n_203),
.B2(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_156),
.B1(n_136),
.B2(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_193),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_100),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_122),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_201),
.C(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_132),
.C(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_154),
.C(n_123),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_148),
.B(n_56),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_57),
.B(n_173),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_164),
.B(n_177),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_164),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_176),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_166),
.B1(n_175),
.B2(n_168),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_215),
.B1(n_221),
.B2(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_159),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_200),
.C(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_220),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

OAI322xp33_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_174),
.A3(n_179),
.B1(n_172),
.B2(n_165),
.C1(n_186),
.C2(n_175),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_189),
.C(n_199),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_172),
.B1(n_169),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_197),
.B1(n_206),
.B2(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_224),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_220),
.B(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_194),
.B1(n_191),
.B2(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_243),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_219),
.C(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_198),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_222),
.B1(n_196),
.B2(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_194),
.C(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

AOI31xp67_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_227),
.A3(n_229),
.B(n_214),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_251),
.A3(n_234),
.B(n_240),
.Y(n_261)
);

AOI31xp67_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_225),
.A3(n_190),
.B(n_212),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_167),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_216),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_228),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_236),
.C(n_244),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_260),
.B(n_264),
.Y(n_269)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_239),
.B1(n_233),
.B2(n_231),
.C(n_238),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_236),
.B(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_202),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_267),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_241),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_249),
.B(n_246),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_269),
.B(n_231),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_256),
.C(n_250),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

AOI321xp33_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_274),
.A3(n_257),
.B1(n_277),
.B2(n_256),
.C(n_279),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.C(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_272),
.Y(n_281)
);


endmodule