module fake_netlist_1_293_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_3), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_5), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_8), .B(n_0), .Y(n_12) );
NAND2xp33_ASAP7_75t_R g13 ( .A(n_6), .B(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_12), .B(n_0), .Y(n_15) );
BUFx2_ASAP7_75t_SL g16 ( .A(n_13), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_16), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_14), .B(n_11), .C(n_10), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_9), .Y(n_20) );
BUFx8_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
XNOR2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_4), .Y(n_23) );
endmodule