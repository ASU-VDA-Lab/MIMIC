module fake_jpeg_25312_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_15),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_25),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_41),
.B1(n_35),
.B2(n_16),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_61),
.B1(n_16),
.B2(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_45),
.Y(n_84)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_21),
.B1(n_17),
.B2(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_21),
.B1(n_17),
.B2(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_80),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_36),
.B1(n_45),
.B2(n_33),
.C(n_29),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_18),
.C(n_20),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_63),
.Y(n_108)
);

INVxp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_33),
.B1(n_23),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_25),
.B1(n_23),
.B2(n_29),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_62),
.B1(n_64),
.B2(n_57),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_104),
.B1(n_109),
.B2(n_70),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_37),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_62),
.B1(n_51),
.B2(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_119),
.Y(n_128)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_62),
.B1(n_83),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_43),
.B1(n_51),
.B2(n_92),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_81),
.C(n_77),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_140),
.C(n_143),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_39),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_136),
.B(n_142),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_33),
.A3(n_80),
.B1(n_89),
.B2(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_133),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_132),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_72),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_71),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_150),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_39),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_105),
.B1(n_111),
.B2(n_120),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_70),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_39),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_97),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_147),
.B1(n_122),
.B2(n_50),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_37),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_103),
.C(n_31),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_94),
.B1(n_43),
.B2(n_52),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_59),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_91),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_96),
.B(n_23),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_26),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_154),
.A2(n_166),
.B1(n_181),
.B2(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_159),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_162),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_119),
.B1(n_50),
.B2(n_52),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_158),
.A2(n_124),
.B(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_163),
.B(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_121),
.B1(n_115),
.B2(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_115),
.B1(n_107),
.B2(n_106),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_173),
.B1(n_142),
.B2(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_18),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_103),
.B1(n_86),
.B2(n_26),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_27),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_187),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_103),
.B1(n_86),
.B2(n_31),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_31),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_123),
.B(n_19),
.C(n_20),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_198),
.B1(n_206),
.B2(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_195),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_124),
.C(n_137),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_187),
.C(n_183),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_146),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_208),
.Y(n_224)
);

AO21x1_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_20),
.B(n_151),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_151),
.B1(n_27),
.B2(n_22),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_19),
.B(n_1),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_210),
.B(n_172),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_27),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_22),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_165),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_14),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_214)
);

AO22x2_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_155),
.B1(n_168),
.B2(n_184),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_220),
.B1(n_230),
.B2(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_156),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_181),
.B1(n_170),
.B2(n_186),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_235),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_163),
.B1(n_177),
.B2(n_164),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_180),
.C(n_167),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_205),
.C(n_192),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_157),
.B1(n_172),
.B2(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_185),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_240),
.B1(n_242),
.B2(n_203),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_178),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_160),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_160),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_222),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_250),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_253),
.B1(n_257),
.B2(n_262),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_212),
.C(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_254),
.C(n_256),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_211),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_200),
.B1(n_212),
.B2(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_201),
.C(n_211),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_200),
.C(n_199),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_233),
.B1(n_217),
.B2(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_14),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_204),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_193),
.B(n_190),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_236),
.B(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_210),
.B1(n_197),
.B2(n_214),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_13),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_252),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_231),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_241),
.C(n_239),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_271),
.C(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_220),
.C(n_221),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_272),
.B(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_13),
.C(n_12),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_13),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_7),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_5),
.C(n_6),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_254),
.C(n_248),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_251),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_291),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_245),
.B(n_261),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_266),
.B(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_250),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_295),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_7),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_7),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_265),
.B1(n_268),
.B2(n_275),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_285),
.B1(n_282),
.B2(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_288),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_9),
.B(n_10),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_8),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_310),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_311),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_282),
.B1(n_288),
.B2(n_10),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_8),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_302),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_8),
.C(n_9),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_9),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_299),
.B(n_304),
.Y(n_321)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_320),
.B(n_322),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_310),
.B(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_319),
.B(n_325),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_297),
.C(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_297),
.C(n_9),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_10),
.B(n_318),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule