module fake_jpeg_1222_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_31),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx12_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_28),
.B1(n_32),
.B2(n_20),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_23),
.B1(n_9),
.B2(n_30),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_9),
.B(n_19),
.C(n_18),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_27),
.B(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_3),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_56),
.B1(n_46),
.B2(n_52),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.C(n_34),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_47),
.B1(n_42),
.B2(n_50),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_47),
.B1(n_55),
.B2(n_53),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_58),
.B(n_40),
.C(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_61),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_33),
.B(n_41),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_41),
.Y(n_72)
);


endmodule