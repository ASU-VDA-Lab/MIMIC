module fake_jpeg_1476_n_393 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_55),
.B(n_30),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_63),
.Y(n_117)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_19),
.A2(n_1),
.B(n_3),
.Y(n_62)
);

NAND2x2_ASAP7_75t_SL g169 ( 
.A(n_62),
.B(n_51),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_24),
.B(n_1),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_75),
.Y(n_128)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g170 ( 
.A(n_70),
.Y(n_170)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_98),
.Y(n_115)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_84),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_94),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_5),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_104),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_11),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_32),
.B(n_12),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_36),
.B(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_34),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_110),
.Y(n_120)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_34),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_35),
.B1(n_45),
.B2(n_33),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_116),
.A2(n_145),
.B1(n_158),
.B2(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_30),
.B1(n_33),
.B2(n_53),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_180),
.B1(n_118),
.B2(n_133),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_127),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_53),
.Y(n_127)
);

BUFx2_ASAP7_75t_R g130 ( 
.A(n_55),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_132),
.B(n_133),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_44),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_136),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_44),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_56),
.A2(n_49),
.B1(n_46),
.B2(n_43),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_152),
.Y(n_229)
);

AO22x2_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_49),
.B1(n_46),
.B2(n_43),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_157),
.B(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_58),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_67),
.B(n_51),
.C(n_49),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_132),
.C(n_168),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g168 ( 
.A(n_70),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_168),
.Y(n_182)
);

OR2x2_ASAP7_75t_SL g227 ( 
.A(n_169),
.B(n_62),
.Y(n_227)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_88),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_177),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_66),
.B(n_77),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_85),
.B(n_91),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_92),
.A2(n_73),
.B1(n_79),
.B2(n_74),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_93),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_70),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_92),
.B1(n_177),
.B2(n_149),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_184),
.A2(n_185),
.B1(n_224),
.B2(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_155),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_187),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_128),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_169),
.B1(n_174),
.B2(n_139),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_190),
.A2(n_233),
.B1(n_184),
.B2(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_192),
.B(n_213),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_146),
.B(n_128),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_115),
.B(n_153),
.CI(n_164),
.CON(n_198),
.SN(n_198)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_198),
.B(n_219),
.Y(n_256)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_201),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_150),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_225),
.C(n_182),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_146),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_208),
.B(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_212),
.B(n_200),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_131),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_145),
.B(n_141),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_129),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_122),
.B(n_121),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_137),
.A2(n_123),
.B(n_135),
.C(n_129),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_230),
.B(n_229),
.C(n_200),
.D(n_212),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_160),
.B(n_147),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_223),
.B(n_226),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_156),
.A2(n_165),
.B1(n_163),
.B2(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_138),
.B(n_140),
.C(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_120),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_198),
.C(n_205),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_133),
.B(n_55),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_117),
.B(n_155),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_232),
.B(n_237),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_177),
.B1(n_118),
.B2(n_127),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_238),
.Y(n_254)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_117),
.B(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_197),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_276),
.C(n_224),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_242),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_245),
.A2(n_263),
.B1(n_265),
.B2(n_260),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_246),
.B(n_218),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_234),
.B(n_228),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_190),
.A2(n_229),
.B1(n_185),
.B2(n_202),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_202),
.B1(n_227),
.B2(n_235),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_207),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_206),
.A2(n_225),
.B1(n_201),
.B2(n_182),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_189),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_215),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_221),
.B(n_209),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_220),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_286),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_236),
.B1(n_199),
.B2(n_203),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_295),
.B1(n_303),
.B2(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_284),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_215),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_256),
.B(n_195),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_194),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_241),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_253),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_276),
.B1(n_268),
.B2(n_263),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_275),
.B(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_261),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_248),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_265),
.A2(n_242),
.B1(n_247),
.B2(n_262),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_255),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_267),
.B1(n_271),
.B2(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_272),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_251),
.B(n_243),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_277),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_244),
.B(n_240),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_321),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_324),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_282),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_240),
.B(n_273),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_303),
.B(n_301),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_284),
.B(n_288),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_331),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

AOI22x1_ASAP7_75t_L g331 ( 
.A1(n_321),
.A2(n_308),
.B1(n_305),
.B2(n_302),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_292),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_333),
.C(n_336),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_292),
.C(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_334),
.B(n_335),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_289),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_287),
.C(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_294),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_338),
.B(n_315),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_299),
.C(n_280),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_316),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_297),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_318),
.C(n_319),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_326),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_350),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_349),
.B(n_316),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_320),
.B1(n_322),
.B2(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_354),
.B(n_322),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_332),
.Y(n_359)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_345),
.A2(n_308),
.B1(n_305),
.B2(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_357),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_360),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_333),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_336),
.C(n_340),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_367),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_339),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_363),
.C(n_331),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_341),
.C(n_356),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_368),
.B(n_314),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_369),
.B(n_310),
.Y(n_381)
);

OAI21x1_ASAP7_75t_SL g370 ( 
.A1(n_366),
.A2(n_352),
.B(n_346),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_374),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_367),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_364),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_314),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_361),
.A2(n_358),
.B(n_345),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_376),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_364),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_379),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_381),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_371),
.B(n_310),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_373),
.B(n_362),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_382),
.B(n_376),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_347),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_384),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_383),
.B(n_351),
.Y(n_388)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_388),
.A2(n_389),
.A3(n_324),
.B1(n_323),
.B2(n_363),
.C1(n_358),
.C2(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_390),
.Y(n_393)
);


endmodule