module fake_aes_2809_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_SL g3 ( .A(n_2), .B(n_0), .Y(n_3) );
AOI21x1_ASAP7_75t_L g4 ( .A1(n_2), .A2(n_0), .B(n_1), .Y(n_4) );
CKINVDCx20_ASAP7_75t_R g5 ( .A(n_3), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
BUFx6f_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
OAI221xp5_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_8), .B1(n_1), .B2(n_2), .C(n_0), .Y(n_10) );
NOR3xp33_ASAP7_75t_L g11 ( .A(n_10), .B(n_9), .C(n_1), .Y(n_11) );
AOI211xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_7), .B(n_10), .C(n_8), .Y(n_12) );
NAND2x1p5_ASAP7_75t_L g13 ( .A(n_12), .B(n_7), .Y(n_13) );
endmodule