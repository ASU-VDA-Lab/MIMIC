module fake_jpeg_8995_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_20),
.B1(n_10),
.B2(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_19),
.B1(n_16),
.B2(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_3),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_28),
.C(n_22),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_13),
.C(n_10),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_40),
.C(n_43),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_13),
.C(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_33),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_14),
.C(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_3),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_14),
.B(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_6),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_50),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_52),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_19),
.B1(n_4),
.B2(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_7),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_31),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_8),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_18),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_12),
.C(n_14),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_30),
.B1(n_36),
.B2(n_12),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_36),
.B1(n_12),
.B2(n_14),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_75),
.B(n_76),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_36),
.B1(n_18),
.B2(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_31),
.B1(n_18),
.B2(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_65),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_62),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_61),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_59),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

AO221x1_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_59),
.B1(n_66),
.B2(n_68),
.C(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_70),
.C(n_67),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_80),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_54),
.B(n_63),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_92),
.A3(n_88),
.B1(n_81),
.B2(n_89),
.C1(n_93),
.C2(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_102),
.Y(n_103)
);

XOR2x2_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_81),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_105),
.A3(n_95),
.B1(n_57),
.B2(n_56),
.C1(n_60),
.C2(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_95),
.B1(n_83),
.B2(n_56),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_107),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_104),
.Y(n_109)
);


endmodule