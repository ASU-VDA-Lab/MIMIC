module real_jpeg_11651_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_2),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_52),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_3),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_4),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_4),
.B(n_23),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_4),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_7),
.B(n_52),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_47),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_11),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_12),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_12),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_12),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_33),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_78),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_53),
.B2(n_54),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.C(n_40),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_48),
.B(n_121),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_67),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.C(n_75),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.C(n_87),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_80),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_95),
.C(n_100),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_133),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.CI(n_86),
.CON(n_83),
.SN(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_105),
.B(n_136),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_102),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_130),
.B(n_135),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_118),
.B(n_129),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_116),
.C(n_117),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_124),
.B(n_128),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);


endmodule