module fake_jpeg_14205_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_21),
.C(n_10),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_20),
.B1(n_10),
.B2(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_7),
.B1(n_13),
.B2(n_16),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_16),
.B(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_30),
.B1(n_20),
.B2(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_11),
.B(n_14),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_17),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_41),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_33),
.B1(n_28),
.B2(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_21),
.Y(n_41)
);

MAJx2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_34),
.C(n_41),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_35),
.C(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_51),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.C(n_47),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_15),
.C(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_44),
.B(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI21x1_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_52),
.B(n_56),
.Y(n_58)
);


endmodule