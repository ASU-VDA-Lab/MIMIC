module fake_jpeg_5172_n_147 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_147);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_25),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_39),
.B1(n_44),
.B2(n_54),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_19),
.B1(n_18),
.B2(n_24),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_53),
.B1(n_46),
.B2(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_36),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_53),
.B1(n_56),
.B2(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_81),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_62),
.B(n_65),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_45),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_58),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_73),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_89),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_95),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_67),
.C(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_44),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_53),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_84),
.B(n_83),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_79),
.B1(n_61),
.B2(n_72),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_83),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_71),
.B(n_86),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_76),
.B1(n_70),
.B2(n_78),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_115),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_64),
.B(n_49),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_77),
.B1(n_81),
.B2(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_99),
.B1(n_94),
.B2(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_118),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_80),
.B1(n_64),
.B2(n_16),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_104),
.B1(n_107),
.B2(n_111),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_52),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_41),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_80),
.C(n_75),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_110),
.C(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_131),
.B(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_133),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_103),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_123),
.B1(n_116),
.B2(n_13),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_128),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_2),
.C(n_3),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_126),
.B(n_132),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_135),
.B(n_136),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_134),
.B(n_137),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_142),
.C(n_143),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_2),
.B(n_4),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_7),
.C(n_8),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_9),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_10),
.Y(n_147)
);


endmodule