module real_aes_7087_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_725, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_725;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g466 ( .A1(n_0), .A2(n_204), .B(n_467), .C(n_470), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_1), .B(n_461), .Y(n_471) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g239 ( .A(n_3), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_4), .B(n_156), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_456), .B(n_544), .Y(n_543) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_6), .A2(n_179), .B(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_7), .A2(n_38), .B1(n_149), .B2(n_173), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_8), .B(n_179), .Y(n_251) );
AND2x6_ASAP7_75t_L g164 ( .A(n_9), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_10), .A2(n_164), .B(n_447), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_11), .B(n_39), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_11), .B(n_39), .Y(n_125) );
INVx1_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_13), .B(n_154), .Y(n_187) );
INVx1_ASAP7_75t_L g231 ( .A(n_14), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_15), .A2(n_75), .B1(n_715), .B2(n_716), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_15), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_16), .B(n_156), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_17), .B(n_180), .Y(n_218) );
AO32x2_ASAP7_75t_L g201 ( .A1(n_18), .A2(n_178), .A3(n_179), .B1(n_202), .B2(n_206), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_19), .B(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_20), .B(n_180), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_21), .A2(n_55), .B1(n_149), .B2(n_173), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g176 ( .A1(n_22), .A2(n_82), .B1(n_149), .B2(n_154), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_23), .B(n_149), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_24), .A2(n_178), .B(n_447), .C(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_25), .A2(n_178), .B(n_447), .C(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_26), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_27), .B(n_141), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g701 ( .A1(n_28), .A2(n_94), .B1(n_702), .B2(n_703), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_28), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_29), .A2(n_700), .B1(n_701), .B2(n_704), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_29), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_30), .A2(n_456), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_31), .B(n_141), .Y(n_166) );
INVx2_ASAP7_75t_L g151 ( .A(n_32), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_33), .A2(n_453), .B(n_479), .C(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_34), .B(n_149), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_35), .B(n_141), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_36), .A2(n_43), .B1(n_437), .B2(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_36), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_37), .B(n_189), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_40), .B(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_41), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_42), .B(n_156), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_43), .A2(n_132), .B1(n_437), .B2(n_438), .Y(n_131) );
INVx1_ASAP7_75t_L g437 ( .A(n_43), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_44), .B(n_456), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_45), .A2(n_453), .B(n_479), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_46), .B(n_149), .Y(n_246) );
INVx1_ASAP7_75t_L g468 ( .A(n_47), .Y(n_468) );
AOI22xp5_ASAP7_75t_SL g127 ( .A1(n_48), .A2(n_123), .B1(n_128), .B2(n_707), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_49), .A2(n_92), .B1(n_173), .B2(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g531 ( .A(n_50), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_51), .B(n_149), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_52), .B(n_149), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_53), .B(n_456), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_54), .B(n_237), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_56), .A2(n_60), .B1(n_149), .B2(n_154), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_57), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_58), .B(n_149), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_59), .B(n_149), .Y(n_259) );
INVx1_ASAP7_75t_L g165 ( .A(n_61), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_62), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_63), .B(n_461), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_64), .A2(n_234), .B(n_237), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_65), .B(n_149), .Y(n_240) );
INVx1_ASAP7_75t_L g144 ( .A(n_66), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_68), .B(n_156), .Y(n_484) );
AO32x2_ASAP7_75t_L g170 ( .A1(n_69), .A2(n_171), .A3(n_177), .B1(n_178), .B2(n_179), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_70), .B(n_157), .Y(n_521) );
INVx1_ASAP7_75t_L g258 ( .A(n_71), .Y(n_258) );
INVx1_ASAP7_75t_L g152 ( .A(n_72), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_73), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_74), .B(n_483), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_75), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_76), .A2(n_447), .B(n_449), .C(n_453), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_77), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_78), .B(n_154), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_79), .Y(n_545) );
INVx1_ASAP7_75t_L g114 ( .A(n_80), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_81), .B(n_482), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_83), .B(n_173), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_84), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_85), .B(n_154), .Y(n_161) );
INVx2_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_87), .A2(n_105), .B1(n_115), .B2(n_722), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_88), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_89), .B(n_175), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_90), .B(n_154), .Y(n_247) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_91), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g122 ( .A(n_91), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_93), .A2(n_103), .B1(n_154), .B2(n_155), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_94), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_95), .B(n_456), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_96), .Y(n_481) );
INVxp67_ASAP7_75t_L g548 ( .A(n_97), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_98), .B(n_154), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g450 ( .A(n_100), .Y(n_450) );
INVx1_ASAP7_75t_L g517 ( .A(n_101), .Y(n_517) );
AND2x2_ASAP7_75t_L g533 ( .A(n_102), .B(n_141), .Y(n_533) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g723 ( .A(n_108), .Y(n_723) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g124 ( .A(n_111), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_127), .B1(n_710), .B2(n_711), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g710 ( .A(n_118), .Y(n_710) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_120), .A2(n_712), .B(n_721), .Y(n_711) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g721 ( .A(n_122), .Y(n_721) );
NOR2x2_ASAP7_75t_L g709 ( .A(n_123), .B(n_130), .Y(n_709) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp33_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_699), .B1(n_705), .B2(n_706), .Y(n_128) );
INVx1_ASAP7_75t_L g705 ( .A(n_129), .Y(n_705) );
AO22x2_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_131), .B1(n_439), .B2(n_698), .Y(n_129) );
INVx1_ASAP7_75t_L g698 ( .A(n_130), .Y(n_698) );
INVx1_ASAP7_75t_L g438 ( .A(n_132), .Y(n_438) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_132), .A2(n_438), .B1(n_718), .B2(n_719), .Y(n_717) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_358), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_307), .C(n_349), .Y(n_133) );
AOI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_212), .B(n_261), .C(n_283), .Y(n_134) );
OAI211xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_167), .B(n_195), .C(n_207), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_137), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g370 ( .A(n_137), .B(n_287), .Y(n_370) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g272 ( .A(n_138), .B(n_198), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_138), .B(n_183), .Y(n_389) );
INVx1_ASAP7_75t_L g407 ( .A(n_138), .Y(n_407) );
AND2x2_ASAP7_75t_L g416 ( .A(n_138), .B(n_304), .Y(n_416) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g299 ( .A(n_139), .B(n_183), .Y(n_299) );
AND2x2_ASAP7_75t_L g357 ( .A(n_139), .B(n_304), .Y(n_357) );
INVx1_ASAP7_75t_L g401 ( .A(n_139), .Y(n_401) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g278 ( .A(n_140), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g286 ( .A(n_140), .Y(n_286) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_140), .Y(n_326) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_166), .Y(n_140) );
INVx2_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_141), .A2(n_184), .B(n_194), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_141), .A2(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g500 ( .A(n_141), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_141), .A2(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g180 ( .A(n_142), .B(n_143), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_159), .B(n_164), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_SL g147 ( .A1(n_148), .A2(n_152), .B(n_153), .C(n_156), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_149), .Y(n_452) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
AND2x6_ASAP7_75t_L g447 ( .A(n_150), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g155 ( .A(n_151), .Y(n_155) );
INVx1_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
INVx2_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_156), .A2(n_246), .B(n_247), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_156), .A2(n_255), .B(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_156), .B(n_548), .Y(n_547) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_157), .A2(n_172), .B1(n_175), .B2(n_176), .Y(n_171) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_158), .Y(n_163) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx1_ASAP7_75t_L g448 ( .A(n_158), .Y(n_448) );
AND2x2_ASAP7_75t_L g457 ( .A(n_158), .B(n_238), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g234 ( .A(n_162), .Y(n_234) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g483 ( .A(n_163), .Y(n_483) );
BUFx3_ASAP7_75t_L g178 ( .A(n_164), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_164), .A2(n_185), .B(n_190), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_164), .A2(n_230), .B(n_235), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_164), .A2(n_245), .B(n_248), .Y(n_244) );
INVx4_ASAP7_75t_SL g454 ( .A(n_164), .Y(n_454) );
AND2x4_ASAP7_75t_L g456 ( .A(n_164), .B(n_457), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_164), .B(n_457), .Y(n_518) );
INVxp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_181), .Y(n_168) );
AND2x2_ASAP7_75t_L g265 ( .A(n_169), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g298 ( .A(n_169), .Y(n_298) );
OR2x2_ASAP7_75t_L g424 ( .A(n_169), .B(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_169), .B(n_183), .Y(n_428) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
INVx1_ASAP7_75t_L g210 ( .A(n_170), .Y(n_210) );
AND2x2_ASAP7_75t_L g287 ( .A(n_170), .B(n_200), .Y(n_287) );
AND2x2_ASAP7_75t_L g327 ( .A(n_170), .B(n_201), .Y(n_327) );
INVx2_ASAP7_75t_L g470 ( .A(n_174), .Y(n_470) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_174), .Y(n_485) );
INVx2_ASAP7_75t_L g193 ( .A(n_175), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_175), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_175), .A2(n_204), .B1(n_221), .B2(n_222), .Y(n_220) );
INVx4_ASAP7_75t_L g469 ( .A(n_175), .Y(n_469) );
INVx1_ASAP7_75t_L g497 ( .A(n_177), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_178), .B(n_220), .C(n_223), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_178), .A2(n_254), .B(n_257), .Y(n_253) );
INVx4_ASAP7_75t_L g223 ( .A(n_179), .Y(n_223) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_179), .A2(n_244), .B(n_251), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_179), .A2(n_507), .B(n_508), .Y(n_506) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_179), .Y(n_542) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g206 ( .A(n_180), .Y(n_206) );
INVxp67_ASAP7_75t_L g369 ( .A(n_181), .Y(n_369) );
AND2x4_ASAP7_75t_L g394 ( .A(n_181), .B(n_287), .Y(n_394) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_182), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g199 ( .A(n_183), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g273 ( .A(n_183), .B(n_201), .Y(n_273) );
INVx1_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
INVx2_ASAP7_75t_L g305 ( .A(n_183), .Y(n_305) );
AND2x2_ASAP7_75t_L g321 ( .A(n_183), .B(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .Y(n_185) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
O2A1O1Ixp5_ASAP7_75t_L g257 ( .A1(n_193), .A2(n_236), .B(n_258), .C(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_196), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g276 ( .A(n_198), .Y(n_276) );
AND2x2_ASAP7_75t_L g384 ( .A(n_198), .B(n_200), .Y(n_384) );
AND2x2_ASAP7_75t_L g301 ( .A(n_199), .B(n_286), .Y(n_301) );
AND2x2_ASAP7_75t_L g400 ( .A(n_199), .B(n_401), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_200), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g425 ( .A(n_200), .B(n_286), .Y(n_425) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g211 ( .A(n_201), .Y(n_211) );
AND2x2_ASAP7_75t_L g304 ( .A(n_201), .B(n_305), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_204), .A2(n_236), .B(n_239), .C(n_240), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_204), .A2(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g228 ( .A(n_206), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_206), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
AND2x2_ASAP7_75t_L g350 ( .A(n_209), .B(n_285), .Y(n_350) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_210), .B(n_286), .Y(n_335) );
INVx2_ASAP7_75t_L g334 ( .A(n_211), .Y(n_334) );
OAI222xp33_ASAP7_75t_L g338 ( .A1(n_211), .A2(n_278), .B1(n_339), .B2(n_341), .C1(n_342), .C2(n_345), .Y(n_338) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g263 ( .A(n_216), .Y(n_263) );
OR2x2_ASAP7_75t_L g374 ( .A(n_216), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g296 ( .A(n_217), .Y(n_296) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_217), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_217), .B(n_267), .Y(n_353) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
AO21x1_ASAP7_75t_L g313 ( .A1(n_220), .A2(n_223), .B(n_314), .Y(n_313) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_223), .A2(n_445), .B(n_458), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_223), .B(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g461 ( .A(n_223), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_223), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_223), .A2(n_516), .B(n_523), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_224), .A2(n_317), .B1(n_356), .B2(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_242), .Y(n_224) );
INVx3_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
OR2x2_ASAP7_75t_L g422 ( .A(n_225), .B(n_298), .Y(n_422) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g295 ( .A(n_226), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_226), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_226), .B(n_267), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_226), .B(n_243), .Y(n_375) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g266 ( .A(n_227), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g270 ( .A(n_227), .B(n_243), .Y(n_270) );
AND2x2_ASAP7_75t_L g346 ( .A(n_227), .B(n_293), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_227), .B(n_252), .Y(n_386) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_241), .Y(n_227) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_228), .A2(n_253), .B(n_260), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .C(n_234), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_232), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_232), .A2(n_521), .B(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_234), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_236), .A2(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_242), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g302 ( .A(n_242), .B(n_263), .Y(n_302) );
AND2x2_ASAP7_75t_L g306 ( .A(n_242), .B(n_296), .Y(n_306) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
INVx3_ASAP7_75t_L g267 ( .A(n_243), .Y(n_267) );
AND2x2_ASAP7_75t_L g292 ( .A(n_243), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g427 ( .A(n_243), .B(n_410), .Y(n_427) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
INVx2_ASAP7_75t_L g293 ( .A(n_252), .Y(n_293) );
AND2x2_ASAP7_75t_L g337 ( .A(n_252), .B(n_313), .Y(n_337) );
INVx1_ASAP7_75t_L g380 ( .A(n_252), .Y(n_380) );
OR2x2_ASAP7_75t_L g411 ( .A(n_252), .B(n_313), .Y(n_411) );
AND2x2_ASAP7_75t_L g431 ( .A(n_252), .B(n_267), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_268), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g269 ( .A(n_263), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_263), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g388 ( .A(n_265), .Y(n_388) );
INVx2_ASAP7_75t_SL g282 ( .A(n_266), .Y(n_282) );
AND2x2_ASAP7_75t_L g402 ( .A(n_266), .B(n_296), .Y(n_402) );
INVx2_ASAP7_75t_L g348 ( .A(n_267), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_267), .B(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B1(n_274), .B2(n_280), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_270), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g436 ( .A(n_270), .Y(n_436) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g361 ( .A(n_272), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_272), .B(n_304), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_273), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g377 ( .A(n_273), .B(n_326), .Y(n_377) );
INVx2_ASAP7_75t_L g433 ( .A(n_273), .Y(n_433) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_276), .B(n_321), .Y(n_354) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_278), .B(n_298), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g415 ( .A(n_281), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_SL g365 ( .A1(n_282), .A2(n_366), .B(n_368), .C(n_371), .Y(n_365) );
OR2x2_ASAP7_75t_L g392 ( .A(n_282), .B(n_296), .Y(n_392) );
OAI221xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_288), .B1(n_290), .B2(n_297), .C(n_300), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_285), .B(n_334), .Y(n_341) );
AND2x2_ASAP7_75t_L g383 ( .A(n_285), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g419 ( .A(n_285), .Y(n_419) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
INVx1_ASAP7_75t_L g323 ( .A(n_286), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_289), .B(n_344), .Y(n_343) );
INVxp67_ASAP7_75t_L g397 ( .A(n_289), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_289), .B(n_337), .Y(n_413) );
INVx2_ASAP7_75t_L g399 ( .A(n_290), .Y(n_399) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g340 ( .A(n_292), .B(n_311), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_292), .A2(n_308), .B(n_350), .C(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g318 ( .A(n_293), .B(n_313), .Y(n_318) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_297), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g366 ( .A(n_298), .B(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_303), .B2(n_306), .Y(n_300) );
INVx1_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
INVx1_ASAP7_75t_L g367 ( .A(n_304), .Y(n_367) );
INVx1_ASAP7_75t_L g418 ( .A(n_306), .Y(n_418) );
AOI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_311), .B(n_315), .C(n_338), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g330 ( .A(n_310), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g381 ( .A(n_311), .Y(n_381) );
AND2x2_ASAP7_75t_L g430 ( .A(n_311), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI21xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B(n_328), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_318), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g336 ( .A(n_319), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g412 ( .A(n_319), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_319), .A2(n_371), .A3(n_378), .B1(n_419), .B2(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_SL g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_SL g391 ( .A(n_321), .Y(n_391) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g331 ( .A(n_327), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B(n_336), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_330), .A2(n_378), .B1(n_404), .B2(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_334), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g364 ( .A(n_348), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_399), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_398) );
NAND5xp2_ASAP7_75t_L g358 ( .A(n_359), .B(n_382), .C(n_398), .D(n_408), .E(n_426), .Y(n_358) );
AOI211xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_365), .C(n_372), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g429 ( .A(n_366), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_376), .B2(n_378), .Y(n_372) );
INVx1_ASAP7_75t_SL g405 ( .A(n_375), .Y(n_405) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI322xp33_ASAP7_75t_L g387 ( .A1(n_378), .A2(n_388), .A3(n_389), .B1(n_390), .B2(n_391), .C1(n_392), .C2(n_393), .Y(n_387) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g390 ( .A(n_380), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_380), .B(n_405), .Y(n_404) );
AOI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_387), .C(n_395), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_391), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_416), .B1(n_417), .B2(n_421), .C(n_423), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_412), .B(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g435 ( .A(n_411), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_429), .B2(n_430), .C(n_432), .Y(n_426) );
AOI21xp33_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_641), .Y(n_439) );
AND4x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_581), .C(n_596), .D(n_621), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g441 ( .A(n_442), .B(n_554), .Y(n_441) );
OAI21xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_472), .B(n_534), .Y(n_442) );
AND2x2_ASAP7_75t_L g584 ( .A(n_443), .B(n_489), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_443), .B(n_488), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_443), .B(n_473), .Y(n_647) );
INVx1_ASAP7_75t_L g651 ( .A(n_443), .Y(n_651) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_460), .Y(n_443) );
INVx2_ASAP7_75t_L g568 ( .A(n_444), .Y(n_568) );
BUFx2_ASAP7_75t_L g595 ( .A(n_444), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
INVx5_ASAP7_75t_L g465 ( .A(n_447), .Y(n_465) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_SL g463 ( .A1(n_454), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_454), .A2(n_465), .B(n_545), .C(n_546), .Y(n_544) );
BUFx2_ASAP7_75t_L g492 ( .A(n_456), .Y(n_492) );
AND2x2_ASAP7_75t_L g535 ( .A(n_460), .B(n_489), .Y(n_535) );
INVx2_ASAP7_75t_L g551 ( .A(n_460), .Y(n_551) );
AND2x2_ASAP7_75t_L g560 ( .A(n_460), .B(n_488), .Y(n_560) );
AND2x2_ASAP7_75t_L g639 ( .A(n_460), .B(n_568), .Y(n_639) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_471), .Y(n_460) );
INVx2_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_501), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_473), .B(n_566), .Y(n_604) );
INVx1_ASAP7_75t_L g692 ( .A(n_473), .Y(n_692) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_488), .Y(n_473) );
AND2x2_ASAP7_75t_L g550 ( .A(n_474), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g564 ( .A(n_474), .B(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_474), .Y(n_593) );
OR2x2_ASAP7_75t_L g625 ( .A(n_474), .B(n_567), .Y(n_625) );
AND2x2_ASAP7_75t_L g633 ( .A(n_474), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g666 ( .A(n_474), .B(n_635), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_474), .B(n_535), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_474), .B(n_595), .Y(n_691) );
AND2x2_ASAP7_75t_L g697 ( .A(n_474), .B(n_584), .Y(n_697) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g557 ( .A(n_475), .Y(n_557) );
AND2x2_ASAP7_75t_L g587 ( .A(n_475), .B(n_567), .Y(n_587) );
AND2x2_ASAP7_75t_L g620 ( .A(n_475), .B(n_580), .Y(n_620) );
AND2x2_ASAP7_75t_L g640 ( .A(n_475), .B(n_489), .Y(n_640) );
AND2x2_ASAP7_75t_L g674 ( .A(n_475), .B(n_540), .Y(n_674) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_484), .C(n_485), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_482), .A2(n_485), .B(n_531), .C(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g580 ( .A(n_488), .B(n_551), .Y(n_580) );
AND2x2_ASAP7_75t_L g591 ( .A(n_488), .B(n_587), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_488), .B(n_567), .Y(n_630) );
INVx2_ASAP7_75t_L g645 ( .A(n_488), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_488), .B(n_579), .Y(n_668) );
AND2x2_ASAP7_75t_L g687 ( .A(n_488), .B(n_639), .Y(n_687) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_489), .Y(n_586) );
AND2x2_ASAP7_75t_L g594 ( .A(n_489), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g635 ( .A(n_489), .B(n_551), .Y(n_635) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
AOI21xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
AND2x2_ASAP7_75t_L g558 ( .A(n_503), .B(n_541), .Y(n_558) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_504), .B(n_515), .Y(n_538) );
OR2x2_ASAP7_75t_L g571 ( .A(n_504), .B(n_541), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_504), .B(n_541), .Y(n_576) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_540), .Y(n_603) );
AND2x2_ASAP7_75t_L g655 ( .A(n_504), .B(n_514), .Y(n_655) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_505), .B(n_525), .Y(n_563) );
AND2x2_ASAP7_75t_L g599 ( .A(n_505), .B(n_515), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_512), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_571), .Y(n_589) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_525), .Y(n_513) );
OAI322xp33_ASAP7_75t_L g554 ( .A1(n_514), .A2(n_555), .A3(n_559), .B1(n_561), .B2(n_564), .C1(n_569), .C2(n_577), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_514), .B(n_540), .Y(n_562) );
OR2x2_ASAP7_75t_L g572 ( .A(n_514), .B(n_526), .Y(n_572) );
AND2x2_ASAP7_75t_L g574 ( .A(n_514), .B(n_526), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_514), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_514), .B(n_541), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_514), .B(n_670), .Y(n_669) );
INVx5_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_515), .B(n_558), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_525), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g552 ( .A(n_525), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_525), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g614 ( .A(n_525), .B(n_541), .Y(n_614) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_525), .A2(n_643), .B(n_646), .C(n_658), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_525), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g680 ( .A(n_525), .B(n_655), .Y(n_680) );
INVx5_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g608 ( .A(n_526), .B(n_541), .Y(n_608) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
AND2x2_ASAP7_75t_L g657 ( .A(n_526), .B(n_655), .Y(n_657) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_526), .B(n_558), .Y(n_688) );
AND2x2_ASAP7_75t_L g695 ( .A(n_526), .B(n_654), .Y(n_695) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_550), .B2(n_552), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_535), .B(n_557), .Y(n_605) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g553 ( .A(n_538), .Y(n_553) );
OR2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g661 ( .A1(n_538), .A2(n_662), .B1(n_664), .B2(n_665), .C(n_667), .Y(n_661) );
INVx2_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
AND2x2_ASAP7_75t_L g573 ( .A(n_540), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g663 ( .A(n_540), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_540), .B(n_655), .Y(n_676) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVxp67_ASAP7_75t_L g618 ( .A(n_541), .Y(n_618) );
AND2x2_ASAP7_75t_L g654 ( .A(n_541), .B(n_655), .Y(n_654) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g656 ( .A(n_550), .B(n_595), .Y(n_656) );
AND2x2_ASAP7_75t_L g566 ( .A(n_551), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_551), .B(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g637 ( .A(n_553), .B(n_600), .Y(n_637) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g643 ( .A(n_556), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OR2x2_ASAP7_75t_L g629 ( .A(n_557), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g694 ( .A(n_557), .B(n_639), .Y(n_694) );
INVx2_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
NAND4xp25_ASAP7_75t_SL g690 ( .A(n_559), .B(n_691), .C(n_692), .D(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_560), .B(n_624), .Y(n_659) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_SL g696 ( .A(n_563), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_SL g658 ( .A1(n_564), .A2(n_627), .B(n_631), .C(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g653 ( .A(n_566), .B(n_645), .Y(n_653) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_567), .Y(n_579) );
INVx1_ASAP7_75t_L g634 ( .A(n_567), .Y(n_634) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_568), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B(n_573), .C(n_575), .Y(n_569) );
AND2x2_ASAP7_75t_L g590 ( .A(n_570), .B(n_574), .Y(n_590) );
OAI322xp33_ASAP7_75t_SL g628 ( .A1(n_570), .A2(n_629), .A3(n_631), .B1(n_632), .B2(n_636), .C1(n_637), .C2(n_638), .Y(n_628) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g650 ( .A(n_572), .B(n_576), .Y(n_650) );
INVx1_ASAP7_75t_L g631 ( .A(n_574), .Y(n_631) );
INVx1_ASAP7_75t_SL g649 ( .A(n_576), .Y(n_649) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_588), .B1(n_590), .B2(n_591), .C1(n_592), .C2(n_725), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .Y(n_582) );
OAI322xp33_ASAP7_75t_L g671 ( .A1(n_583), .A2(n_645), .A3(n_650), .B1(n_672), .B2(n_673), .C1(n_675), .C2(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_584), .A2(n_598), .B1(n_622), .B2(n_626), .C(n_628), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g601 ( .A1(n_589), .A2(n_602), .B1(n_604), .B2(n_605), .C1(n_606), .C2(n_609), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_591), .A2(n_598), .B1(n_668), .B2(n_669), .Y(n_667) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_601), .C(n_612), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_598), .A2(n_635), .B(n_678), .C(n_681), .Y(n_677) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g607 ( .A(n_599), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g670 ( .A(n_603), .Y(n_670) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_610), .B(n_635), .Y(n_664) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_619), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_613), .A2(n_682), .B1(n_683), .B2(n_684), .C(n_685), .Y(n_681) );
INVxp33_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_617), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_624), .B(n_635), .Y(n_675) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g686 ( .A(n_639), .B(n_645), .Y(n_686) );
AND4x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_660), .C(n_677), .D(n_689), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_648), .B1(n_650), .B2(n_651), .C(n_652), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g682 ( .A(n_653), .Y(n_682) );
INVx1_ASAP7_75t_SL g672 ( .A(n_657), .Y(n_672) );
NOR2xp33_ASAP7_75t_SL g660 ( .A(n_661), .B(n_671), .Y(n_660) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_673), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g706 ( .A(n_699), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx3_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
XNOR2xp5_ASAP7_75t_SL g713 ( .A(n_714), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
endmodule