module fake_jpeg_9864_n_15 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_15);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_15;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_9;

OAI22xp33_ASAP7_75t_SL g9 ( 
.A1(n_7),
.A2(n_0),
.B1(n_6),
.B2(n_3),
.Y(n_9)
);

OA22x2_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_4),
.B1(n_0),
.B2(n_5),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

HB1xp67_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_13),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_1),
.B(n_9),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_10),
.Y(n_15)
);


endmodule