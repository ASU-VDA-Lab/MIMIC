module fake_jpeg_20943_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_25),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_31),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_49),
.B1(n_37),
.B2(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_43),
.B1(n_26),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_22),
.B(n_21),
.C(n_32),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_31),
.B(n_25),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_85),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_20),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_27),
.CI(n_3),
.CON(n_122),
.SN(n_122)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_42),
.B1(n_32),
.B2(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_94),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_30),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_104),
.B1(n_62),
.B2(n_59),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_31),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_25),
.B1(n_27),
.B2(n_16),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_25),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_93),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_52),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_123),
.B(n_98),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_62),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_80),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_66),
.B(n_67),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_71),
.B1(n_77),
.B2(n_92),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_131),
.B(n_129),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_111),
.B1(n_115),
.B2(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_136),
.B1(n_147),
.B2(n_151),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_84),
.B1(n_75),
.B2(n_105),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_113),
.B1(n_129),
.B2(n_131),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_86),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_122),
.C(n_121),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_105),
.B(n_100),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_143),
.B(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_100),
.B(n_97),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_117),
.B1(n_113),
.B2(n_110),
.Y(n_147)
);

NAND2xp67_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_122),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_95),
.B1(n_106),
.B2(n_101),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_108),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_73),
.B1(n_74),
.B2(n_97),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_2),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_118),
.B1(n_124),
.B2(n_123),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

OAI221xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.C(n_142),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_112),
.B(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_160),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_134),
.B1(n_169),
.B2(n_144),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_112),
.B(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_157),
.C(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_108),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_182),
.B1(n_155),
.B2(n_167),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_164),
.B(n_168),
.Y(n_194)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_152),
.A3(n_148),
.B1(n_139),
.B2(n_149),
.C(n_138),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_166),
.A3(n_161),
.B1(n_120),
.B2(n_156),
.C1(n_158),
.C2(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_185),
.C(n_186),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_143),
.B1(n_149),
.B2(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_144),
.B1(n_149),
.B2(n_141),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_141),
.C(n_116),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_116),
.C(n_126),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_185),
.B(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_191),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_153),
.B(n_160),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_187),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_153),
.C(n_163),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_196),
.B(n_198),
.Y(n_202)
);

AOI31xp67_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_184),
.A3(n_182),
.B(n_173),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_161),
.B(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_14),
.A3(n_13),
.B1(n_109),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_5),
.C(n_6),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_5),
.C(n_8),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_191),
.C(n_190),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_192),
.C(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_218),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_201),
.Y(n_214)
);

OAI31xp33_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_8),
.A3(n_9),
.B(n_12),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_207),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_12),
.B(n_202),
.C(n_203),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_213),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_220),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_224),
.CI(n_221),
.CON(n_227),
.SN(n_227)
);


endmodule