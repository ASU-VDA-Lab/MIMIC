module real_jpeg_7261_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_0),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_0),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_0),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_0),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_0),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_119),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_0),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_1),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_1),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_1),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_2),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_2),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_2),
.Y(n_386)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_3),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_4),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_5),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_5),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_5),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_6),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_6),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_6),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_6),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_6),
.B(n_342),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_6),
.B(n_290),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_6),
.B(n_422),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_7),
.Y(n_413)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_9),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_9),
.Y(n_383)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_13),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_13),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_13),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_13),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_14),
.B(n_50),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_14),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_14),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_14),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_14),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_14),
.B(n_106),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_14),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_15),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_15),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_15),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_15),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_15),
.B(n_233),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_15),
.B(n_34),
.Y(n_398)
);

AND2x6_ASAP7_75t_SL g412 ( 
.A(n_15),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_16),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_16),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_16),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_16),
.B(n_48),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_16),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_16),
.B(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_16),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_16),
.B(n_383),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_17),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_17),
.B(n_99),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_17),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_17),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_290),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_17),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_17),
.B(n_226),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_17),
.B(n_233),
.Y(n_419)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_19),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_19),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_19),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_19),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_19),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_19),
.B(n_121),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_19),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_19),
.B(n_427),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_538),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_22),
.Y(n_539)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_46),
.B(n_81),
.C(n_537),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_51),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_27),
.B(n_51),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_44),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.C(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_29),
.A2(n_33),
.B1(n_45),
.B2(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_31),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_55),
.C(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_35),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_36),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_36),
.Y(n_309)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_36),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_77),
.C(n_79),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_52),
.B(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.C(n_69),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_62),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_55),
.A2(n_61),
.B1(n_73),
.B2(n_123),
.Y(n_127)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_58),
.Y(n_221)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.C(n_73),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_71),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_73),
.A2(n_117),
.B1(n_118),
.B2(n_123),
.Y(n_510)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_76),
.Y(n_236)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_76),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_134),
.B(n_536),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_131),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_83),
.B(n_131),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_128),
.C(n_129),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_84),
.A2(n_85),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_111),
.C(n_124),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_86),
.A2(n_87),
.B1(n_514),
.B2(n_516),
.Y(n_513)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_97),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_92),
.C(n_97),
.Y(n_128)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_107),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_98),
.B(n_505),
.Y(n_504)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_505)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_105),
.B(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_111),
.A2(n_124),
.B1(n_125),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_111),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_123),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_112),
.B(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_116),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_117),
.A2(n_118),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_118),
.B(n_209),
.C(n_213),
.Y(n_511)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_122),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_122),
.Y(n_371)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_128),
.B(n_129),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_530),
.B(n_535),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_498),
.B(n_527),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_310),
.B(n_497),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_264),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_138),
.B(n_264),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_206),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_139),
.B(n_207),
.C(n_239),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_180),
.C(n_190),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_140),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_153),
.C(n_167),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_141),
.B(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_148),
.C(n_152),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_146),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_153),
.A2(n_154),
.B1(n_167),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_163),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_155),
.B(n_163),
.Y(n_473)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_158),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_162),
.Y(n_366)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_162),
.Y(n_422)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_167),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_176),
.B2(n_177),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_171),
.B(n_176),
.C(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_175),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_175),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_176),
.A2(n_177),
.B1(n_213),
.B2(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_176),
.B(n_213),
.C(n_243),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_179),
.Y(n_333)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_179),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_190),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_184),
.A2(n_188),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_184),
.B(n_187),
.C(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_184),
.B(n_256),
.C(n_260),
.Y(n_506)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_199),
.C(n_203),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_191),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.C(n_197),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_192),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_197),
.Y(n_276)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_199),
.B(n_203),
.Y(n_296)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_202),
.Y(n_328)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_239),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_217),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_208),
.B(n_218),
.C(n_238),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_227),
.B1(n_237),
.B2(n_238),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_223),
.Y(n_252)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_228),
.B(n_232),
.C(n_234),
.Y(n_512)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_253),
.B2(n_254),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_240),
.B(n_255),
.C(n_262),
.Y(n_523)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.C(n_251),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_271),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_266),
.B(n_269),
.Y(n_493)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_271),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_294),
.C(n_297),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_273),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.C(n_284),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_274),
.A2(n_275),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_277),
.A2(n_278),
.B(n_280),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_277),
.B(n_284),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.C(n_292),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_441)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_292),
.B(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_382),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_294),
.A2(n_295),
.B1(n_297),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_297),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_306),
.C(n_307),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_299),
.B(n_475),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_300),
.B(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_302),
.Y(n_454)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_306),
.B(n_307),
.Y(n_475)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_491),
.B(n_496),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_478),
.B(n_490),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_460),
.B(n_477),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_434),
.B(n_459),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_403),
.B(n_433),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_374),
.B(n_402),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_355),
.B(n_373),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_335),
.B(n_354),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_329),
.B(n_334),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_326),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_323),
.Y(n_336)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_337),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_346),
.C(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_341),
.Y(n_361)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_349),
.B2(n_350),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_372),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_372),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_361),
.C(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_360),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_393),
.C(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_377),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_391),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_392),
.C(n_395),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_381),
.C(n_384),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_385),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_390),
.Y(n_414)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_399),
.C(n_400),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_398),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_432),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_432),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_416),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_415),
.C(n_458),
.Y(n_457)
);

XNOR2x1_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_414),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_412),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_448),
.C(n_449),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_416),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_423),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_425),
.C(n_430),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_420),
.C(n_421),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_430),
.B2(n_431),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_428),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_457),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_457),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_446),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_438),
.C(n_446),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_442),
.B2(n_443),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_469),
.C(n_470),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_451),
.C(n_456),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_455),
.B2(n_456),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_452),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_476),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_476),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_467),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_466),
.C(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_468),
.B(n_471),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_472),
.C(n_474),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_488),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_488),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_485),
.C(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_494),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_494),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_524),
.Y(n_498)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_499),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_518),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_518),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_507),
.B2(n_517),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_508),
.C(n_513),
.Y(n_534)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.C(n_506),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_520),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_506),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_513),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.C(n_512),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_522),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_512),
.Y(n_522)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_514),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.C(n_523),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g525 ( 
.A(n_519),
.B(n_521),
.CI(n_523),
.CON(n_525),
.SN(n_525)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_526),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_525),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);


endmodule