module fake_jpeg_13634_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_18),
.Y(n_22)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_14),
.B1(n_19),
.B2(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_17),
.B(n_12),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_23),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_21),
.B1(n_29),
.B2(n_31),
.Y(n_33)
);


endmodule