module fake_jpeg_23971_n_159 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_159);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_0),
.B(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_13),
.B2(n_23),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_51),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_13),
.B1(n_23),
.B2(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_18),
.B2(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_23),
.B1(n_13),
.B2(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_36),
.B1(n_27),
.B2(n_26),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AO21x2_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_16),
.B(n_3),
.Y(n_65)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_63),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_64),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_36),
.B1(n_18),
.B2(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_67),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_20),
.B1(n_24),
.B2(n_15),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_38),
.B(n_51),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_72),
.B(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_50),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_41),
.C(n_39),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_65),
.C(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_85),
.B1(n_59),
.B2(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_79),
.C(n_82),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_65),
.B(n_64),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_81),
.B(n_82),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_96),
.B(n_20),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_97),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_76),
.B1(n_83),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_112),
.B1(n_95),
.B2(n_92),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_82),
.C(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.C(n_114),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_19),
.B(n_3),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_2),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_120),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_90),
.B(n_98),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_94),
.C(n_89),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_129),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_131),
.C(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_114),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_113),
.B(n_4),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_124),
.B1(n_118),
.B2(n_117),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_131),
.C(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_119),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_139),
.B(n_141),
.Y(n_147)
);

OA21x2_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_122),
.B(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_142),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_130),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_132),
.C(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_147),
.B(n_8),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_153),
.B1(n_10),
.B2(n_11),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_10),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_156),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_151),
.A2(n_5),
.B1(n_6),
.B2(n_152),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_155),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_157),
.Y(n_159)
);


endmodule