module fake_jpeg_22650_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_17),
.B1(n_35),
.B2(n_20),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_65),
.B(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_29),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_17),
.B1(n_35),
.B2(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_17),
.B1(n_31),
.B2(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_29),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_67),
.B1(n_48),
.B2(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_78),
.B1(n_81),
.B2(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_42),
.B(n_39),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_60),
.B(n_69),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_40),
.B1(n_20),
.B2(n_35),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_40),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_1),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_31),
.B1(n_21),
.B2(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_86),
.B1(n_24),
.B2(n_30),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_22),
.B1(n_31),
.B2(n_36),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_90),
.B1(n_97),
.B2(n_24),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_31),
.B1(n_21),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_36),
.B1(n_40),
.B2(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_18),
.B(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_26),
.B1(n_18),
.B2(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_77),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_100),
.B(n_103),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_84),
.Y(n_133)
);

FAx1_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_71),
.CI(n_93),
.CON(n_103),
.SN(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_83),
.B1(n_78),
.B2(n_86),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_107),
.B1(n_97),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_62),
.B1(n_66),
.B2(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_115),
.Y(n_157)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_32),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_32),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_124),
.Y(n_147)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_127),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_45),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_18),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_32),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_79),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_137),
.B1(n_146),
.B2(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_72),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_101),
.B1(n_110),
.B2(n_122),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_76),
.B1(n_98),
.B2(n_85),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_80),
.C(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_148),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_98),
.B1(n_75),
.B2(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_105),
.B1(n_124),
.B2(n_116),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_100),
.B(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_50),
.B1(n_47),
.B2(n_75),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_95),
.C(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_73),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_29),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_167),
.B1(n_172),
.B2(n_176),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_180),
.B(n_183),
.Y(n_214)
);

XOR2x2_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_103),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_133),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_169),
.B(n_179),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_100),
.B(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_188),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_123),
.B1(n_104),
.B2(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_186),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_123),
.B1(n_126),
.B2(n_111),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_192),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_104),
.B(n_123),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_104),
.B1(n_126),
.B2(n_111),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_92),
.B1(n_119),
.B2(n_117),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_191),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_30),
.B(n_24),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_119),
.B1(n_112),
.B2(n_128),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_112),
.B1(n_128),
.B2(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_128),
.B(n_33),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_190),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_128),
.B(n_33),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_1),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_209),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_138),
.B1(n_149),
.B2(n_143),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_206),
.B1(n_176),
.B2(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_145),
.B1(n_134),
.B2(n_152),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_212),
.B1(n_19),
.B2(n_2),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_152),
.B1(n_142),
.B2(n_151),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_145),
.C(n_139),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_210),
.C(n_218),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_157),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_145),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_28),
.B(n_25),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_131),
.C(n_129),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_131),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_129),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_43),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_165),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_195),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_174),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_240),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_219),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_186),
.C(n_166),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_231),
.C(n_233),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_163),
.C(n_183),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_192),
.C(n_160),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_202),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_185),
.C(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_242),
.C(n_195),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_180),
.B1(n_188),
.B2(n_187),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_10),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_9),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_25),
.B1(n_19),
.B2(n_28),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_28),
.C(n_25),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_201),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_9),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_249),
.B(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_214),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_199),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_214),
.B(n_206),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_235),
.B(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_196),
.C(n_197),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_196),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_197),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_247),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_270),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_251),
.B1(n_239),
.B2(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_250),
.B1(n_227),
.B2(n_257),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_275),
.B(n_285),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_243),
.B(n_229),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_262),
.B1(n_233),
.B2(n_231),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_284),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_230),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_289),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_253),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_253),
.B(n_266),
.C(n_258),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_250),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_9),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_272),
.B(n_270),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_19),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_3),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_282),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_2),
.C(n_3),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_283),
.C(n_276),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_313),
.C(n_300),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_297),
.B(n_289),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_272),
.B1(n_273),
.B2(n_282),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_274),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_274),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_3),
.C(n_4),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_12),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_321),
.B1(n_8),
.B2(n_14),
.Y(n_327)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_323),
.C(n_324),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_307),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_308),
.A2(n_10),
.B(n_15),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_305),
.A3(n_303),
.B1(n_306),
.B2(n_313),
.C1(n_10),
.C2(n_12),
.Y(n_325)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_328),
.A3(n_331),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_330),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_327),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_14),
.C1(n_16),
.C2(n_323),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_319),
.B(n_5),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_4),
.B1(n_6),
.B2(n_329),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_325),
.Y(n_337)
);


endmodule