module fake_jpeg_25708_n_276 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_44),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_3),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_5),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_19),
.B(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_37),
.B1(n_38),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_63),
.B1(n_74),
.B2(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_28),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_78),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_32),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_70),
.A2(n_80),
.B(n_67),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_88),
.B(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_29),
.B1(n_23),
.B2(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_86),
.Y(n_96)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_55),
.B1(n_47),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_5),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_31),
.B1(n_25),
.B2(n_36),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_43),
.C(n_54),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_105),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_43),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_141)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_25),
.B1(n_20),
.B2(n_7),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_85),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_43),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_108),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_121),
.B1(n_89),
.B2(n_10),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_53),
.C(n_20),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_20),
.B1(n_48),
.B2(n_7),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_77),
.B1(n_64),
.B2(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_5),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_140),
.B(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_101),
.B1(n_123),
.B2(n_118),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_85),
.B1(n_64),
.B2(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_149),
.B1(n_123),
.B2(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_65),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_90),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_65),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_102),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_6),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_105),
.B1(n_96),
.B2(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_104),
.B1(n_122),
.B2(n_108),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_89),
.B1(n_9),
.B2(n_10),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_152),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_8),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_102),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_165),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_119),
.B1(n_110),
.B2(n_94),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_104),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_170),
.B1(n_132),
.B2(n_138),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_103),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_99),
.B1(n_97),
.B2(n_112),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_99),
.C(n_112),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_140),
.C(n_141),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_177),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_13),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_89),
.B1(n_14),
.B2(n_15),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_136),
.B1(n_127),
.B2(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_147),
.B1(n_134),
.B2(n_125),
.C(n_141),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_154),
.B1(n_130),
.B2(n_132),
.C(n_166),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_164),
.C(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_135),
.B(n_134),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_196),
.B(n_160),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_162),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_142),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_156),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_199),
.B1(n_193),
.B2(n_187),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_135),
.B(n_142),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_178),
.B(n_165),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_217),
.C(n_194),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_207),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_216),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_200),
.B1(n_198),
.B2(n_158),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_218),
.B1(n_220),
.B2(n_222),
.Y(n_235)
);

OAI322xp33_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_156),
.A3(n_180),
.B1(n_155),
.B2(n_169),
.C1(n_143),
.C2(n_150),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_130),
.C(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_155),
.C(n_175),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_154),
.B1(n_179),
.B2(n_166),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_208),
.B(n_222),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_203),
.B(n_210),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_217),
.B(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_182),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_196),
.B1(n_187),
.B2(n_181),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_209),
.B1(n_207),
.B2(n_211),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_205),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_248),
.C(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_234),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_206),
.B(n_215),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_182),
.B1(n_181),
.B2(n_192),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_245),
.Y(n_251)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_153),
.C(n_89),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_230),
.C(n_227),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_13),
.C(n_16),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_225),
.B1(n_229),
.B2(n_226),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_257),
.B1(n_238),
.B2(n_16),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_255),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_233),
.B1(n_223),
.B2(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_239),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_254),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_255),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_253),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_237),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_237),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_253),
.B(n_260),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_268),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_272),
.C(n_267),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_16),
.B(n_17),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_17),
.Y(n_276)
);


endmodule