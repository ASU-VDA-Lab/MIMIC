module fake_jpeg_1473_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.C(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_11),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_8),
.B1(n_24),
.B2(n_20),
.C(n_22),
.Y(n_30)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_4),
.B(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_9),
.B1(n_10),
.B2(n_7),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_33),
.B(n_31),
.Y(n_38)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_38),
.B1(n_30),
.B2(n_33),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_32),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_42),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_45),
.C(n_43),
.Y(n_47)
);


endmodule