module fake_jpeg_9444_n_80 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_35),
.B1(n_3),
.B2(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_54),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_20),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_13),
.B(n_15),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_70),
.C(n_66),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.C(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_65),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_59),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_62),
.C(n_47),
.Y(n_76)
);

NOR2xp67_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_62),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_47),
.B(n_52),
.Y(n_78)
);

OAI33xp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_68),
.A3(n_69),
.B1(n_50),
.B2(n_22),
.B3(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_21),
.Y(n_80)
);


endmodule