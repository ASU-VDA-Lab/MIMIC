module fake_aes_10955_n_666 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_666);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_627;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g83 ( .A(n_66), .Y(n_83) );
BUFx10_ASAP7_75t_L g84 ( .A(n_71), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_81), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_46), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_29), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_62), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_40), .Y(n_94) );
INVx1_ASAP7_75t_SL g95 ( .A(n_78), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_31), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_32), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_43), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_79), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_24), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_63), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_20), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_82), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_48), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
INVx4_ASAP7_75t_R g114 ( .A(n_8), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_34), .B(n_18), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_10), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_1), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_64), .Y(n_119) );
BUFx5_ASAP7_75t_L g120 ( .A(n_58), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_16), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_11), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_17), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_41), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_88), .B(n_37), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_91), .B(n_0), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_120), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_103), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_98), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_91), .B(n_3), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_98), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_90), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_93), .A2(n_39), .B(n_80), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_132), .A2(n_103), .B1(n_123), .B2(n_108), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_133), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_130), .B(n_99), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_127), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_141), .B(n_109), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_132), .A2(n_123), .B1(n_125), .B2(n_116), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_130), .B(n_100), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_127), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_148), .Y(n_168) );
NOR3xp33_ASAP7_75t_L g169 ( .A(n_143), .B(n_122), .C(n_121), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_151), .B(n_111), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_130), .B(n_99), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_141), .B(n_111), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_130), .A2(n_117), .B1(n_102), .B2(n_89), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_130), .B(n_102), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_151), .B(n_113), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_128), .B(n_113), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_129), .B(n_101), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_129), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_155), .A2(n_129), .B1(n_152), .B2(n_154), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_171), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_179), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_161), .B(n_129), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_168), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_168), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_165), .A2(n_152), .B1(n_154), .B2(n_128), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_187), .B(n_146), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_187), .B(n_131), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_186), .B(n_131), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
INVx6_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_182), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
OR2x2_ASAP7_75t_SL g213 ( .A(n_167), .B(n_146), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_166), .B(n_134), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_164), .B(n_146), .Y(n_216) );
AO22x1_ASAP7_75t_L g217 ( .A1(n_169), .A2(n_143), .B1(n_136), .B2(n_94), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_175), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_180), .B(n_142), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_166), .B(n_138), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_174), .B(n_138), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_163), .B(n_149), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_174), .B(n_134), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_184), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_174), .A2(n_139), .B1(n_140), .B2(n_145), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_184), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_159), .B(n_139), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_174), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_163), .B(n_149), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_203), .B(n_174), .Y(n_235) );
BUFx12f_ASAP7_75t_L g236 ( .A(n_199), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_210), .B(n_173), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_192), .Y(n_238) );
OAI221xp5_ASAP7_75t_L g239 ( .A1(n_202), .A2(n_140), .B1(n_145), .B2(n_185), .C(n_183), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_203), .B(n_184), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_194), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
BUFx12f_ASAP7_75t_L g245 ( .A(n_199), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_184), .B1(n_136), .B2(n_149), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_221), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_207), .B(n_172), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_205), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_225), .A2(n_185), .B(n_183), .Y(n_253) );
AOI21x1_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_178), .B(n_172), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_189), .Y(n_255) );
BUFx12f_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_150), .B(n_160), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_190), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_209), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_233), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_221), .Y(n_266) );
CKINVDCx11_ASAP7_75t_R g267 ( .A(n_200), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_222), .B(n_178), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_222), .B(n_153), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_224), .B(n_86), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_233), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_229), .Y(n_273) );
INVx4_ASAP7_75t_SL g274 ( .A(n_229), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_215), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
AOI21x1_ASAP7_75t_L g277 ( .A1(n_217), .A2(n_150), .B(n_158), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_197), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_256), .A2(n_218), .B1(n_224), .B2(n_197), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_247), .B(n_213), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_242), .Y(n_281) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_256), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_241), .Y(n_283) );
AOI221xp5_ASAP7_75t_SL g284 ( .A1(n_239), .A2(n_213), .B1(n_214), .B2(n_206), .C(n_204), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_256), .A2(n_218), .B1(n_216), .B2(n_226), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_242), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_239), .A2(n_193), .B1(n_228), .B2(n_231), .C(n_226), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_268), .A2(n_216), .B1(n_227), .B2(n_208), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_268), .B(n_216), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_260), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_241), .Y(n_293) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_249), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_278), .A2(n_231), .B1(n_136), .B2(n_211), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_278), .A2(n_231), .B1(n_220), .B2(n_208), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_255), .A2(n_83), .B1(n_118), .B2(n_105), .C(n_153), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_231), .B1(n_136), .B2(n_227), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_269), .B(n_208), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_244), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_249), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_271), .A2(n_230), .B(n_232), .C(n_223), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_269), .B(n_229), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_258), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_248), .A2(n_223), .B1(n_215), .B2(n_229), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_250), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_269), .B(n_232), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_250), .B(n_207), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_292), .B(n_248), .Y(n_317) );
AOI222xp33_ASAP7_75t_L g318 ( .A1(n_291), .A2(n_245), .B1(n_236), .B2(n_255), .C1(n_262), .C2(n_261), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_281), .A2(n_263), .B(n_276), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_288), .A2(n_252), .B1(n_243), .B2(n_238), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_291), .A2(n_252), .B1(n_243), .B2(n_238), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_254), .B(n_257), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_284), .A2(n_240), .B1(n_235), .B2(n_246), .C(n_261), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_238), .B(n_243), .C(n_240), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_280), .A2(n_262), .B1(n_264), .B2(n_265), .C(n_272), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_282), .A2(n_236), .B1(n_245), .B2(n_238), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_281), .A2(n_254), .B(n_257), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_282), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_280), .A2(n_236), .B1(n_245), .B2(n_235), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_293), .A2(n_237), .B1(n_264), .B2(n_272), .Y(n_331) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_299), .A2(n_246), .B(n_126), .C(n_243), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_279), .A2(n_237), .B1(n_136), .B2(n_265), .Y(n_333) );
AO31x2_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_253), .A3(n_276), .B(n_258), .Y(n_334) );
BUFx5_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_293), .A2(n_237), .B1(n_136), .B2(n_234), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_294), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_295), .A2(n_237), .B1(n_136), .B2(n_234), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
AO31x2_ASAP7_75t_L g340 ( .A1(n_286), .A2(n_253), .A3(n_276), .B(n_263), .Y(n_340) );
INVx5_ASAP7_75t_SL g341 ( .A(n_308), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_295), .A2(n_237), .B1(n_136), .B2(n_234), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_285), .A2(n_237), .B1(n_275), .B2(n_234), .C(n_124), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_303), .A2(n_136), .B1(n_147), .B2(n_135), .Y(n_344) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_296), .A2(n_277), .B(n_257), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_282), .A2(n_275), .B1(n_266), .B2(n_259), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_339), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_316), .Y(n_348) );
INVx5_ASAP7_75t_L g349 ( .A(n_341), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_289), .B1(n_303), .B2(n_282), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_331), .A2(n_305), .B(n_300), .Y(n_351) );
OAI21xp5_ASAP7_75t_SL g352 ( .A1(n_327), .A2(n_287), .B(n_308), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_330), .A2(n_307), .B1(n_297), .B2(n_300), .C(n_296), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_326), .Y(n_354) );
OAI211xp5_ASAP7_75t_SL g355 ( .A1(n_325), .A2(n_119), .B(n_106), .C(n_104), .Y(n_355) );
NAND2xp33_ASAP7_75t_R g356 ( .A(n_337), .B(n_287), .Y(n_356) );
INVx5_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_335), .B(n_286), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_335), .B(n_290), .Y(n_359) );
OAI31xp33_ASAP7_75t_L g360 ( .A1(n_343), .A2(n_292), .A3(n_287), .B(n_304), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_324), .A2(n_301), .B(n_306), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_317), .A2(n_294), .B1(n_292), .B2(n_308), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_335), .B(n_290), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_335), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_320), .A2(n_294), .B1(n_308), .B2(n_287), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
OA222x2_ASAP7_75t_L g369 ( .A1(n_335), .A2(n_290), .B1(n_298), .B2(n_302), .C1(n_312), .C2(n_309), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_323), .A2(n_314), .B1(n_308), .B2(n_298), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_321), .A2(n_298), .B1(n_302), .B2(n_309), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_319), .A2(n_302), .B(n_312), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_331), .B(n_312), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_277), .B(n_124), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_115), .B1(n_314), .B2(n_147), .C(n_135), .Y(n_375) );
AOI211x1_ASAP7_75t_SL g376 ( .A1(n_355), .A2(n_107), .B(n_112), .C(n_135), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_368), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g378 ( .A1(n_352), .A2(n_329), .B(n_308), .C(n_95), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_358), .B(n_335), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_358), .B(n_345), .Y(n_380) );
NAND3xp33_ASAP7_75t_L g381 ( .A(n_367), .B(n_333), .C(n_135), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_341), .B1(n_107), .B2(n_112), .C1(n_336), .C2(n_338), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_359), .B(n_334), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_356), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_348), .B(n_334), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_363), .A2(n_342), .B(n_338), .C(n_336), .Y(n_387) );
NOR2xp33_ASAP7_75t_SL g388 ( .A(n_349), .B(n_313), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_350), .A2(n_342), .B(n_344), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
AOI31xp33_ASAP7_75t_L g392 ( .A1(n_350), .A2(n_346), .A3(n_315), .B(n_344), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_351), .A2(n_135), .B(n_144), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_374), .A2(n_361), .B(n_328), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_364), .B(n_334), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_349), .B(n_313), .Y(n_396) );
OAI33xp33_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_153), .A3(n_114), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_360), .A2(n_96), .B1(n_135), .B2(n_144), .C(n_147), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_364), .B(n_340), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_375), .B(n_144), .C(n_135), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_351), .A2(n_147), .B1(n_144), .B2(n_188), .C(n_177), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_370), .A2(n_263), .B1(n_270), .B2(n_5), .C(n_6), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_347), .B(n_340), .Y(n_408) );
AOI31xp33_ASAP7_75t_L g409 ( .A1(n_369), .A2(n_315), .A3(n_311), .B(n_313), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_371), .A2(n_310), .B(n_313), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_383), .B(n_373), .Y(n_411) );
AOI21x1_ASAP7_75t_L g412 ( .A1(n_381), .A2(n_372), .B(n_369), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_401), .B(n_373), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_378), .B(n_357), .C(n_349), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_383), .B(n_373), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_401), .B(n_374), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_395), .B(n_374), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_366), .B1(n_357), .B2(n_349), .C(n_362), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_385), .B(n_3), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_395), .B(n_362), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_357), .B1(n_349), .B2(n_120), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_403), .B(n_362), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_400), .B(n_362), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_400), .B(n_362), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_380), .B(n_120), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_380), .B(n_120), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_384), .B(n_120), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_403), .B(n_340), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_379), .B(n_340), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_406), .B(n_357), .C(n_144), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_382), .B(n_357), .C(n_144), .Y(n_434) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_409), .B(n_310), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_379), .B(n_144), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_386), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_408), .B(n_310), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_390), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_407), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_408), .B(n_310), .Y(n_442) );
BUFx12f_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_390), .B(n_147), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_147), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_398), .B(n_147), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_377), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_150), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_391), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_409), .B(n_310), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_391), .B(n_150), .Y(n_452) );
NOR3xp33_ASAP7_75t_SL g453 ( .A(n_387), .B(n_4), .C(n_7), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_150), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_394), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_392), .B(n_4), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_394), .B(n_9), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_394), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_410), .B(n_9), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_457), .B(n_397), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_420), .B(n_393), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_456), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_427), .B(n_381), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_420), .B(n_393), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_443), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_443), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_457), .A2(n_399), .B1(n_388), .B2(n_402), .C(n_376), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_428), .B(n_376), .Y(n_473) );
AND3x2_ASAP7_75t_L g474 ( .A(n_419), .B(n_388), .C(n_396), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_428), .B(n_396), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_430), .B(n_10), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_440), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_424), .B(n_404), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_424), .B(n_11), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_418), .A2(n_402), .B1(n_310), .B2(n_266), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_426), .B(n_12), .Y(n_481) );
AOI21xp5_ASAP7_75t_SL g482 ( .A1(n_418), .A2(n_315), .B(n_273), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_411), .B(n_12), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_435), .B(n_250), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_430), .B(n_13), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_414), .B(n_266), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_443), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_437), .B(n_14), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_436), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_413), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_426), .B(n_15), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_411), .B(n_15), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_423), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_415), .B(n_16), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_413), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_417), .B(n_18), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_425), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_417), .B(n_19), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_438), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_415), .B(n_19), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_431), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_432), .B(n_20), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_458), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_422), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_432), .B(n_21), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g513 ( .A1(n_450), .A2(n_188), .B(n_170), .C(n_176), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_422), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_446), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_416), .B(n_21), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_416), .B(n_22), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_446), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_438), .B(n_22), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_449), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_467), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_468), .A2(n_435), .B1(n_434), .B2(n_433), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_468), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_490), .B(n_434), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_492), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_463), .B(n_470), .Y(n_526) );
NOR2xp67_ASAP7_75t_L g527 ( .A(n_468), .B(n_433), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_471), .B(n_438), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_472), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_495), .B(n_449), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_461), .B(n_460), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_500), .B(n_451), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_461), .B(n_460), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_465), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_504), .B(n_451), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
NAND2xp33_ASAP7_75t_SL g539 ( .A(n_468), .B(n_453), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_487), .B(n_438), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_465), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_482), .B(n_485), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_484), .B(n_421), .Y(n_543) );
AOI321xp33_ASAP7_75t_L g544 ( .A1(n_497), .A2(n_421), .A3(n_455), .B1(n_445), .B2(n_459), .C(n_447), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_482), .B(n_445), .Y(n_545) );
NAND2x1_ASAP7_75t_L g546 ( .A(n_489), .B(n_444), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_509), .A2(n_453), .B1(n_455), .B2(n_459), .C(n_447), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_507), .Y(n_548) );
NAND3xp33_ASAP7_75t_SL g549 ( .A(n_513), .B(n_444), .C(n_429), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_508), .B(n_429), .Y(n_550) );
XNOR2xp5_ASAP7_75t_L g551 ( .A(n_497), .B(n_442), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_499), .A2(n_442), .B1(n_439), .B2(n_425), .Y(n_552) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_485), .B(n_425), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_508), .B(n_439), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_505), .B(n_442), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_499), .A2(n_412), .B(n_459), .C(n_448), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g558 ( .A1(n_510), .A2(n_442), .B(n_448), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_512), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_515), .B(n_412), .Y(n_560) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_474), .B(n_454), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_483), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_493), .B(n_454), .C(n_452), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
XNOR2xp5_ASAP7_75t_L g565 ( .A(n_479), .B(n_452), .Y(n_565) );
XNOR2x2_ASAP7_75t_L g566 ( .A(n_479), .B(n_251), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_481), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_518), .B(n_160), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_475), .A2(n_266), .B1(n_259), .B2(n_250), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_481), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_514), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_506), .B(n_23), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_494), .B(n_26), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_501), .B(n_27), .Y(n_574) );
OAI21xp33_ASAP7_75t_L g575 ( .A1(n_496), .A2(n_158), .B(n_188), .Y(n_575) );
XNOR2x1_ASAP7_75t_L g576 ( .A(n_496), .B(n_519), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_483), .B(n_188), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_498), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_503), .A2(n_170), .B1(n_176), .B2(n_188), .C(n_177), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_516), .B(n_177), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_517), .B(n_177), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_502), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_502), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_478), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_478), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_462), .B(n_28), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_469), .A2(n_170), .B1(n_176), .B2(n_177), .Y(n_588) );
AOI311xp33_ASAP7_75t_L g589 ( .A1(n_476), .A2(n_30), .A3(n_33), .B(n_35), .C(n_38), .Y(n_589) );
AOI31xp33_ASAP7_75t_L g590 ( .A1(n_480), .A2(n_270), .A3(n_274), .B(n_47), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_486), .B(n_44), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_473), .B(n_45), .Y(n_592) );
OAI32xp33_ASAP7_75t_L g593 ( .A1(n_464), .A2(n_266), .A3(n_259), .B1(n_273), .B2(n_270), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_462), .B(n_49), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_466), .Y(n_595) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_466), .A2(n_250), .B(n_259), .C(n_176), .Y(n_596) );
XNOR2x1_ASAP7_75t_L g597 ( .A(n_480), .B(n_50), .Y(n_597) );
AND2x4_ASAP7_75t_SL g598 ( .A(n_468), .B(n_176), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_504), .B(n_170), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_461), .A2(n_170), .B1(n_274), .B2(n_54), .Y(n_601) );
NOR2xp33_ASAP7_75t_R g602 ( .A(n_468), .B(n_51), .Y(n_602) );
OA22x2_ASAP7_75t_L g603 ( .A1(n_490), .A2(n_53), .B1(n_55), .B2(n_56), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g604 ( .A1(n_482), .A2(n_207), .B(n_60), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_463), .B(n_57), .Y(n_605) );
NAND3xp33_ASAP7_75t_SL g606 ( .A(n_490), .B(n_65), .C(n_69), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g607 ( .A1(n_482), .A2(n_207), .B(n_74), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_461), .A2(n_274), .B1(n_75), .B2(n_76), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_463), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_463), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_522), .A2(n_557), .B(n_531), .C(n_533), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_539), .B(n_547), .C(n_522), .Y(n_612) );
OAI22xp33_ASAP7_75t_SL g613 ( .A1(n_521), .A2(n_542), .B1(n_567), .B2(n_546), .Y(n_613) );
NOR2xp33_ASAP7_75t_R g614 ( .A(n_606), .B(n_523), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_586), .B(n_585), .Y(n_615) );
AOI22x1_ASAP7_75t_L g616 ( .A1(n_607), .A2(n_604), .B1(n_544), .B2(n_610), .Y(n_616) );
BUFx2_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
AND4x1_ASAP7_75t_L g618 ( .A(n_589), .B(n_604), .C(n_607), .D(n_547), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_524), .A2(n_567), .B1(n_559), .B2(n_543), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_527), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_541), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_545), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_609), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_576), .A2(n_570), .B1(n_551), .B2(n_565), .Y(n_624) );
OR3x1_ASAP7_75t_L g625 ( .A(n_549), .B(n_558), .C(n_594), .Y(n_625) );
NAND4xp75_ASAP7_75t_L g626 ( .A(n_587), .B(n_526), .C(n_605), .D(n_560), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_603), .A2(n_590), .B(n_549), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_561), .B(n_603), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_559), .A2(n_557), .B1(n_595), .B2(n_571), .C(n_564), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_548), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_563), .A2(n_525), .B1(n_599), .B2(n_550), .C(n_554), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_575), .A2(n_597), .B1(n_563), .B2(n_588), .C(n_552), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_624), .B(n_538), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_623), .Y(n_635) );
OAI321xp33_ASAP7_75t_L g636 ( .A1(n_624), .A2(n_608), .A3(n_601), .B1(n_592), .B2(n_574), .C(n_572), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_612), .A2(n_596), .B(n_591), .C(n_569), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_627), .A2(n_553), .B(n_580), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_631), .B(n_529), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_613), .A2(n_593), .B(n_540), .C(n_528), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_611), .A2(n_535), .B1(n_536), .B2(n_530), .C(n_532), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_573), .B(n_582), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_625), .A2(n_556), .B1(n_537), .B2(n_579), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_632), .B(n_581), .C(n_600), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_616), .A2(n_600), .B(n_566), .C(n_568), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_621), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_635), .Y(n_647) );
AND3x2_ASAP7_75t_L g648 ( .A(n_634), .B(n_620), .C(n_622), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_646), .Y(n_649) );
OAI222xp33_ASAP7_75t_L g650 ( .A1(n_643), .A2(n_619), .B1(n_632), .B2(n_617), .C1(n_615), .C2(n_630), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_644), .B(n_629), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_641), .A2(n_645), .B1(n_638), .B2(n_642), .C(n_637), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_641), .B(n_618), .C(n_614), .Y(n_653) );
NOR4xp25_ASAP7_75t_L g654 ( .A(n_653), .B(n_639), .C(n_636), .D(n_633), .Y(n_654) );
OA22x2_ASAP7_75t_L g655 ( .A1(n_648), .A2(n_615), .B1(n_640), .B2(n_626), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_652), .B(n_577), .C(n_579), .Y(n_656) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_651), .B(n_598), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_654), .B(n_647), .C(n_650), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_656), .A2(n_647), .B(n_649), .C(n_577), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_657), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_660), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_658), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_662), .A2(n_655), .B1(n_659), .B2(n_541), .C(n_584), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g665 ( .A(n_663), .B(n_583), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_664), .B1(n_578), .B2(n_562), .C(n_534), .Y(n_666) );
endmodule