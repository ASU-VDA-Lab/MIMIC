module real_jpeg_27528_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_73;
wire n_65;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_58;
wire n_49;
wire n_31;
wire n_52;
wire n_76;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_75;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_11;
wire n_14;
wire n_71;
wire n_45;
wire n_25;
wire n_51;
wire n_61;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_39;
wire n_36;
wire n_40;
wire n_70;
wire n_74;
wire n_41;
wire n_32;
wire n_20;
wire n_48;
wire n_27;
wire n_19;
wire n_26;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_0),
.A2(n_15),
.B1(n_20),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_0),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_31),
.B(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_31),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_15),
.B1(n_20),
.B2(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_15),
.B1(n_20),
.B2(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g40 ( 
.A1(n_5),
.A2(n_20),
.A3(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_15),
.B1(n_20),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_58),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_44),
.B(n_57),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_27),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_13),
.B(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_13)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_19),
.A2(n_26),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_47),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_25),
.Y(n_75)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_40),
.B2(n_43),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_28),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B(n_56),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_76),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_62),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_72),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);


endmodule