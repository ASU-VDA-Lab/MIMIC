module fake_netlist_5_346_n_524 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_524);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_524;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_483;
wire n_467;
wire n_423;
wire n_501;
wire n_245;
wire n_284;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_373;
wire n_307;
wire n_439;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_492;
wire n_171;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_297;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_223;
wire n_392;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_344;
wire n_287;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_258;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_463;
wire n_488;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_404;
wire n_233;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_426;
wire n_520;
wire n_409;
wire n_500;
wire n_300;
wire n_435;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_13),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_25),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_92),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_24),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_23),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_99),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_60),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_44),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_78),
.B(n_108),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_54),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVxp33_ASAP7_75t_SL g213 ( 
.A(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_56),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_45),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_83),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_39),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_85),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_58),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_50),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_64),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_97),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_125),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_61),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_148),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_66),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_43),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_95),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_47),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_70),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_130),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_79),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_126),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_17),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_65),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_90),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g256 ( 
.A(n_42),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_93),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_123),
.Y(n_259)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_67),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_142),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_133),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_105),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_122),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_89),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_131),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_151),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_26),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_10),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_96),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_106),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_118),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_100),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_155),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_145),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_129),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_124),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_55),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_141),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_115),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_186),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_164),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_165),
.Y(n_292)
);

CKINVDCx8_ASAP7_75t_R g293 ( 
.A(n_176),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_167),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_234),
.B(n_0),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_194),
.B(n_0),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_179),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_201),
.B(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_238),
.B(n_4),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_179),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_6),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_168),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_169),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_170),
.B(n_11),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_163),
.A2(n_14),
.B(n_15),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_173),
.B(n_16),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_172),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_174),
.B(n_19),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_177),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_188),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_203),
.B(n_20),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_183),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_188),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_162),
.B(n_21),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_R g322 ( 
.A(n_184),
.B(n_22),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_185),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_189),
.B(n_29),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_166),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_187),
.B(n_34),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_191),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_171),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_192),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_193),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_271),
.B(n_37),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_195),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_204),
.B(n_40),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_180),
.B(n_41),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_199),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_273),
.B(n_46),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_181),
.B(n_48),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_200),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_205),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_220),
.B(n_49),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_272),
.B(n_276),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_206),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_208),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_52),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_178),
.B(n_57),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_211),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_331),
.A2(n_260),
.B1(n_190),
.B2(n_213),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_256),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_347),
.A2(n_270),
.B1(n_265),
.B2(n_226),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_283),
.B1(n_281),
.B2(n_268),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_293),
.B(n_197),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_302),
.B(n_259),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_212),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_298),
.B(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_297),
.B(n_214),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_216),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_313),
.B(n_215),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_219),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_217),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_223),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_218),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_294),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_230),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_229),
.B(n_247),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_224),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_225),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_248),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_348),
.B(n_236),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_255),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_317),
.B(n_320),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_324),
.B(n_243),
.Y(n_380)
);

OR2x6_ASAP7_75t_L g381 ( 
.A(n_289),
.B(n_237),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_291),
.B(n_288),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_280),
.C(n_267),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g385 ( 
.A(n_325),
.B(n_250),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_252),
.B1(n_221),
.B2(n_240),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_351),
.A2(n_210),
.B1(n_343),
.B2(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

AO22x1_ASAP7_75t_L g390 ( 
.A1(n_371),
.A2(n_321),
.B1(n_318),
.B2(n_222),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_321),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_306),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_364),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_307),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

AO22x1_ASAP7_75t_L g400 ( 
.A1(n_367),
.A2(n_321),
.B1(n_254),
.B2(n_258),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_311),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_349),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_362),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_337),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_315),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_319),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_314),
.Y(n_414)
);

AO221x1_ASAP7_75t_L g415 ( 
.A1(n_372),
.A2(n_263),
.B1(n_249),
.B2(n_246),
.C(n_253),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_396),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_393),
.A2(n_353),
.B1(n_354),
.B2(n_387),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_388),
.A2(n_363),
.B1(n_310),
.B2(n_335),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_397),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_398),
.B(n_274),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_401),
.A2(n_373),
.B1(n_375),
.B2(n_374),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_355),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_394),
.B(n_368),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_384),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_350),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_341),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_333),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_235),
.B1(n_242),
.B2(n_241),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_414),
.A2(n_232),
.B1(n_233),
.B2(n_231),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_392),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_385),
.Y(n_437)
);

CKINVDCx11_ASAP7_75t_R g438 ( 
.A(n_409),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_403),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_413),
.B1(n_402),
.B2(n_257),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_431),
.Y(n_441)
);

BUFx2_ASAP7_75t_R g442 ( 
.A(n_425),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_400),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_395),
.Y(n_444)
);

CKINVDCx6p67_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_422),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_432),
.Y(n_447)
);

INVx4_ASAP7_75t_SL g448 ( 
.A(n_426),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_309),
.B(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_390),
.B(n_228),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_415),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_346),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_416),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_437),
.Y(n_456)
);

AOI221xp5_ASAP7_75t_L g457 ( 
.A1(n_440),
.A2(n_418),
.B1(n_434),
.B2(n_435),
.C(n_423),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_455),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_428),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_449),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_428),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_438),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_467),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_459),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_453),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_462),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_466),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_465),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_452),
.B(n_443),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_443),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

AOI221xp5_ASAP7_75t_L g483 ( 
.A1(n_469),
.A2(n_327),
.B1(n_345),
.B2(n_342),
.C(n_279),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_460),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_287),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_478),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_322),
.B1(n_286),
.B2(n_285),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_262),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_266),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_470),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_486),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_474),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_479),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_485),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_492),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_490),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_493),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_484),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_481),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_489),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_483),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_503),
.A2(n_482),
.B(n_269),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_261),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

AO21x1_ASAP7_75t_L g508 ( 
.A1(n_506),
.A2(n_502),
.B(n_500),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_497),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_282),
.B(n_275),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_507),
.B(n_482),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_251),
.C(n_227),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_508),
.Y(n_513)
);

AOI21xp33_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_284),
.B(n_244),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_511),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_76),
.C(n_80),
.Y(n_516)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_513),
.C(n_84),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_82),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_518),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_517),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_101),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

O2A1O1Ixp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_521),
.B(n_520),
.C(n_112),
.Y(n_524)
);


endmodule