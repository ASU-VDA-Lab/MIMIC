module fake_ariane_2132_n_1618 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1618);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1618;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_77),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_65),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_43),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_29),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_30),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_53),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_57),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_79),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_119),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_49),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_98),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_90),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_67),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_78),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_49),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_16),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_10),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_34),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_10),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_45),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_5),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_57),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_103),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_123),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_2),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_81),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_96),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_74),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_40),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_104),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_73),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_47),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_28),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_45),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_18),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_72),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_129),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_4),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_33),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_93),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_89),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_46),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_34),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_18),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_76),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_20),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_134),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_1),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_58),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_31),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_80),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_136),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_44),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_35),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_110),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_108),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_20),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_41),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_91),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_19),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_50),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_130),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_92),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_82),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_29),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_102),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_118),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_86),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_150),
.B(n_3),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_177),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_154),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_152),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_186),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_228),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_156),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_159),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_3),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_173),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_151),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_194),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_207),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_208),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_6),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_210),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_145),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_151),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_163),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_206),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_176),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_227),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_236),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_236),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_179),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_182),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_236),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_232),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_236),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_214),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_191),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_214),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_241),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_180),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_248),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_197),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_201),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_205),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_205),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_257),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_218),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_219),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_149),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_158),
.B(n_7),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_264),
.B(n_8),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_289),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_289),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_315),
.A2(n_168),
.B(n_162),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_184),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_313),
.A2(n_237),
.B1(n_268),
.B2(n_243),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_315),
.B(n_160),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_295),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_294),
.B(n_169),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_296),
.B(n_283),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_264),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_298),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_309),
.B(n_172),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_174),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_310),
.B(n_178),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_157),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_316),
.B(n_318),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_183),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_305),
.B(n_189),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_303),
.B(n_276),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_319),
.B(n_195),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_211),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_212),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_359),
.B(n_184),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_286),
.B(n_276),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_350),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_400),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_410),
.A2(n_353),
.B1(n_324),
.B2(n_357),
.Y(n_433)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_423),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_419),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_410),
.B(n_329),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_394),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_378),
.B(n_330),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_366),
.B(n_301),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_384),
.B(n_333),
.Y(n_444)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_358),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_371),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_387),
.B(n_306),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_336),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

AND3x2_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_343),
.C(n_317),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_385),
.B(n_344),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_385),
.B(n_345),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_377),
.Y(n_464)
);

AO22x2_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_306),
.B1(n_200),
.B2(n_261),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_384),
.B(n_354),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_366),
.B(n_355),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_403),
.A2(n_356),
.B1(n_300),
.B2(n_153),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_360),
.B1(n_193),
.B2(n_185),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_413),
.B(n_302),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_387),
.B(n_358),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_422),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_423),
.B(n_304),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_407),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_377),
.B(n_311),
.Y(n_485)
);

INVx8_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_420),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_413),
.A2(n_267),
.B1(n_244),
.B2(n_234),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_414),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_424),
.B(n_314),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_407),
.B(n_165),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_424),
.B(n_144),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_407),
.A2(n_199),
.B1(n_170),
.B2(n_282),
.Y(n_503)
);

NOR2x1p5_ASAP7_75t_L g504 ( 
.A(n_429),
.B(n_163),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_337),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_417),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_390),
.B(n_288),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_390),
.A2(n_164),
.B1(n_254),
.B2(n_255),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_423),
.B(n_144),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_363),
.B(n_146),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_363),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_423),
.B(n_146),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_394),
.B(n_337),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_412),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_394),
.B(n_339),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_394),
.B(n_147),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_394),
.B(n_339),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_364),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_364),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_412),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_365),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_402),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_365),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_412),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_416),
.B(n_340),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_340),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_369),
.Y(n_531)
);

OAI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_418),
.A2(n_164),
.B1(n_255),
.B2(n_272),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_367),
.B(n_293),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_402),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_342),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_389),
.B(n_147),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_367),
.Y(n_538)
);

NOR2x1p5_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_254),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_370),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_389),
.B(n_148),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_426),
.B(n_181),
.C(n_175),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_412),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_370),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_369),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_342),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_412),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_374),
.B(n_148),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_374),
.B(n_307),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_379),
.B(n_155),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_402),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_379),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_380),
.B(n_272),
.C(n_265),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_412),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_380),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_381),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_428),
.B(n_347),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_381),
.Y(n_560)
);

NOR3xp33_ASAP7_75t_L g561 ( 
.A(n_392),
.B(n_274),
.C(n_275),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_386),
.B(n_308),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_386),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_402),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_388),
.B(n_155),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_388),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_368),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_368),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_368),
.B(n_347),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_392),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_369),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_391),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_448),
.B(n_508),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_441),
.B(n_396),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_448),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_396),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_463),
.A2(n_401),
.B1(n_406),
.B2(n_404),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_571),
.B(n_398),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_540),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_431),
.B(n_398),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_454),
.B(n_404),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_480),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_431),
.B(n_406),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_457),
.B(n_401),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_436),
.B(n_439),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_485),
.B(n_312),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_436),
.B(n_369),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_472),
.B(n_369),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_522),
.B(n_369),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_463),
.A2(n_161),
.B1(n_166),
.B2(n_284),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_439),
.B(n_480),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_522),
.B(n_369),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_554),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_480),
.B(n_373),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_529),
.B(n_373),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_529),
.B(n_373),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_529),
.B(n_530),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_522),
.B(n_435),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_472),
.B(n_373),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_529),
.B(n_373),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_530),
.B(n_373),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_530),
.B(n_373),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_530),
.B(n_375),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_501),
.B(n_375),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_554),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_501),
.B(n_375),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_533),
.B(n_320),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_551),
.B(n_323),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_494),
.B(n_280),
.C(n_223),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_562),
.B(n_326),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_435),
.B(n_375),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_484),
.B(n_427),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_511),
.B(n_375),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_472),
.B(n_375),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_L g620 ( 
.A(n_478),
.B(n_213),
.C(n_220),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_484),
.B(n_375),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_438),
.A2(n_161),
.B1(n_284),
.B2(n_278),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_518),
.B(n_427),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_556),
.B(n_427),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_518),
.B(n_427),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_444),
.B(n_427),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_467),
.B(n_427),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_537),
.B(n_226),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_488),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_488),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_556),
.B(n_166),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_521),
.B(n_167),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_256),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_482),
.B(n_256),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_442),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_487),
.B(n_258),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_504),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_493),
.Y(n_638)
);

AND2x6_ASAP7_75t_SL g639 ( 
.A(n_516),
.B(n_235),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_516),
.B(n_273),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_263),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_430),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_493),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_541),
.B(n_238),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_443),
.B(n_332),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_498),
.B(n_263),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_445),
.B(n_250),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_445),
.B(n_266),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_248),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_433),
.B(n_277),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_445),
.B(n_251),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_280),
.C(n_278),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_495),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_485),
.B(n_279),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_531),
.B(n_277),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_539),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_442),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_531),
.B(n_216),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_449),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_276),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_470),
.B(n_524),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_449),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_496),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_452),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_445),
.B(n_231),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_516),
.B(n_408),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_519),
.B(n_240),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_532),
.B(n_245),
.C(n_249),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_452),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_440),
.B(n_408),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_506),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_547),
.B(n_262),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_507),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_477),
.B(n_415),
.C(n_421),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_483),
.B(n_171),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_497),
.B(n_408),
.Y(n_679)
);

INVx8_ASAP7_75t_L g680 ( 
.A(n_505),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_505),
.B(n_411),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_415),
.C(n_421),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_499),
.B(n_13),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_505),
.B(n_15),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_453),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_555),
.B(n_550),
.C(n_513),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_507),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_453),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_547),
.B(n_415),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_455),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_505),
.B(n_16),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_547),
.B(n_415),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_486),
.A2(n_421),
.B(n_411),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_455),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_514),
.A2(n_573),
.B1(n_538),
.B2(n_527),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_446),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_514),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_489),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_547),
.B(n_415),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_489),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_440),
.B(n_411),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_535),
.B(n_459),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_465),
.B(n_383),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_440),
.B(n_415),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_511),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_490),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_490),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_535),
.B(n_383),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_492),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_492),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_459),
.B(n_17),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_468),
.B(n_415),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_471),
.B(n_383),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_456),
.B(n_397),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_469),
.B(n_180),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_502),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_502),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_552),
.B(n_229),
.C(n_187),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_503),
.B(n_397),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_437),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_437),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_523),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_469),
.B(n_180),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_491),
.B(n_190),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_491),
.B(n_233),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_523),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_491),
.B(n_180),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_184),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_548),
.B(n_397),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_465),
.A2(n_376),
.B1(n_399),
.B2(n_184),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_447),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_525),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_525),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_574),
.A2(n_465),
.B1(n_500),
.B2(n_471),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_587),
.B(n_500),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_583),
.A2(n_486),
.B(n_569),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_585),
.B(n_548),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_645),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_575),
.A2(n_584),
.B(n_586),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_629),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_L g742 ( 
.A1(n_575),
.A2(n_568),
.B(n_569),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_588),
.A2(n_566),
.B(n_546),
.C(n_563),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_630),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_680),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_672),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_584),
.A2(n_557),
.B1(n_558),
.B2(n_567),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_663),
.B(n_517),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_638),
.A2(n_557),
.B1(n_558),
.B2(n_567),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_663),
.B(n_517),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_576),
.A2(n_528),
.B1(n_545),
.B2(n_549),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_621),
.A2(n_486),
.B(n_568),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_577),
.B(n_560),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_611),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_643),
.A2(n_560),
.B1(n_563),
.B2(n_475),
.Y(n_755)
);

AO21x1_ASAP7_75t_L g756 ( 
.A1(n_678),
.A2(n_447),
.B(n_450),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_612),
.Y(n_757)
);

BUFx4f_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_642),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_590),
.A2(n_486),
.B(n_432),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_653),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_595),
.B(n_579),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_673),
.A2(n_432),
.B(n_451),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_640),
.B(n_548),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_647),
.A2(n_528),
.B1(n_545),
.B2(n_549),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_703),
.B(n_601),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_654),
.B(n_464),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_655),
.Y(n_768)
);

OAI21xp33_ASAP7_75t_L g769 ( 
.A1(n_628),
.A2(n_460),
.B(n_458),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_432),
.B(n_451),
.Y(n_770)
);

NAND2x1_ASAP7_75t_L g771 ( 
.A(n_618),
.B(n_553),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_705),
.A2(n_451),
.B(n_512),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_705),
.A2(n_515),
.B(n_520),
.Y(n_773)
);

NOR2x1_ASAP7_75t_R g774 ( 
.A(n_615),
.B(n_559),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_661),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_713),
.A2(n_520),
.B(n_526),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_649),
.B(n_458),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_716),
.A2(n_473),
.B(n_543),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_665),
.A2(n_510),
.B1(n_553),
.B2(n_564),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_667),
.B(n_670),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_642),
.B(n_559),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_685),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_668),
.A2(n_553),
.B1(n_564),
.B2(n_462),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_680),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_628),
.A2(n_462),
.B(n_479),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_713),
.A2(n_526),
.B(n_534),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_647),
.B(n_461),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_592),
.A2(n_534),
.B(n_536),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_580),
.B(n_564),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_724),
.A2(n_728),
.B(n_598),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_581),
.B(n_565),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_623),
.A2(n_479),
.B(n_466),
.C(n_476),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_625),
.A2(n_476),
.B(n_466),
.C(n_570),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_592),
.A2(n_543),
.B(n_536),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_580),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_684),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_688),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_683),
.A2(n_572),
.B(n_570),
.C(n_464),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_714),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_676),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_670),
.B(n_570),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_580),
.B(n_572),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_580),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_596),
.A2(n_434),
.B(n_202),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_651),
.B(n_544),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_651),
.B(n_632),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_644),
.A2(n_198),
.B(n_196),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_593),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_683),
.A2(n_399),
.B(n_203),
.C(n_242),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_704),
.A2(n_399),
.B1(n_376),
.B2(n_184),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_631),
.A2(n_17),
.B(n_19),
.C(n_21),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_687),
.B(n_209),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_681),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_697),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_689),
.A2(n_376),
.B(n_434),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_723),
.B(n_215),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_696),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_724),
.A2(n_376),
.B(n_246),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_589),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_582),
.B(n_597),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_593),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_727),
.A2(n_247),
.B1(n_285),
.B2(n_253),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_733),
.B(n_252),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_609),
.B(n_21),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_591),
.A2(n_239),
.B(n_230),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_631),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_591),
.A2(n_619),
.B(n_603),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_714),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_734),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_618),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_603),
.A2(n_225),
.B(n_217),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_686),
.B(n_22),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_709),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_650),
.B(n_23),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_695),
.A2(n_27),
.B(n_28),
.C(n_32),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_640),
.B(n_27),
.Y(n_837)
);

AOI21x1_ASAP7_75t_L g838 ( 
.A1(n_692),
.A2(n_376),
.B(n_399),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_650),
.B(n_32),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_696),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_662),
.B(n_33),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_637),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_652),
.B(n_70),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_593),
.B(n_399),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_728),
.A2(n_692),
.B(n_699),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_646),
.B(n_36),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_730),
.B(n_37),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_593),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_614),
.B(n_180),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_644),
.B(n_37),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_684),
.B(n_180),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_699),
.A2(n_376),
.B(n_180),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_608),
.A2(n_376),
.B(n_180),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_691),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_657),
.Y(n_855)
);

NOR2x1_ASAP7_75t_L g856 ( 
.A(n_719),
.B(n_376),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_599),
.A2(n_85),
.B(n_142),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_691),
.B(n_42),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_610),
.A2(n_75),
.B(n_140),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_600),
.A2(n_62),
.B(n_138),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_616),
.A2(n_143),
.B(n_135),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_690),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_721),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_604),
.A2(n_128),
.B(n_121),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_633),
.B(n_42),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_634),
.B(n_44),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_46),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_694),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_731),
.B(n_47),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_636),
.B(n_50),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

O2A1O1Ixp5_ASAP7_75t_L g872 ( 
.A1(n_656),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_605),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_648),
.B(n_56),
.Y(n_874)
);

NOR2x1_ASAP7_75t_L g875 ( 
.A(n_613),
.B(n_602),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_594),
.B(n_622),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_641),
.A2(n_712),
.B(n_698),
.C(n_711),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_725),
.A2(n_726),
.B(n_718),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_712),
.B(n_732),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_694),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_700),
.A2(n_710),
.B(n_717),
.Y(n_881)
);

O2A1O1Ixp5_ASAP7_75t_L g882 ( 
.A1(n_656),
.A2(n_624),
.B(n_627),
.C(n_626),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_721),
.B(n_732),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_578),
.A2(n_606),
.B1(n_607),
.B2(n_617),
.Y(n_884)
);

INVx11_ASAP7_75t_L g885 ( 
.A(n_729),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_614),
.B(n_702),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_602),
.A2(n_624),
.B(n_659),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_722),
.A2(n_708),
.B(n_707),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_722),
.A2(n_693),
.B(n_614),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_669),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_620),
.B(n_671),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_626),
.B(n_627),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_682),
.A2(n_704),
.B1(n_675),
.B2(n_659),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_635),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_702),
.B(n_706),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_679),
.B(n_720),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_677),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_702),
.A2(n_617),
.B(n_664),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_658),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_702),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_618),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_660),
.A2(n_666),
.B(n_675),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_762),
.B(n_731),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_746),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_741),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_807),
.A2(n_639),
.B(n_618),
.C(n_706),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_835),
.A2(n_706),
.B(n_618),
.C(n_729),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_758),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_744),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_742),
.A2(n_706),
.B(n_729),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_757),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_858),
.B(n_729),
.C(n_706),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_758),
.B(n_784),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_736),
.A2(n_729),
.B(n_828),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_780),
.A2(n_876),
.B1(n_754),
.B2(n_797),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_762),
.B(n_834),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_869),
.A2(n_767),
.B1(n_814),
.B2(n_835),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_869),
.A2(n_797),
.B1(n_753),
.B2(n_850),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_839),
.A2(n_874),
.B(n_777),
.C(n_802),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_892),
.A2(n_747),
.B(n_878),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_833),
.A2(n_879),
.B1(n_787),
.B2(n_801),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_739),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_737),
.A2(n_752),
.B(n_763),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_761),
.Y(n_924)
);

INVxp33_ASAP7_75t_SL g925 ( 
.A(n_774),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_768),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_775),
.A2(n_815),
.B1(n_830),
.B2(n_749),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_764),
.B(n_814),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_770),
.A2(n_889),
.B(n_895),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_845),
.A2(n_794),
.B(n_789),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_777),
.B(n_896),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_882),
.A2(n_791),
.B(n_884),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_894),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_764),
.B(n_745),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_899),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_766),
.B(n_890),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_839),
.A2(n_735),
.B1(n_891),
.B2(n_874),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_766),
.A2(n_820),
.B1(n_738),
.B2(n_800),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_738),
.B(n_800),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_863),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_745),
.B(n_784),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_831),
.B(n_901),
.Y(n_942)
);

OR2x2_ASAP7_75t_SL g943 ( 
.A(n_806),
.B(n_841),
.Y(n_943)
);

AO32x1_ASAP7_75t_L g944 ( 
.A1(n_783),
.A2(n_755),
.A3(n_779),
.B1(n_867),
.B2(n_862),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_865),
.A2(n_870),
.B1(n_866),
.B2(n_799),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_821),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_808),
.B(n_873),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_829),
.A2(n_825),
.B1(n_781),
.B2(n_875),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_846),
.A2(n_756),
.B(n_882),
.C(n_851),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_821),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_SL g951 ( 
.A(n_831),
.B(n_901),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_831),
.B(n_901),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_854),
.A2(n_836),
.B(n_812),
.C(n_827),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_873),
.B(n_883),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_759),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_782),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_837),
.A2(n_811),
.B1(n_825),
.B2(n_765),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_798),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_796),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_795),
.A2(n_743),
.B(n_776),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_759),
.B(n_818),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_897),
.Y(n_962)
);

BUFx2_ASAP7_75t_R g963 ( 
.A(n_842),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_897),
.B(n_818),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_840),
.B(n_813),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_769),
.A2(n_877),
.B(n_785),
.C(n_843),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_868),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_880),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_796),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_871),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_840),
.B(n_809),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_888),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_817),
.B(n_824),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_792),
.B(n_748),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_751),
.A2(n_792),
.B1(n_893),
.B2(n_900),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_855),
.A2(n_811),
.B1(n_864),
.B2(n_857),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_810),
.A2(n_872),
.B(n_788),
.C(n_823),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_750),
.B(n_848),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_786),
.A2(n_773),
.B(n_772),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_871),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_796),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_849),
.A2(n_887),
.B(n_803),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_796),
.B(n_822),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_804),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_760),
.A2(n_803),
.B(n_790),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_SL g986 ( 
.A1(n_860),
.A2(n_822),
.B1(n_900),
.B2(n_809),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_SL g987 ( 
.A1(n_819),
.A2(n_832),
.B1(n_826),
.B2(n_872),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_804),
.B(n_900),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_881),
.A2(n_902),
.B1(n_849),
.B2(n_778),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_804),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_804),
.B(n_809),
.Y(n_991)
);

AO32x2_ASAP7_75t_L g992 ( 
.A1(n_886),
.A2(n_793),
.A3(n_861),
.B1(n_853),
.B2(n_838),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_898),
.A2(n_844),
.B(n_771),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_809),
.B(n_822),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_852),
.A2(n_844),
.B(n_856),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_822),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_805),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_885),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_859),
.A2(n_584),
.B(n_575),
.C(n_591),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_816),
.B(n_762),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_762),
.B(n_574),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_762),
.B(n_574),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_762),
.B(n_574),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_797),
.B(n_301),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_SL g1007 ( 
.A1(n_740),
.A2(n_584),
.B(n_575),
.C(n_591),
.Y(n_1007)
);

AO32x2_ASAP7_75t_L g1008 ( 
.A1(n_747),
.A2(n_884),
.A3(n_749),
.B1(n_695),
.B2(n_755),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_741),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_757),
.A2(n_410),
.B1(n_443),
.B2(n_574),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_R g1012 ( 
.A(n_757),
.B(n_443),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_767),
.B(n_574),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_740),
.A2(n_587),
.B(n_839),
.C(n_835),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_740),
.A2(n_587),
.B(n_839),
.C(n_835),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_797),
.B(n_301),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_797),
.B(n_301),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_780),
.B(n_443),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_758),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_780),
.B(n_443),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_740),
.A2(n_587),
.B(n_839),
.C(n_835),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_741),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_869),
.A2(n_464),
.B1(n_767),
.B2(n_485),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_797),
.B(n_301),
.Y(n_1026)
);

OR2x6_ASAP7_75t_SL g1027 ( 
.A(n_757),
.B(n_301),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_764),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_807),
.A2(n_740),
.B(n_850),
.C(n_478),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_780),
.B(n_443),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_740),
.A2(n_587),
.B(n_839),
.C(n_835),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_740),
.A2(n_742),
.B(n_736),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_762),
.B(n_574),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_740),
.A2(n_587),
.B(n_839),
.C(n_835),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_762),
.B(n_574),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_764),
.B(n_680),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_757),
.Y(n_1039)
);

AO21x1_ASAP7_75t_L g1040 ( 
.A1(n_740),
.A2(n_802),
.B(n_850),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_929),
.A2(n_930),
.B(n_960),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_922),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_923),
.A2(n_979),
.B(n_985),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1032),
.A2(n_1036),
.B(n_919),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_918),
.B(n_976),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_932),
.A2(n_1005),
.B(n_1002),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_999),
.A2(n_920),
.B(n_1007),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_921),
.A2(n_918),
.B(n_937),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_911),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1020),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_1034),
.B(n_1033),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_904),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1013),
.B(n_1025),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_905),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_932),
.A2(n_949),
.B(n_1040),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_993),
.A2(n_995),
.B(n_982),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_995),
.A2(n_910),
.B(n_914),
.Y(n_1058)
);

INVx6_ASAP7_75t_SL g1059 ( 
.A(n_1038),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_1006),
.B(n_1016),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1017),
.B(n_1026),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_909),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_908),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1004),
.B(n_1035),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_945),
.B(n_1030),
.C(n_1011),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1037),
.A2(n_931),
.B1(n_916),
.B2(n_917),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_973),
.A2(n_965),
.B(n_971),
.C(n_961),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_SL g1068 ( 
.A1(n_1012),
.A2(n_957),
.B1(n_903),
.B2(n_947),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1000),
.A2(n_986),
.B(n_951),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_924),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_989),
.A2(n_972),
.B(n_975),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_942),
.A2(n_952),
.B(n_977),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_907),
.A2(n_957),
.A3(n_927),
.B(n_940),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_908),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_1039),
.B(n_981),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_1038),
.B(n_934),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_944),
.A2(n_950),
.B(n_946),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_944),
.A2(n_964),
.B(n_994),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_936),
.B(n_1031),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_962),
.A2(n_958),
.A3(n_968),
.B(n_956),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_983),
.A2(n_1021),
.B(n_1018),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_997),
.A2(n_987),
.B(n_988),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_925),
.A2(n_967),
.B1(n_935),
.B2(n_933),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_997),
.A2(n_955),
.B(n_974),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_955),
.A2(n_984),
.B(n_906),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_953),
.A2(n_990),
.B(n_912),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_954),
.A2(n_948),
.B(n_996),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_915),
.B(n_938),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_1027),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_990),
.A2(n_969),
.B(n_991),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_969),
.A2(n_1024),
.B(n_1009),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_969),
.A2(n_926),
.B(n_1008),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_943),
.Y(n_1093)
);

AO21x1_ASAP7_75t_L g1094 ( 
.A1(n_939),
.A2(n_978),
.B(n_1008),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_970),
.A2(n_980),
.B(n_913),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_992),
.A2(n_998),
.A3(n_959),
.B(n_980),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_928),
.Y(n_1097)
);

AOI211x1_ASAP7_75t_L g1098 ( 
.A1(n_913),
.A2(n_992),
.B(n_941),
.C(n_959),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_992),
.A2(n_959),
.A3(n_1029),
.B(n_934),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1038),
.A2(n_934),
.B(n_941),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1019),
.A2(n_908),
.B(n_963),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1006),
.B(n_472),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_919),
.A2(n_1014),
.B(n_1022),
.C(n_1015),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_928),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_1014),
.A2(n_1015),
.B(n_1032),
.C(n_1022),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_922),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1013),
.B(n_1025),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_918),
.A2(n_937),
.B1(n_410),
.B2(n_869),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_SL g1109 ( 
.A(n_911),
.B(n_1039),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_922),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_919),
.A2(n_1014),
.B(n_1022),
.C(n_1015),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_966),
.A2(n_923),
.B(n_945),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1113)
);

NAND2x1_ASAP7_75t_L g1114 ( 
.A(n_970),
.B(n_871),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_932),
.A2(n_930),
.B(n_923),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1040),
.A2(n_945),
.A3(n_756),
.B(n_966),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_922),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_908),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_905),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1014),
.A2(n_1022),
.B(n_1015),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_905),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_905),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1013),
.B(n_767),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_904),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1014),
.A2(n_1022),
.B1(n_1032),
.B2(n_1015),
.Y(n_1129)
);

AO32x2_ASAP7_75t_L g1130 ( 
.A1(n_921),
.A2(n_918),
.A3(n_986),
.B1(n_945),
.B2(n_927),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_1013),
.B(n_1025),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1040),
.A2(n_945),
.A3(n_756),
.B(n_966),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_928),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_919),
.A2(n_1014),
.B(n_1022),
.C(n_1015),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_918),
.A2(n_937),
.B1(n_410),
.B2(n_869),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_SL g1138 ( 
.A(n_1001),
.B(n_663),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_908),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1014),
.A2(n_1015),
.B1(n_1032),
.B2(n_1022),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1038),
.B(n_934),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_929),
.A2(n_930),
.B(n_960),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_922),
.Y(n_1147)
);

AO32x2_ASAP7_75t_L g1148 ( 
.A1(n_921),
.A2(n_918),
.A3(n_986),
.B1(n_945),
.B2(n_927),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_922),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1013),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_929),
.A2(n_930),
.B(n_960),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_904),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_928),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_904),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_SL g1155 ( 
.A1(n_921),
.A2(n_918),
.B(n_1040),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_911),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1014),
.A2(n_1022),
.B(n_1032),
.C(n_1015),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_905),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_911),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1014),
.A2(n_740),
.B(n_1015),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_919),
.A2(n_1014),
.B(n_1022),
.C(n_1015),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_1049),
.B2(n_1046),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1130),
.B(n_1148),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1153),
.Y(n_1167)
);

AOI22x1_ASAP7_75t_L g1168 ( 
.A1(n_1113),
.A2(n_1162),
.B1(n_1117),
.B2(n_1156),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1046),
.A2(n_1049),
.B1(n_1068),
.B2(n_1093),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_1110),
.Y(n_1170)
);

BUFx8_ASAP7_75t_L g1171 ( 
.A(n_1147),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1065),
.A2(n_1054),
.B1(n_1107),
.B2(n_1131),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1062),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1070),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1088),
.A2(n_1127),
.B1(n_1065),
.B2(n_1066),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1096),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1123),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_1075),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1066),
.A2(n_1152),
.B1(n_1154),
.B2(n_1053),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_R g1180 ( 
.A1(n_1102),
.A2(n_1105),
.B1(n_1158),
.B2(n_1141),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1042),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1089),
.A2(n_1133),
.B1(n_1150),
.B2(n_1134),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_1161),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1125),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1103),
.A2(n_1136),
.B1(n_1164),
.B2(n_1111),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1161),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1130),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1044),
.B(n_1064),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1155),
.A2(n_1045),
.B1(n_1129),
.B2(n_1124),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1121),
.A2(n_1146),
.B1(n_1139),
.B2(n_1144),
.Y(n_1190)
);

BUFx8_ASAP7_75t_SL g1191 ( 
.A(n_1106),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1128),
.A2(n_1083),
.B1(n_1159),
.B2(n_1143),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1130),
.B(n_1148),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1138),
.A2(n_1104),
.B1(n_1097),
.B2(n_1135),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1148),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1084),
.B(n_1079),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1119),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1097),
.A2(n_1135),
.B1(n_1104),
.B2(n_1094),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1118),
.A2(n_1120),
.B(n_1163),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1050),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1126),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1099),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1087),
.A2(n_1081),
.B1(n_1059),
.B2(n_1076),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1073),
.B(n_1092),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1149),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1160),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1142),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1080),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1074),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1073),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1073),
.B(n_1077),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1112),
.A2(n_1056),
.B1(n_1069),
.B2(n_1100),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1063),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_SL g1215 ( 
.A(n_1157),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1101),
.A2(n_1112),
.B1(n_1091),
.B2(n_1086),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1056),
.A2(n_1071),
.B1(n_1082),
.B2(n_1085),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1109),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1078),
.A2(n_1140),
.B1(n_1122),
.B2(n_1072),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1140),
.A2(n_1090),
.B1(n_1047),
.B2(n_1048),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1067),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1047),
.A2(n_1115),
.B1(n_1095),
.B2(n_1058),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1115),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1057),
.A2(n_1114),
.B1(n_1051),
.B2(n_1052),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1116),
.B(n_1132),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1098),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1116),
.B(n_1132),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1041),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1145),
.B(n_1151),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1043),
.B(n_1130),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_1110),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1108),
.A2(n_1025),
.B1(n_1137),
.B2(n_611),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1142),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1161),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1096),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_1060),
.B2(n_1061),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1046),
.A2(n_869),
.B1(n_410),
.B2(n_611),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1108),
.A2(n_1025),
.B1(n_1137),
.B2(n_611),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_410),
.B2(n_1046),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1096),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1074),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1074),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1110),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1055),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1044),
.B(n_1064),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1108),
.A2(n_1025),
.B1(n_1137),
.B2(n_611),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1108),
.A2(n_1025),
.B1(n_1137),
.B2(n_611),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1142),
.Y(n_1248)
);

CKINVDCx14_ASAP7_75t_R g1249 ( 
.A(n_1075),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1055),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_410),
.B2(n_1046),
.Y(n_1251)
);

BUFx8_ASAP7_75t_L g1252 ( 
.A(n_1147),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1108),
.A2(n_1025),
.B1(n_1137),
.B2(n_611),
.Y(n_1253)
);

BUFx2_ASAP7_75t_SL g1254 ( 
.A(n_1093),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_SL g1255 ( 
.A(n_1074),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1130),
.B(n_1148),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1046),
.A2(n_869),
.B1(n_410),
.B2(n_611),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1076),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_410),
.B2(n_1046),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1046),
.A2(n_869),
.B1(n_410),
.B2(n_611),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1096),
.Y(n_1261)
);

CKINVDCx11_ASAP7_75t_R g1262 ( 
.A(n_1110),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1108),
.A2(n_1137),
.B1(n_410),
.B2(n_1046),
.Y(n_1263)
);

BUFx2_ASAP7_75t_R g1264 ( 
.A(n_1089),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1209),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1167),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1210),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1227),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1166),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1237),
.A2(n_1260),
.B1(n_1257),
.B2(n_1239),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1193),
.B(n_1256),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1193),
.B(n_1256),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1187),
.B(n_1195),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1187),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1195),
.B(n_1230),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1211),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1225),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1170),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1251),
.A2(n_1263),
.B(n_1259),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1207),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1225),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1236),
.A2(n_1169),
.B(n_1238),
.C(n_1246),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1210),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1228),
.Y(n_1285)
);

BUFx4f_ASAP7_75t_SL g1286 ( 
.A(n_1218),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1173),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1212),
.B(n_1205),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1228),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1174),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1221),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1184),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1201),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1223),
.B(n_1165),
.Y(n_1295)
);

INVx8_ASAP7_75t_L g1296 ( 
.A(n_1221),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1244),
.B(n_1250),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1176),
.B(n_1235),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1189),
.B(n_1261),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1229),
.A2(n_1168),
.B(n_1199),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1197),
.B(n_1206),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1226),
.B(n_1203),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1170),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1168),
.A2(n_1224),
.B(n_1222),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_1245),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1220),
.A2(n_1240),
.B(n_1219),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1185),
.A2(n_1216),
.B(n_1247),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1240),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1261),
.A2(n_1196),
.B(n_1198),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1213),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1217),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1179),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1232),
.B(n_1253),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1172),
.B(n_1254),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1180),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1274),
.B(n_1254),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1274),
.B(n_1182),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1277),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1276),
.B(n_1194),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1267),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1277),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1272),
.B(n_1204),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1286),
.B(n_1200),
.Y(n_1324)
);

AOI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1316),
.A2(n_1192),
.B1(n_1215),
.B2(n_1200),
.C(n_1241),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1300),
.A2(n_1248),
.B(n_1233),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1267),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1272),
.B(n_1214),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1284),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1278),
.B(n_1282),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1273),
.B(n_1208),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1283),
.A2(n_1249),
.B(n_1178),
.C(n_1241),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1316),
.A2(n_1178),
.B1(n_1249),
.B2(n_1218),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1285),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1279),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1305),
.B(n_1181),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1308),
.A2(n_1242),
.B(n_1202),
.C(n_1258),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1281),
.B(n_1181),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1270),
.A2(n_1255),
.B(n_1191),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1301),
.B(n_1191),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1306),
.A2(n_1215),
.B(n_1255),
.C(n_1264),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_SL g1343 ( 
.A1(n_1303),
.A2(n_1231),
.B(n_1243),
.C(n_1262),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1265),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_SL g1345 ( 
.A1(n_1266),
.A2(n_1231),
.B(n_1243),
.C(n_1262),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1288),
.B(n_1183),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1269),
.B(n_1271),
.Y(n_1347)
);

INVx5_ASAP7_75t_SL g1348 ( 
.A(n_1280),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1269),
.B(n_1271),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1299),
.B(n_1186),
.Y(n_1350)
);

NAND4xp25_ASAP7_75t_L g1351 ( 
.A(n_1315),
.B(n_1186),
.C(n_1234),
.D(n_1171),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1284),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1287),
.B(n_1234),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1171),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1297),
.B(n_1252),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1275),
.B(n_1252),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1297),
.B(n_1268),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1280),
.A2(n_1314),
.B1(n_1295),
.B2(n_1315),
.Y(n_1358)
);

AOI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1312),
.A2(n_1311),
.B1(n_1295),
.B2(n_1314),
.C(n_1292),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1300),
.A2(n_1304),
.B(n_1311),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1313),
.A2(n_1307),
.B(n_1296),
.C(n_1298),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1304),
.A2(n_1307),
.B(n_1309),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1359),
.A2(n_1313),
.B1(n_1310),
.B2(n_1302),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1319),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1326),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1322),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1347),
.B(n_1289),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1347),
.B(n_1289),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1349),
.B(n_1289),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1326),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1337),
.B(n_1291),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1326),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1318),
.B(n_1290),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1349),
.B(n_1289),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1344),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1357),
.B(n_1328),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1318),
.B(n_1357),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1334),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1334),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1358),
.B(n_1293),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1336),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1330),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1378),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1376),
.B(n_1367),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1379),
.B(n_1331),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1378),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1378),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1381),
.B(n_1302),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1366),
.Y(n_1391)
);

AO221x2_ASAP7_75t_L g1392 ( 
.A1(n_1383),
.A2(n_1340),
.B1(n_1333),
.B2(n_1339),
.C(n_1355),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1378),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1367),
.B(n_1362),
.Y(n_1394)
);

AND4x1_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1332),
.C(n_1342),
.D(n_1354),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1363),
.A2(n_1325),
.B1(n_1348),
.B2(n_1354),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1381),
.A2(n_1361),
.B1(n_1338),
.B2(n_1351),
.C(n_1356),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1370),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1380),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1365),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1364),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1379),
.B(n_1348),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1365),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1371),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1375),
.B(n_1320),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1382),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1369),
.B(n_1374),
.Y(n_1409)
);

AND4x1_ASAP7_75t_L g1410 ( 
.A(n_1371),
.B(n_1324),
.C(n_1341),
.D(n_1350),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1375),
.B(n_1294),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1411),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1411),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1391),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1410),
.B(n_1379),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1410),
.B(n_1343),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1410),
.B(n_1335),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1399),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1399),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1391),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1399),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1385),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1385),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1401),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1407),
.B(n_1373),
.Y(n_1425)
);

AND2x2_ASAP7_75t_SL g1426 ( 
.A(n_1395),
.B(n_1381),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1386),
.B(n_1409),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1365),
.Y(n_1428)
);

NAND2x1_ASAP7_75t_L g1429 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1395),
.A2(n_1381),
.B1(n_1379),
.B2(n_1372),
.C(n_1365),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1403),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1403),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1399),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1377),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1408),
.B(n_1373),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1394),
.B(n_1369),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1387),
.B(n_1377),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1394),
.B(n_1369),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1406),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1387),
.B(n_1377),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1441)
);

NOR3xp33_ASAP7_75t_L g1442 ( 
.A(n_1397),
.B(n_1351),
.C(n_1372),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1440),
.B(n_1377),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1414),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1422),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1414),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1427),
.B(n_1401),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1420),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1423),
.B(n_1398),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1420),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1440),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1440),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1423),
.B(n_1422),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1437),
.B(n_1387),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1437),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1398),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1431),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1435),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1441),
.B(n_1400),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1430),
.A2(n_1396),
.B1(n_1415),
.B2(n_1397),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1426),
.A2(n_1396),
.B1(n_1390),
.B2(n_1404),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1412),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1439),
.B(n_1335),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1442),
.B(n_1441),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1412),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1413),
.Y(n_1469)
);

OAI21xp33_ASAP7_75t_L g1470 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1401),
.Y(n_1470)
);

NAND2x1_ASAP7_75t_L g1471 ( 
.A(n_1424),
.B(n_1384),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1413),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1417),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1442),
.A2(n_1395),
.B(n_1396),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1434),
.B(n_1373),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1431),
.Y(n_1476)
);

NOR2xp67_ASAP7_75t_L g1477 ( 
.A(n_1441),
.B(n_1389),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1427),
.B(n_1400),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1439),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1418),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1418),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1434),
.B(n_1373),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1418),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1432),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1461),
.B(n_1425),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1452),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1458),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1445),
.B(n_1452),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1479),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1458),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1444),
.B(n_1425),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1476),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1416),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1465),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1480),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1471),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1474),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1446),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1460),
.B(n_1427),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1460),
.B(n_1436),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1447),
.B(n_1424),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1484),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1480),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1448),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1447),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1462),
.A2(n_1390),
.B1(n_1404),
.B2(n_1392),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1481),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1424),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1450),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1459),
.B(n_1432),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1478),
.B(n_1436),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1451),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1481),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1345),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1438),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1453),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1464),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1466),
.A2(n_1406),
.B1(n_1404),
.B2(n_1390),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1489),
.B(n_1454),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1457),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1494),
.B(n_1456),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1487),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1487),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1506),
.A2(n_1470),
.B1(n_1463),
.B2(n_1494),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1497),
.A2(n_1392),
.B1(n_1390),
.B2(n_1350),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1486),
.B(n_1449),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1492),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1438),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1516),
.A2(n_1443),
.B1(n_1455),
.B2(n_1471),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1493),
.A2(n_1429),
.B(n_1392),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

OAI32xp33_ASAP7_75t_L g1539 ( 
.A1(n_1519),
.A2(n_1455),
.A3(n_1443),
.B1(n_1482),
.B2(n_1475),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1519),
.A2(n_1392),
.B1(n_1390),
.B2(n_1483),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1515),
.B(n_1429),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1475),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1502),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1530),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1537),
.A2(n_1488),
.B(n_1498),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1523),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1543),
.B(n_1488),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1530),
.A2(n_1498),
.B(n_1501),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1524),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1538),
.Y(n_1551)
);

AO22x1_ASAP7_75t_L g1552 ( 
.A1(n_1531),
.A2(n_1486),
.B1(n_1538),
.B2(n_1541),
.Y(n_1552)
);

OAI322xp33_ASAP7_75t_L g1553 ( 
.A1(n_1525),
.A2(n_1520),
.A3(n_1521),
.B1(n_1486),
.B2(n_1522),
.C1(n_1533),
.C2(n_1540),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1532),
.A2(n_1501),
.B1(n_1496),
.B2(n_1511),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1536),
.A2(n_1513),
.B1(n_1495),
.B2(n_1507),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1527),
.B(n_1512),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1539),
.A2(n_1518),
.B1(n_1517),
.B2(n_1512),
.C(n_1509),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1541),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1514),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1531),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1531),
.B(n_1496),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1517),
.C(n_1509),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1534),
.A2(n_1508),
.B(n_1504),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1545),
.Y(n_1564)
);

AOI32xp33_ASAP7_75t_L g1565 ( 
.A1(n_1557),
.A2(n_1544),
.A3(n_1542),
.B1(n_1526),
.B2(n_1528),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1559),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1551),
.B(n_1518),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1555),
.A2(n_1485),
.B1(n_1491),
.B2(n_1513),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_L g1569 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1548),
.B(n_1508),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1556),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1546),
.A2(n_1535),
.B(n_1510),
.C(n_1511),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1561),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1562),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1566),
.B(n_1560),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1568),
.B(n_1561),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1564),
.B(n_1558),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1570),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1569),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1573),
.B(n_1553),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1567),
.Y(n_1582)
);

NAND4xp25_ASAP7_75t_L g1583 ( 
.A(n_1574),
.B(n_1571),
.C(n_1572),
.D(n_1567),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1566),
.B(n_1552),
.Y(n_1584)
);

NAND4xp25_ASAP7_75t_L g1585 ( 
.A(n_1578),
.B(n_1563),
.C(n_1550),
.D(n_1547),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1579),
.A2(n_1554),
.B1(n_1485),
.B2(n_1510),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1575),
.Y(n_1587)
);

AOI311xp33_ASAP7_75t_L g1588 ( 
.A1(n_1577),
.A2(n_1491),
.A3(n_1468),
.B(n_1469),
.C(n_1472),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1583),
.B(n_1508),
.Y(n_1589)
);

OAI32xp33_ASAP7_75t_L g1590 ( 
.A1(n_1581),
.A2(n_1513),
.A3(n_1507),
.B1(n_1503),
.B2(n_1495),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1584),
.A2(n_1582),
.B1(n_1577),
.B2(n_1580),
.C(n_1576),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1589),
.A2(n_1507),
.B1(n_1503),
.B2(n_1495),
.Y(n_1592)
);

OAI211xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1587),
.A2(n_1586),
.B(n_1591),
.C(n_1588),
.Y(n_1593)
);

AOI211xp5_ASAP7_75t_L g1594 ( 
.A1(n_1585),
.A2(n_1508),
.B(n_1535),
.C(n_1511),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1590),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1587),
.Y(n_1596)
);

AOI221x1_ASAP7_75t_L g1597 ( 
.A1(n_1585),
.A2(n_1503),
.B1(n_1483),
.B2(n_1424),
.C(n_1428),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_1595),
.B(n_1500),
.C(n_1353),
.Y(n_1598)
);

NAND4xp75_ASAP7_75t_L g1599 ( 
.A(n_1597),
.B(n_1500),
.C(n_1499),
.D(n_1346),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1596),
.Y(n_1600)
);

XNOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1592),
.B(n_1356),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1594),
.B(n_1499),
.Y(n_1602)
);

XOR2xp5_ASAP7_75t_L g1603 ( 
.A(n_1601),
.B(n_1593),
.Y(n_1603)
);

NOR4xp75_ASAP7_75t_L g1604 ( 
.A(n_1599),
.B(n_1389),
.C(n_1405),
.D(n_1402),
.Y(n_1604)
);

NOR4xp25_ASAP7_75t_L g1605 ( 
.A(n_1600),
.B(n_1602),
.C(n_1598),
.D(n_1421),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1603),
.Y(n_1606)
);

AO22x2_ASAP7_75t_L g1607 ( 
.A1(n_1606),
.A2(n_1605),
.B1(n_1604),
.B2(n_1428),
.Y(n_1607)
);

NOR2x1_ASAP7_75t_L g1608 ( 
.A(n_1607),
.B(n_1424),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1607),
.A2(n_1424),
.B(n_1428),
.Y(n_1609)
);

AOI22x1_ASAP7_75t_L g1610 ( 
.A1(n_1608),
.A2(n_1428),
.B1(n_1388),
.B2(n_1393),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1609),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1610),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1611),
.A2(n_1419),
.B1(n_1421),
.B2(n_1433),
.C(n_1428),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1612),
.A2(n_1482),
.B(n_1421),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_1613),
.B(n_1408),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1321),
.B1(n_1327),
.B2(n_1329),
.Y(n_1616)
);

OAI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1616),
.A2(n_1327),
.B1(n_1321),
.B2(n_1352),
.C(n_1329),
.Y(n_1617)
);

AOI211xp5_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1352),
.B(n_1291),
.C(n_1346),
.Y(n_1618)
);


endmodule