module fake_netlist_6_4796_n_110 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_110);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_110;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp67_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_22),
.B(n_32),
.C(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_33),
.B(n_43),
.C(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_34),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2x1p5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_47),
.B(n_46),
.Y(n_61)
);

AO31x2_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_60),
.A3(n_28),
.B(n_24),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_48),
.B(n_53),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_54),
.B1(n_39),
.B2(n_49),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_18),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_67)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_52),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_0),
.C(n_4),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_66),
.B(n_8),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_64),
.Y(n_73)
);

NOR2xp67_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_72),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_67),
.C(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_82),
.B1(n_84),
.B2(n_83),
.Y(n_95)
);

OAI211xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_84),
.B(n_90),
.C(n_5),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_91),
.C(n_92),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_92),
.B1(n_68),
.B2(n_63),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_63),
.B(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_5),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_103),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_101),
.B1(n_102),
.B2(n_7),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_102),
.B(n_65),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_104),
.B1(n_107),
.B2(n_61),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_61),
.C(n_62),
.Y(n_110)
);


endmodule