module fake_jpeg_20770_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_16),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_8),
.B1(n_13),
.B2(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_11),
.B1(n_10),
.B2(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_17),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_10),
.C(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_25),
.B1(n_13),
.B2(n_11),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_8),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_28),
.C(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_30),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_37),
.C(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_35),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_34),
.B(n_33),
.C(n_14),
.D(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_7),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_44),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_50),
.B1(n_49),
.B2(n_3),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.C(n_54),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_0),
.C(n_1),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_0),
.C(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_4),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_6),
.Y(n_62)
);


endmodule