module fake_ariane_2355_n_2279 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2279);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2279;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_212),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_43),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_87),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_165),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_126),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_92),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_83),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_85),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_55),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_64),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_182),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_164),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_133),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_171),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_76),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_116),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_166),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_106),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_127),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_123),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_168),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_60),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_54),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_134),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_2),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_58),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_13),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_178),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_136),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_47),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_185),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_203),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_73),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_55),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_70),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_45),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_172),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_163),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_190),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_72),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_191),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_47),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_156),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_74),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_111),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_64),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_66),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_115),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_200),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_181),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_90),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_63),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_52),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_152),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_77),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_141),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_88),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_41),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_32),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_5),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_148),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_27),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_154),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_173),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_71),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_221),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_80),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_59),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_66),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_59),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_175),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_29),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_135),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_25),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_81),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_13),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_35),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_99),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_137),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_187),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_62),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_22),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_15),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_197),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_24),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_101),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_31),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_161),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_176),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_78),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_193),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_142),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_54),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_51),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_206),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_60),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_20),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_43),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_42),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_195),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_79),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_26),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_104),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_73),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_39),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_63),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_149),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_145),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_125),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_113),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_52),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_89),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_216),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_109),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_95),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_2),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_44),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_97),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_34),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_108),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_103),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_84),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_37),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_122),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_72),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_131),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_21),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_140),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_58),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_67),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_138),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_202),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_158),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_17),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_14),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_75),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_45),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_18),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_204),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_67),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_68),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_143),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_57),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_207),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_147),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_198),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_36),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_0),
.Y(n_421)
);

BUFx8_ASAP7_75t_SL g422 ( 
.A(n_5),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_4),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_128),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_19),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_114),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_8),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_78),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_28),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_4),
.Y(n_430)
);

BUFx2_ASAP7_75t_R g431 ( 
.A(n_186),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_6),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_177),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_57),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_170),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_196),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_209),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_224),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_422),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_366),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_242),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_239),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_224),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_245),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_334),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_333),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_235),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_381),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_243),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_347),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_243),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_249),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_333),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_326),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_242),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_249),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_250),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_387),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_391),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_250),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_242),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_417),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_242),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_226),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_233),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_251),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_226),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_236),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_251),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_252),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_236),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_369),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_316),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_244),
.B(n_0),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_297),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_329),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_297),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_340),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_340),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_238),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_247),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_415),
.B(n_1),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_385),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_252),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_259),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_415),
.B(n_6),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_354),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_372),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_263),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_R g497 ( 
.A(n_222),
.B(n_82),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_390),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_333),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_278),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_231),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_256),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_279),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_421),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_256),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_283),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_260),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_398),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_363),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_260),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_225),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_346),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_287),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_268),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_268),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_288),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_398),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_272),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_272),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_289),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_242),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_292),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_286),
.B(n_8),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_346),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_225),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_246),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_273),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_273),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_346),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_299),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_246),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_368),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_280),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_368),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_280),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_303),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_301),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_303),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_302),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_311),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_311),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_335),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_307),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_242),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_335),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_368),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_349),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_257),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_257),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_367),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_286),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_286),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_310),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_269),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_444),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_443),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_349),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_465),
.A2(n_281),
.B(n_351),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_351),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_448),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_465),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_440),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_451),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_446),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_462),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_463),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_469),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_466),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_445),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_458),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_441),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_467),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_447),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_478),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_552),
.A2(n_281),
.B(n_357),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_485),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_486),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_481),
.B(n_431),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_490),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_552),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_447),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_450),
.A2(n_281),
.B(n_357),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_496),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_498),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_452),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_454),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_494),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_359),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_473),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_501),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_495),
.B(n_313),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_460),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_461),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_517),
.B(n_282),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_464),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_504),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_513),
.B(n_359),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_464),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_470),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_507),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_470),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_514),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_499),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_474),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_475),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_548),
.B(n_244),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_518),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_489),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_505),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_548),
.B(n_364),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_489),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_506),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_508),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_487),
.B(n_367),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_522),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_508),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_511),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_511),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_532),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_515),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_516),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_516),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_439),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_541),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_545),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_601),
.B(n_439),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_613),
.B(n_449),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_627),
.A2(n_442),
.B1(n_492),
.B2(n_472),
.Y(n_654)
);

INVxp33_ASAP7_75t_SL g655 ( 
.A(n_585),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_566),
.B(n_502),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_576),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_558),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_558),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_566),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_566),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_597),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_627),
.B(n_456),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_578),
.B(n_364),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_566),
.B(n_502),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_581),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_592),
.B(n_453),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_597),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_597),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_613),
.B(n_500),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_566),
.B(n_509),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_519),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_648),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_581),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_627),
.A2(n_472),
.B1(n_525),
.B2(n_477),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_453),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_459),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_591),
.B(n_459),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_574),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_586),
.A2(n_488),
.B1(n_555),
.B2(n_482),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_588),
.A2(n_488),
.B1(n_556),
.B2(n_457),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_594),
.A2(n_479),
.B1(n_483),
.B2(n_480),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_591),
.B(n_520),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_591),
.B(n_521),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_596),
.B(n_617),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_627),
.B(n_517),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_597),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_592),
.B(n_438),
.C(n_491),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_597),
.Y(n_697)
);

NAND2x1p5_ASAP7_75t_L g698 ( 
.A(n_593),
.B(n_561),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_564),
.Y(n_699)
);

INVxp33_ASAP7_75t_L g700 ( 
.A(n_607),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_590),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_595),
.B(n_484),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_564),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_604),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_603),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_615),
.B(n_526),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_574),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_608),
.B(n_493),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_627),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_559),
.Y(n_710)
);

AND3x2_ASAP7_75t_L g711 ( 
.A(n_608),
.B(n_493),
.C(n_524),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_619),
.A2(n_479),
.B1(n_318),
.B2(n_331),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_604),
.B(n_531),
.Y(n_713)
);

INVx3_ASAP7_75t_R g714 ( 
.A(n_568),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_596),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_605),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_367),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_605),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_617),
.B(n_521),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_534),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_610),
.B(n_374),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_638),
.A2(n_536),
.B1(n_529),
.B2(n_535),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_617),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_617),
.B(n_529),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_579),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_557),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_624),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_559),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_624),
.B(n_530),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_624),
.B(n_530),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_611),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_645),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_565),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_645),
.Y(n_736)
);

NOR2x1p5_ASAP7_75t_L g737 ( 
.A(n_621),
.B(n_628),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_645),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_611),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_559),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_626),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_565),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_565),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_632),
.B(n_539),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_639),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_601),
.B(n_510),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_645),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_632),
.B(n_553),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_643),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_598),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_598),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_568),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_559),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_633),
.B(n_554),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_598),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_602),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_633),
.B(n_634),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_600),
.A2(n_537),
.B1(n_540),
.B2(n_538),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_634),
.B(n_540),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_636),
.B(n_542),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_600),
.A2(n_542),
.B1(n_544),
.B2(n_543),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_650),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_651),
.B(n_543),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_636),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_631),
.A2(n_544),
.B1(n_549),
.B2(n_547),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_637),
.B(n_640),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_606),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_637),
.B(n_547),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_602),
.B(n_512),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_607),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_563),
.B(n_570),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_606),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_640),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_593),
.B(n_549),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_606),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_631),
.B(n_527),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_609),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_609),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_569),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_641),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_616),
.B(n_528),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_641),
.B(n_356),
.C(n_261),
.Y(n_785)
);

INVx6_ASAP7_75t_L g786 ( 
.A(n_559),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_616),
.A2(n_261),
.B1(n_284),
.B2(n_282),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_609),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_642),
.B(n_284),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_642),
.B(n_533),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_644),
.B(n_550),
.Y(n_791)
);

CKINVDCx11_ASAP7_75t_R g792 ( 
.A(n_648),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_644),
.B(n_551),
.Y(n_793)
);

BUFx4f_ASAP7_75t_L g794 ( 
.A(n_646),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_612),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_646),
.B(n_269),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_569),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_612),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_647),
.B(n_323),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_577),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_SL g801 ( 
.A(n_647),
.B(n_497),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_559),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_560),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_266),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_583),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_649),
.B(n_336),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_577),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_612),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_571),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_583),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_803),
.B(n_560),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_794),
.B(n_664),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_789),
.A2(n_562),
.B1(n_618),
.B2(n_614),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_683),
.B(n_572),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_803),
.B(n_562),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_754),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_685),
.B(n_789),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_SL g818 ( 
.A1(n_655),
.A2(n_599),
.B1(n_630),
.B2(n_622),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_730),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_745),
.B(n_750),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_794),
.B(n_614),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_683),
.B(n_573),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_779),
.B(n_614),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_713),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_684),
.B(n_618),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_758),
.B(n_575),
.C(n_275),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_794),
.B(n_618),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_620),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_708),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_777),
.B(n_620),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_664),
.B(n_620),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_779),
.B(n_623),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_801),
.A2(n_625),
.B1(n_629),
.B2(n_623),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_730),
.A2(n_625),
.B(n_629),
.C(n_623),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_784),
.B(n_629),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_664),
.B(n_635),
.Y(n_836)
);

NOR3x1_ASAP7_75t_L g837 ( 
.A(n_745),
.B(n_275),
.C(n_274),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_666),
.B(n_635),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_750),
.B(n_635),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_784),
.B(n_308),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_666),
.B(n_593),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_666),
.B(n_561),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_766),
.B(n_343),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_748),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_723),
.B(n_234),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_730),
.B(n_561),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_734),
.Y(n_847)
);

OAI221xp5_ASAP7_75t_L g848 ( 
.A1(n_787),
.A2(n_682),
.B1(n_654),
.B2(n_744),
.C(n_785),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_721),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_777),
.B(n_367),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_668),
.B(n_338),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_668),
.B(n_274),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_801),
.A2(n_286),
.B1(n_367),
.B2(n_296),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_668),
.B(n_433),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_761),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_793),
.B(n_296),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_709),
.A2(n_317),
.B1(n_380),
.B2(n_374),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_L g858 ( 
.A1(n_772),
.A2(n_402),
.B1(n_389),
.B2(n_293),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_677),
.B(n_389),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_L g860 ( 
.A1(n_760),
.A2(n_377),
.B1(n_379),
.B2(n_348),
.C(n_384),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_772),
.B(n_587),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_763),
.B(n_402),
.Y(n_862)
);

O2A1O1Ixp5_ASAP7_75t_L g863 ( 
.A1(n_734),
.A2(n_380),
.B(n_397),
.C(n_386),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_386),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_765),
.B(n_293),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_771),
.B(n_397),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_771),
.B(n_404),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_769),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_708),
.B(n_587),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_769),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_672),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_672),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_686),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_709),
.B(n_404),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_715),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_669),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_782),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_707),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_678),
.B(n_295),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_659),
.B(n_350),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_715),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_797),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_653),
.B(n_295),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_797),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_653),
.B(n_309),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_800),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_804),
.B(n_309),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_715),
.B(n_312),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_SL g890 ( 
.A1(n_655),
.A2(n_630),
.B1(n_622),
.B2(n_599),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_724),
.B(n_312),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_746),
.Y(n_892)
);

BUFx6f_ASAP7_75t_SL g893 ( 
.A(n_705),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_724),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_726),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_746),
.B(n_315),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_759),
.B(n_315),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_800),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_670),
.A2(n_320),
.B1(n_270),
.B2(n_383),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_736),
.B(n_747),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_736),
.B(n_584),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_749),
.A2(n_330),
.B(n_420),
.C(n_348),
.Y(n_902)
);

CKINVDCx11_ASAP7_75t_R g903 ( 
.A(n_705),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_676),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_756),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_736),
.B(n_324),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_805),
.B(n_324),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_747),
.B(n_584),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_676),
.A2(n_270),
.B1(n_383),
.B2(n_320),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_747),
.B(n_355),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_694),
.B(n_728),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_656),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_694),
.B(n_358),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_705),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_657),
.B(n_330),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_669),
.A2(n_367),
.B1(n_394),
.B2(n_580),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_658),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_728),
.B(n_360),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_660),
.B(n_339),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_665),
.A2(n_370),
.B(n_420),
.C(n_377),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_738),
.B(n_584),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_807),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_770),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_671),
.B(n_339),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_681),
.B(n_341),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_701),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_669),
.A2(n_262),
.B1(n_437),
.B2(n_285),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_770),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_704),
.B(n_341),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_765),
.B(n_345),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_716),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_737),
.B(n_345),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_807),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_719),
.B(n_370),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_733),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_739),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_738),
.B(n_234),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_669),
.A2(n_394),
.B1(n_582),
.B2(n_580),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_810),
.B(n_371),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_741),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_767),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_776),
.B(n_371),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_783),
.B(n_379),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_796),
.B(n_384),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_SL g945 ( 
.A1(n_700),
.A2(n_396),
.B1(n_410),
.B2(n_400),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_752),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_661),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_799),
.B(n_375),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_727),
.B(n_414),
.C(n_392),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_796),
.B(n_392),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_661),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_796),
.B(n_414),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_663),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_693),
.B(n_790),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_727),
.B(n_416),
.C(n_403),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_693),
.B(n_791),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_687),
.B(n_407),
.C(n_378),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_770),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_726),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_663),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_693),
.B(n_416),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_669),
.A2(n_722),
.B1(n_798),
.B2(n_775),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_669),
.Y(n_963)
);

NOR2x1p5_ASAP7_75t_L g964 ( 
.A(n_792),
.B(n_409),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_806),
.B(n_411),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_764),
.B(n_413),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_679),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_696),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_775),
.B(n_423),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_768),
.B(n_775),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_798),
.B(n_425),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_718),
.B(n_241),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_792),
.B(n_427),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_798),
.B(n_428),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_692),
.B(n_429),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_912),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_834),
.A2(n_777),
.B(n_674),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_825),
.B(n_762),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_844),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_830),
.A2(n_674),
.B(n_673),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_817),
.B(n_667),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_845),
.A2(n_722),
.B1(n_752),
.B2(n_757),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_849),
.B(n_809),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_879),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_905),
.A2(n_817),
.B1(n_824),
.B2(n_869),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_690),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_892),
.B(n_706),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_881),
.A2(n_688),
.B1(n_774),
.B2(n_722),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_914),
.B(n_680),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_921),
.A2(n_697),
.B(n_673),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_830),
.A2(n_697),
.B(n_698),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_871),
.A2(n_731),
.B1(n_732),
.B2(n_725),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_900),
.A2(n_698),
.B(n_675),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_917),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_921),
.A2(n_778),
.B(n_757),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_963),
.B(n_923),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_829),
.B(n_680),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_963),
.B(n_667),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_914),
.B(n_702),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_902),
.A2(n_956),
.B(n_954),
.C(n_835),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_850),
.A2(n_698),
.B(n_675),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_962),
.B(n_667),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_926),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_811),
.B(n_691),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_815),
.B(n_720),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_816),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_904),
.B(n_881),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_931),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_850),
.A2(n_841),
.B(n_842),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_841),
.A2(n_675),
.B(n_662),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_842),
.A2(n_695),
.B(n_662),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_823),
.B(n_722),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_902),
.A2(n_808),
.B(n_795),
.C(n_788),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_828),
.B(n_722),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_848),
.A2(n_751),
.B(n_795),
.C(n_788),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_901),
.A2(n_695),
.B(n_662),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_832),
.B(n_722),
.Y(n_1017)
);

AOI21x1_ASAP7_75t_L g1018 ( 
.A1(n_846),
.A2(n_699),
.B(n_679),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_908),
.A2(n_695),
.B(n_717),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_852),
.B(n_751),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_831),
.A2(n_838),
.B(n_836),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_838),
.A2(n_735),
.B(n_717),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_852),
.B(n_751),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_852),
.B(n_780),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_895),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_935),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_906),
.A2(n_712),
.B(n_742),
.C(n_743),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_843),
.A2(n_795),
.B(n_788),
.C(n_781),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_865),
.A2(n_742),
.B(n_743),
.C(n_753),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_872),
.B(n_652),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_846),
.A2(n_753),
.B(n_780),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_814),
.B(n_773),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_821),
.A2(n_781),
.B(n_780),
.C(n_703),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_959),
.B(n_689),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_851),
.B(n_781),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_821),
.A2(n_703),
.B(n_699),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_923),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_812),
.A2(n_667),
.B(n_748),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_863),
.A2(n_729),
.B(n_710),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_843),
.A2(n_281),
.B(n_271),
.C(n_277),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_827),
.A2(n_729),
.B(n_710),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_928),
.A2(n_652),
.B1(n_430),
.B2(n_432),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_873),
.B(n_711),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_819),
.B(n_748),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_969),
.A2(n_786),
.B1(n_802),
.B2(n_755),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_854),
.B(n_748),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_911),
.A2(n_580),
.B(n_577),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_819),
.B(n_755),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_847),
.A2(n_802),
.B(n_755),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_847),
.A2(n_867),
.B(n_911),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_958),
.B(n_755),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_876),
.A2(n_802),
.B(n_729),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_845),
.A2(n_700),
.B1(n_582),
.B2(n_277),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_959),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_969),
.A2(n_786),
.B1(n_802),
.B2(n_434),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_840),
.B(n_786),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_910),
.B(n_802),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_882),
.A2(n_729),
.B(n_710),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_786),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_936),
.Y(n_1061)
);

OAI321xp33_ASAP7_75t_L g1062 ( 
.A1(n_860),
.A2(n_321),
.A3(n_376),
.B1(n_241),
.B2(n_271),
.C(n_290),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_894),
.A2(n_729),
.B(n_710),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_826),
.B(n_918),
.C(n_913),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_855),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_971),
.A2(n_740),
.B(n_227),
.Y(n_1066)
);

AOI33xp33_ASAP7_75t_L g1067 ( 
.A1(n_858),
.A2(n_322),
.A3(n_321),
.B1(n_300),
.B2(n_290),
.B3(n_376),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_813),
.A2(n_322),
.B(n_435),
.C(n_582),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_865),
.B(n_714),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_940),
.A2(n_435),
.B1(n_740),
.B2(n_332),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_877),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_941),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_844),
.B(n_740),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_975),
.A2(n_948),
.B(n_965),
.C(n_839),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_975),
.B(n_223),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_930),
.B(n_228),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_856),
.A2(n_388),
.B(n_436),
.C(n_589),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_897),
.A2(n_388),
.B(n_436),
.C(n_589),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_974),
.A2(n_337),
.B(n_230),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_946),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_865),
.B(n_714),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_937),
.A2(n_589),
.B(n_436),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_844),
.A2(n_328),
.B(n_232),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_822),
.B(n_424),
.C(n_265),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_884),
.A2(n_589),
.B1(n_436),
.B2(n_388),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_820),
.B(n_9),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_918),
.B(n_342),
.C(n_237),
.Y(n_1087)
);

INVx11_ASAP7_75t_L g1088 ( 
.A(n_893),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_970),
.A2(n_864),
.B1(n_866),
.B2(n_868),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_949),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_1090)
);

BUFx12f_ASAP7_75t_L g1091 ( 
.A(n_903),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_877),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_884),
.B(n_229),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_947),
.A2(n_352),
.B(n_248),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_947),
.A2(n_353),
.B(n_253),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_884),
.B(n_240),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_948),
.A2(n_436),
.B(n_388),
.C(n_589),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_903),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_973),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_886),
.B(n_254),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_893),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_877),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_951),
.A2(n_362),
.B(n_258),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_886),
.B(n_888),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_951),
.A2(n_365),
.B(n_264),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_937),
.A2(n_589),
.B(n_436),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_886),
.B(n_255),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_953),
.A2(n_373),
.B(n_426),
.Y(n_1108)
);

AND2x6_ASAP7_75t_L g1109 ( 
.A(n_877),
.B(n_388),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_820),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_953),
.A2(n_361),
.B(n_419),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_878),
.A2(n_589),
.B(n_388),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_820),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_862),
.B(n_267),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_973),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_944),
.B(n_291),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_972),
.A2(n_418),
.B1(n_412),
.B2(n_406),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_861),
.B(n_10),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_960),
.A2(n_405),
.B(n_401),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_972),
.B(n_399),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_932),
.B(n_12),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_889),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_960),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_950),
.B(n_294),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_967),
.A2(n_395),
.B(n_393),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_870),
.B(n_16),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_891),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_818),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_875),
.A2(n_382),
.B(n_344),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_965),
.A2(n_327),
.B1(n_325),
.B2(n_319),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_920),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1131)
);

BUFx8_ASAP7_75t_L g1132 ( 
.A(n_968),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_909),
.A2(n_314),
.B(n_306),
.C(n_305),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_859),
.A2(n_94),
.B(n_217),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_952),
.B(n_304),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_883),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_961),
.B(n_298),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_883),
.A2(n_86),
.B(n_208),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_833),
.B(n_23),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_857),
.A2(n_23),
.B(n_24),
.Y(n_1140)
);

AO22x1_ASAP7_75t_L g1141 ( 
.A1(n_837),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_885),
.A2(n_96),
.B(n_205),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_915),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_896),
.B(n_30),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1104),
.B(n_880),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1006),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1033),
.A2(n_927),
.B(n_899),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_SL g1148 ( 
.A(n_1092),
.B(n_932),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_1132),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_991),
.A2(n_922),
.B(n_885),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_1029),
.A2(n_929),
.B(n_925),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1001),
.A2(n_922),
.B(n_933),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1033),
.A2(n_943),
.B(n_924),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1028),
.A2(n_919),
.B(n_942),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1058),
.A2(n_933),
.B(n_887),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1009),
.A2(n_887),
.B(n_898),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1018),
.A2(n_898),
.B(n_934),
.Y(n_1158)
);

OAI22x1_ASAP7_75t_L g1159 ( 
.A1(n_988),
.A2(n_964),
.B1(n_957),
.B2(n_890),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_1060),
.A2(n_966),
.B(n_920),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_985),
.B(n_907),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1028),
.A2(n_853),
.B(n_938),
.Y(n_1162)
);

AOI221x1_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_955),
.B1(n_945),
.B2(n_916),
.C(n_932),
.Y(n_1163)
);

INVx8_ASAP7_75t_L g1164 ( 
.A(n_1091),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1086),
.A2(n_939),
.B(n_33),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_984),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_983),
.B(n_30),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1039),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_993),
.A2(n_98),
.B(n_199),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1039),
.Y(n_1170)
);

AO22x1_ASAP7_75t_L g1171 ( 
.A1(n_1121),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_978),
.B(n_38),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1036),
.A2(n_100),
.B(n_194),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_982),
.B(n_38),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1015),
.A2(n_39),
.B(n_40),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1064),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1089),
.A2(n_112),
.B(n_184),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1092),
.B(n_1113),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1143),
.B(n_46),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_986),
.A2(n_110),
.B(n_183),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_977),
.A2(n_1048),
.B(n_1112),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_980),
.A2(n_107),
.B(n_179),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1117),
.A2(n_48),
.B(n_49),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1004),
.A2(n_93),
.B(n_174),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1088),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1007),
.B(n_48),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1015),
.A2(n_49),
.A3(n_50),
.B(n_51),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1005),
.A2(n_117),
.B(n_162),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1144),
.B(n_50),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_994),
.B(n_1003),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1008),
.B(n_53),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1032),
.B(n_53),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1025),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1026),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1061),
.B(n_56),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1031),
.A2(n_160),
.B(n_153),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_989),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1092),
.B(n_146),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1019),
.A2(n_130),
.B(n_120),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1128),
.B(n_56),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1072),
.B(n_61),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1121),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1010),
.A2(n_1011),
.B(n_1016),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1132),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1140),
.A2(n_70),
.B(n_75),
.C(n_77),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1050),
.A2(n_118),
.B(n_1074),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1000),
.A2(n_1090),
.B(n_1131),
.C(n_1122),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_995),
.A2(n_1021),
.B(n_1051),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1097),
.A2(n_1068),
.A3(n_1041),
.B(n_1077),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1127),
.B(n_1076),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_989),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_997),
.B(n_1030),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_990),
.A2(n_1106),
.B(n_1082),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1022),
.A2(n_1038),
.B(n_1053),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1110),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_982),
.A2(n_1075),
.B1(n_1117),
.B2(n_1080),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1055),
.B(n_1087),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1054),
.B(n_1069),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1098),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_981),
.A2(n_1002),
.B(n_1040),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1115),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1097),
.A2(n_1068),
.A3(n_1077),
.B(n_1078),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_981),
.A2(n_1066),
.B(n_1042),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1138),
.A2(n_1142),
.B(n_1059),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1045),
.A2(n_1049),
.B(n_1052),
.Y(n_1226)
);

BUFx2_ASAP7_75t_SL g1227 ( 
.A(n_999),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_987),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1045),
.A2(n_1049),
.B(n_1052),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1054),
.B(n_1069),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_979),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1063),
.A2(n_1027),
.B(n_1134),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_979),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1123),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_992),
.A2(n_1073),
.B(n_1046),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1081),
.B(n_1126),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1110),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1073),
.A2(n_1047),
.B(n_1139),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1012),
.A2(n_1014),
.B(n_1017),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_L g1240 ( 
.A1(n_1139),
.A2(n_1120),
.B(n_1013),
.C(n_1122),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1013),
.A2(n_1057),
.B(n_1035),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1120),
.A2(n_1057),
.B(n_998),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_998),
.A2(n_1079),
.B(n_1114),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1081),
.B(n_1084),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1020),
.A2(n_1024),
.B1(n_1023),
.B2(n_1037),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_979),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1084),
.B(n_1118),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1065),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1078),
.A2(n_1136),
.A3(n_1070),
.B(n_1133),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1030),
.B(n_1107),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1067),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1101),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_996),
.A2(n_1102),
.B(n_1071),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1092),
.B(n_1102),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_996),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1129),
.A2(n_1037),
.B(n_1135),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_979),
.B(n_1071),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1094),
.A2(n_1105),
.B(n_1125),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_999),
.B(n_1034),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1116),
.A2(n_1124),
.B(n_1137),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1095),
.A2(n_1103),
.B(n_1119),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1110),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1108),
.A2(n_1111),
.B(n_1056),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1044),
.A2(n_1043),
.B1(n_1086),
.B2(n_1130),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1085),
.A2(n_1083),
.B(n_1100),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1062),
.A2(n_1085),
.B(n_1133),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1109),
.A2(n_1044),
.B(n_1141),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1109),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1109),
.B(n_849),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1109),
.B(n_1092),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1109),
.B(n_686),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_991),
.A2(n_1001),
.B(n_993),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1001),
.A2(n_850),
.B(n_830),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_991),
.A2(n_1001),
.B(n_993),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_991),
.A2(n_1001),
.B(n_993),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_991),
.A2(n_1001),
.B(n_993),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1001),
.A2(n_850),
.B(n_830),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1104),
.B(n_849),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1104),
.B(n_849),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1001),
.A2(n_850),
.B(n_830),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1001),
.A2(n_850),
.B(n_830),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1104),
.B(n_849),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_SL g1284 ( 
.A1(n_1029),
.A2(n_1000),
.B(n_1021),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1091),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1132),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_991),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1104),
.B(n_849),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1104),
.B(n_849),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1104),
.B(n_849),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1033),
.A2(n_834),
.B(n_1028),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1033),
.A2(n_834),
.B(n_1028),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_984),
.B(n_686),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1025),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1025),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_976),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_976),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_976),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1029),
.A2(n_1000),
.B(n_1021),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1001),
.A2(n_850),
.B(n_830),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1294),
.A2(n_1295),
.B(n_1164),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1149),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1168),
.Y(n_1303)
);

CKINVDCx8_ASAP7_75t_R g1304 ( 
.A(n_1164),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1168),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1170),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1146),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1213),
.B(n_1197),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1145),
.B(n_1279),
.Y(n_1309)
);

BUFx2_ASAP7_75t_SL g1310 ( 
.A(n_1185),
.Y(n_1310)
);

AO21x1_ASAP7_75t_L g1311 ( 
.A1(n_1217),
.A2(n_1175),
.B(n_1267),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1156),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1213),
.B(n_1167),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1245),
.B(n_1161),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1174),
.A2(n_1265),
.B1(n_1165),
.B2(n_1260),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1178),
.B(n_1148),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1274),
.A2(n_1281),
.B(n_1278),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1293),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1194),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1174),
.A2(n_1260),
.B1(n_1288),
.B2(n_1280),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1296),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1297),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1251),
.B(n_1212),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1149),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1271),
.Y(n_1325)
);

INVx3_ASAP7_75t_SL g1326 ( 
.A(n_1294),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1178),
.B(n_1209),
.Y(n_1327)
);

AOI222xp33_ASAP7_75t_L g1328 ( 
.A1(n_1202),
.A2(n_1171),
.B1(n_1159),
.B2(n_1200),
.C1(n_1205),
.C2(n_1192),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1172),
.A2(n_1189),
.B(n_1248),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1283),
.B(n_1289),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1260),
.B(n_1170),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1209),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1285),
.B(n_1198),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1222),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1298),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1290),
.B(n_1219),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1166),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1282),
.A2(n_1300),
.B(n_1235),
.Y(n_1338)
);

INVx8_ASAP7_75t_L g1339 ( 
.A(n_1164),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1240),
.A2(n_1261),
.B(n_1205),
.C(n_1183),
.Y(n_1340)
);

INVx5_ASAP7_75t_L g1341 ( 
.A(n_1233),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1176),
.B(n_1163),
.C(n_1207),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1275),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1233),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1190),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1228),
.B(n_1227),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1271),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1207),
.A2(n_1186),
.B(n_1242),
.C(n_1211),
.Y(n_1348)
);

INVx5_ASAP7_75t_L g1349 ( 
.A(n_1233),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1178),
.B(n_1222),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1291),
.A2(n_1292),
.B(n_1181),
.Y(n_1351)
);

INVx8_ASAP7_75t_L g1352 ( 
.A(n_1253),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1198),
.A2(n_1246),
.B(n_1154),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1277),
.A2(n_1208),
.B(n_1206),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1230),
.A2(n_1236),
.B1(n_1252),
.B2(n_1249),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1234),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1271),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1244),
.A2(n_1152),
.B(n_1257),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1256),
.B(n_1237),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1263),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1181),
.A2(n_1243),
.B(n_1241),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1191),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1256),
.B(n_1153),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1215),
.A2(n_1287),
.B(n_1203),
.Y(n_1364)
);

AOI22x1_ASAP7_75t_L g1365 ( 
.A1(n_1226),
.A2(n_1229),
.B1(n_1262),
.B2(n_1151),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1231),
.B(n_1247),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1240),
.A2(n_1239),
.B(n_1238),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1195),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1201),
.Y(n_1369)
);

INVx3_ASAP7_75t_SL g1370 ( 
.A(n_1295),
.Y(n_1370)
);

BUFx2_ASAP7_75t_R g1371 ( 
.A(n_1204),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1287),
.A2(n_1225),
.B(n_1264),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1179),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1220),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1253),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1238),
.A2(n_1221),
.B(n_1147),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1185),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1233),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1204),
.B(n_1286),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1216),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1198),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1162),
.A2(n_1218),
.B1(n_1177),
.B2(n_1269),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1255),
.B(n_1286),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1149),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1231),
.B(n_1247),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1187),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1269),
.A2(n_1180),
.B1(n_1258),
.B2(n_1182),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1268),
.B(n_1255),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1187),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1187),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1225),
.A2(n_1299),
.B(n_1284),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1193),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1193),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1255),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1254),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_1155),
.B(n_1221),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1268),
.B(n_1254),
.Y(n_1398)
);

NOR3xp33_ASAP7_75t_L g1399 ( 
.A(n_1258),
.B(n_1188),
.C(n_1184),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1285),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1266),
.B(n_1250),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1187),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1196),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1266),
.B(n_1224),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1220),
.B(n_1250),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1250),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1158),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1250),
.B(n_1210),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1160),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1160),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1210),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1259),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1259),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1157),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1157),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1210),
.B(n_1223),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1214),
.A2(n_1150),
.B(n_1169),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1199),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1210),
.B(n_1223),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1223),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1223),
.B(n_1214),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1173),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1173),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1178),
.B(n_1148),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1165),
.A2(n_849),
.B1(n_988),
.B2(n_1161),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1174),
.A2(n_1161),
.B1(n_1064),
.B2(n_988),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1174),
.A2(n_845),
.B1(n_849),
.B2(n_462),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1168),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1146),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1197),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1149),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1168),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1220),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1185),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1156),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1213),
.B(n_983),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1274),
.A2(n_850),
.B(n_1278),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1233),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1213),
.B(n_983),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1197),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_SL g1442 ( 
.A(n_1294),
.B(n_959),
.Y(n_1442)
);

AND2x6_ASAP7_75t_L g1443 ( 
.A(n_1198),
.B(n_1271),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1145),
.B(n_978),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1174),
.A2(n_845),
.B1(n_849),
.B2(n_462),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1245),
.B(n_655),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1227),
.B(n_1212),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1178),
.B(n_1148),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1233),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1145),
.B(n_978),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1178),
.B(n_1148),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1145),
.B(n_978),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1209),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1209),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1197),
.B(n_1161),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1279),
.B(n_1280),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1271),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1149),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1245),
.B(n_655),
.Y(n_1459)
);

BUFx4f_ASAP7_75t_L g1460 ( 
.A(n_1149),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1220),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1146),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1206),
.A2(n_1074),
.B(n_1240),
.C(n_1175),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1245),
.B(n_655),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1233),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1315),
.A2(n_1445),
.B1(n_1428),
.B2(n_1446),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1398),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1312),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1303),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1328),
.A2(n_1427),
.B1(n_1426),
.B2(n_1314),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1437),
.B(n_1440),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1401),
.A2(n_1423),
.B(n_1404),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1305),
.Y(n_1473)
);

BUFx2_ASAP7_75t_R g1474 ( 
.A(n_1304),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1375),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1460),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1334),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1459),
.B(n_1464),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1427),
.A2(n_1328),
.B1(n_1333),
.B2(n_1313),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1405),
.B(n_1416),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1342),
.A2(n_1383),
.B1(n_1382),
.B2(n_1443),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1398),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1383),
.A2(n_1382),
.B1(n_1443),
.B2(n_1309),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1395),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1306),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1434),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1319),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1321),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1322),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1329),
.A2(n_1311),
.B1(n_1374),
.B2(n_1320),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1460),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1438),
.A2(n_1353),
.B(n_1338),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1419),
.B(n_1411),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1335),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1323),
.B(n_1444),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1339),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1436),
.Y(n_1498)
);

INVx3_ASAP7_75t_SL g1499 ( 
.A(n_1352),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1458),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1439),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1443),
.A2(n_1309),
.B1(n_1380),
.B2(n_1444),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1429),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1341),
.Y(n_1504)
);

BUFx4f_ASAP7_75t_SL g1505 ( 
.A(n_1400),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1453),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1341),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1408),
.B(n_1308),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1433),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1455),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1356),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1450),
.A2(n_1452),
.B1(n_1348),
.B2(n_1362),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1326),
.B(n_1370),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1331),
.B(n_1420),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1358),
.A2(n_1373),
.B(n_1317),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1345),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1430),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1462),
.Y(n_1518)
);

BUFx2_ASAP7_75t_R g1519 ( 
.A(n_1310),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1389),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1439),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1339),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1341),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1443),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1454),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1368),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1369),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1456),
.A2(n_1330),
.B1(n_1336),
.B2(n_1355),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1439),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1366),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1395),
.Y(n_1531)
);

INVx6_ASAP7_75t_L g1532 ( 
.A(n_1458),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1387),
.B(n_1390),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1325),
.B(n_1347),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1330),
.A2(n_1336),
.B1(n_1452),
.B2(n_1450),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1366),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1344),
.B(n_1349),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1431),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1318),
.A2(n_1409),
.B1(n_1410),
.B2(n_1372),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1386),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1318),
.A2(n_1346),
.B1(n_1441),
.B2(n_1431),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1441),
.A2(n_1424),
.B1(n_1316),
.B2(n_1448),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1332),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1344),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1316),
.A2(n_1451),
.B1(n_1424),
.B2(n_1448),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1386),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1360),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1378),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1451),
.A2(n_1402),
.B1(n_1391),
.B2(n_1447),
.Y(n_1549)
);

INVx3_ASAP7_75t_SL g1550 ( 
.A(n_1352),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1363),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1363),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1421),
.B(n_1406),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1463),
.A2(n_1340),
.B(n_1392),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1380),
.A2(n_1442),
.B1(n_1302),
.B2(n_1324),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1344),
.B(n_1465),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1354),
.A2(n_1397),
.B(n_1392),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1349),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1337),
.B(n_1376),
.Y(n_1559)
);

BUFx2_ASAP7_75t_SL g1560 ( 
.A(n_1400),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1327),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1327),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1350),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1350),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1389),
.B(n_1325),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1447),
.A2(n_1388),
.B1(n_1403),
.B2(n_1385),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1359),
.Y(n_1567)
);

BUFx2_ASAP7_75t_SL g1568 ( 
.A(n_1432),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1447),
.A2(n_1357),
.B1(n_1425),
.B2(n_1347),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1359),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1388),
.A2(n_1403),
.B1(n_1352),
.B2(n_1357),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1425),
.A2(n_1457),
.B1(n_1389),
.B2(n_1384),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1393),
.A2(n_1381),
.B1(n_1395),
.B2(n_1394),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1457),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1384),
.A2(n_1351),
.B1(n_1399),
.B2(n_1393),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1407),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1365),
.A2(n_1351),
.B1(n_1367),
.B2(n_1401),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1339),
.A2(n_1301),
.B1(n_1435),
.B2(n_1378),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1396),
.B(n_1377),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1379),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1371),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1421),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1361),
.B(n_1377),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_R g1584 ( 
.A1(n_1371),
.A2(n_1378),
.B1(n_1435),
.B2(n_1413),
.Y(n_1584)
);

BUFx12f_ASAP7_75t_L g1585 ( 
.A(n_1435),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_SL g1586 ( 
.A(n_1396),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1397),
.A2(n_1367),
.B(n_1413),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1422),
.A2(n_1415),
.B(n_1414),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1361),
.A2(n_1396),
.B1(n_1412),
.B2(n_1418),
.Y(n_1589)
);

CKINVDCx11_ASAP7_75t_R g1590 ( 
.A(n_1379),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1422),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1379),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1417),
.A2(n_1449),
.B(n_1465),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1449),
.A2(n_845),
.B1(n_1328),
.B2(n_1428),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1449),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_SL g1596 ( 
.A1(n_1363),
.A2(n_1175),
.B(n_1348),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_SL g1597 ( 
.A1(n_1363),
.A2(n_1175),
.B(n_1348),
.Y(n_1597)
);

BUFx2_ASAP7_75t_SL g1598 ( 
.A(n_1304),
.Y(n_1598)
);

INVx4_ASAP7_75t_SL g1599 ( 
.A(n_1443),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1439),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1353),
.B(n_1389),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1312),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1314),
.B(n_1437),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1303),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1312),
.Y(n_1605)
);

BUFx12f_ASAP7_75t_L g1606 ( 
.A(n_1375),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1358),
.A2(n_1373),
.B(n_1317),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1343),
.A2(n_1364),
.B(n_1373),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1314),
.B(n_1405),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1314),
.B(n_1405),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1314),
.B(n_1405),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1334),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1460),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1307),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1382),
.B(n_1341),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1315),
.A2(n_1165),
.B(n_988),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1343),
.A2(n_1364),
.B(n_1373),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1312),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1303),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1434),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1315),
.A2(n_1165),
.B1(n_988),
.B2(n_1427),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1305),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1307),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1460),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1328),
.A2(n_845),
.B1(n_1445),
.B2(n_1428),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1312),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_L g1627 ( 
.A(n_1314),
.B(n_1458),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1439),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1398),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1312),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1312),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1307),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1469),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1496),
.B(n_1535),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1485),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1533),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1608),
.A2(n_1617),
.B(n_1557),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1587),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1533),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1576),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1467),
.B(n_1482),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1467),
.B(n_1482),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1554),
.Y(n_1645)
);

CKINVDCx6p67_ASAP7_75t_R g1646 ( 
.A(n_1476),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1603),
.B(n_1512),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1510),
.B(n_1471),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1590),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1530),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1493),
.A2(n_1621),
.B(n_1617),
.Y(n_1651)
);

INVx5_ASAP7_75t_SL g1652 ( 
.A(n_1601),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1536),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1503),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1540),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1546),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1629),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1473),
.B(n_1622),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1629),
.B(n_1609),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1582),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1553),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1553),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1551),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1593),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1552),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1494),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1494),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1588),
.A2(n_1607),
.B(n_1515),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1593),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1538),
.B(n_1509),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1468),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1604),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1543),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1487),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1619),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1489),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1490),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1495),
.Y(n_1679)
);

NAND2x1p5_ASAP7_75t_L g1680 ( 
.A(n_1524),
.B(n_1593),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1498),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1616),
.A2(n_1583),
.B(n_1591),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1547),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1610),
.B(n_1611),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1579),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1590),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1511),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1611),
.B(n_1514),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1602),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1514),
.B(n_1583),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1478),
.B(n_1477),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1605),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1618),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1626),
.B(n_1630),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1526),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1631),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1515),
.A2(n_1607),
.B(n_1589),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1527),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1520),
.B(n_1579),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1591),
.A2(n_1575),
.B(n_1491),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1472),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1565),
.B(n_1579),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1472),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1486),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1472),
.Y(n_1705)
);

CKINVDCx6p67_ASAP7_75t_R g1706 ( 
.A(n_1476),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1528),
.B(n_1516),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1565),
.B(n_1601),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1479),
.A2(n_1517),
.B(n_1518),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1470),
.B(n_1601),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1577),
.B(n_1571),
.Y(n_1711)
);

AO21x1_ASAP7_75t_SL g1712 ( 
.A1(n_1594),
.A2(n_1574),
.B(n_1595),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1625),
.A2(n_1466),
.B1(n_1502),
.B2(n_1481),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1541),
.B(n_1627),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1599),
.B(n_1524),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1483),
.A2(n_1555),
.B1(n_1539),
.B2(n_1519),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1564),
.B(n_1549),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1524),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1534),
.B(n_1506),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1614),
.A2(n_1632),
.B(n_1623),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1534),
.B(n_1529),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1534),
.B(n_1529),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_SL g1723 ( 
.A(n_1474),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1529),
.B(n_1521),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_SL g1725 ( 
.A(n_1581),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1586),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1529),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1529),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1566),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1615),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1615),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1567),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1612),
.B(n_1525),
.Y(n_1733)
);

BUFx12f_ASAP7_75t_L g1734 ( 
.A(n_1486),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1501),
.B(n_1628),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1525),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1561),
.B(n_1563),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1562),
.B(n_1550),
.Y(n_1738)
);

OA21x2_ASAP7_75t_L g1739 ( 
.A1(n_1572),
.A2(n_1569),
.B(n_1592),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1570),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1501),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1500),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1501),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1521),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1521),
.B(n_1600),
.Y(n_1745)
);

AO21x2_ASAP7_75t_L g1746 ( 
.A1(n_1573),
.A2(n_1578),
.B(n_1584),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1600),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1600),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1580),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1628),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1580),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1558),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1504),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1499),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1500),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1558),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1642),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1665),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1649),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1714),
.B(n_1559),
.C(n_1513),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1718),
.Y(n_1762)
);

CKINVDCx6p67_ASAP7_75t_R g1763 ( 
.A(n_1734),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1720),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1718),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1690),
.B(n_1550),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1649),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1690),
.B(n_1499),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1647),
.B(n_1568),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1667),
.B(n_1581),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1667),
.B(n_1542),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1668),
.B(n_1544),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1659),
.B(n_1634),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1691),
.B(n_1606),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1659),
.B(n_1523),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1634),
.B(n_1640),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1640),
.B(n_1523),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1688),
.B(n_1544),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1668),
.B(n_1531),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1688),
.B(n_1548),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1661),
.B(n_1531),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1672),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1636),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1672),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1675),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1682),
.B(n_1548),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1661),
.B(n_1484),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1675),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1682),
.B(n_1558),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1682),
.B(n_1484),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1665),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1658),
.B(n_1654),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1677),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1637),
.B(n_1641),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1637),
.B(n_1641),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1662),
.B(n_1484),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1662),
.B(n_1484),
.Y(n_1797)
);

INVx5_ASAP7_75t_SL g1798 ( 
.A(n_1649),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1677),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1673),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1716),
.A2(n_1620),
.B1(n_1624),
.B2(n_1492),
.C(n_1613),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1678),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1678),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1643),
.B(n_1531),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1643),
.B(n_1531),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1644),
.B(n_1507),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1676),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1683),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1657),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1644),
.B(n_1507),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1649),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1633),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1657),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1633),
.B(n_1532),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1644),
.B(n_1507),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1679),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1674),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1679),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1695),
.B(n_1532),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1681),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1663),
.B(n_1598),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1663),
.B(n_1504),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1644),
.B(n_1702),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1713),
.A2(n_1488),
.B1(n_1545),
.B2(n_1492),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1657),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1736),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1681),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1698),
.B(n_1532),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1684),
.B(n_1537),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1665),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1649),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1671),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1755),
.B(n_1606),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1694),
.B(n_1556),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1734),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1686),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1687),
.B(n_1689),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1670),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1635),
.A2(n_1560),
.B1(n_1620),
.B2(n_1532),
.C(n_1500),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1719),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1692),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1747),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1692),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1773),
.B(n_1651),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1812),
.B(n_1711),
.C(n_1655),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1773),
.B(n_1823),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_SL g1847 ( 
.A(n_1835),
.B(n_1704),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1776),
.B(n_1651),
.Y(n_1848)
);

OAI211xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1783),
.A2(n_1648),
.B(n_1738),
.C(n_1748),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1823),
.B(n_1766),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_L g1851 ( 
.A(n_1769),
.B(n_1711),
.C(n_1655),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1839),
.A2(n_1686),
.B(n_1729),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1762),
.B(n_1742),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1766),
.B(n_1708),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1761),
.B(n_1707),
.C(n_1738),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1800),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1807),
.B(n_1664),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1762),
.B(n_1742),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1824),
.A2(n_1729),
.B1(n_1710),
.B2(n_1746),
.Y(n_1859)
);

NAND3xp33_ASAP7_75t_L g1860 ( 
.A(n_1842),
.B(n_1656),
.C(n_1653),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1808),
.B(n_1664),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1817),
.B(n_1653),
.C(n_1656),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1768),
.B(n_1733),
.Y(n_1863)
);

NAND3xp33_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1650),
.C(n_1666),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_R g1865 ( 
.A(n_1835),
.B(n_1704),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1768),
.B(n_1708),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1824),
.A2(n_1710),
.B1(n_1646),
.B2(n_1706),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1801),
.A2(n_1740),
.B1(n_1650),
.B2(n_1693),
.C(n_1696),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1666),
.C(n_1740),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1771),
.A2(n_1746),
.B1(n_1712),
.B2(n_1709),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1776),
.B(n_1721),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1774),
.A2(n_1686),
.B(n_1838),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1792),
.B(n_1660),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1786),
.B(n_1660),
.C(n_1743),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_R g1875 ( 
.A(n_1763),
.B(n_1723),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_L g1876 ( 
.A1(n_1837),
.A2(n_1696),
.B(n_1693),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1840),
.A2(n_1701),
.B1(n_1705),
.B2(n_1703),
.C(n_1645),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1764),
.A2(n_1669),
.B(n_1638),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1758),
.A2(n_1701),
.B1(n_1705),
.B2(n_1703),
.C(n_1645),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1804),
.B(n_1721),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1786),
.B(n_1741),
.C(n_1743),
.Y(n_1881)
);

NOR2xp67_ASAP7_75t_L g1882 ( 
.A(n_1759),
.B(n_1670),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1821),
.A2(n_1646),
.B1(n_1706),
.B2(n_1725),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1767),
.B(n_1686),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1821),
.A2(n_1686),
.B1(n_1756),
.B2(n_1500),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1826),
.B(n_1645),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1770),
.A2(n_1756),
.B1(n_1652),
.B2(n_1752),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1771),
.A2(n_1746),
.B1(n_1712),
.B2(n_1709),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1837),
.B(n_1639),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1762),
.B(n_1726),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1770),
.A2(n_1670),
.B1(n_1726),
.B2(n_1737),
.C(n_1717),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1763),
.A2(n_1709),
.B1(n_1651),
.B2(n_1717),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1804),
.B(n_1639),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1838),
.A2(n_1715),
.B(n_1754),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_SL g1895 ( 
.A(n_1833),
.B(n_1488),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1822),
.B(n_1741),
.C(n_1744),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1794),
.B(n_1639),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1794),
.B(n_1722),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1814),
.B(n_1749),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1795),
.B(n_1722),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1829),
.A2(n_1652),
.B1(n_1752),
.B2(n_1749),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1805),
.B(n_1727),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1805),
.B(n_1727),
.Y(n_1903)
);

AOI21xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1831),
.A2(n_1780),
.B(n_1777),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1822),
.B(n_1744),
.C(n_1751),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1795),
.B(n_1750),
.Y(n_1906)
);

NAND3xp33_ASAP7_75t_L g1907 ( 
.A(n_1772),
.B(n_1748),
.C(n_1751),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1775),
.B(n_1728),
.Y(n_1908)
);

NOR3xp33_ASAP7_75t_L g1909 ( 
.A(n_1759),
.B(n_1757),
.C(n_1753),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1778),
.B(n_1750),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1775),
.B(n_1728),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1798),
.A2(n_1652),
.B1(n_1749),
.B2(n_1699),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1778),
.B(n_1780),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1790),
.A2(n_1739),
.B1(n_1700),
.B2(n_1737),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1759),
.A2(n_1732),
.B1(n_1680),
.B2(n_1739),
.C(n_1730),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1796),
.B(n_1724),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1777),
.B(n_1735),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1798),
.A2(n_1754),
.B1(n_1757),
.B2(n_1753),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1791),
.A2(n_1830),
.B1(n_1790),
.B2(n_1789),
.C(n_1772),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1796),
.B(n_1724),
.Y(n_1920)
);

NAND3xp33_ASAP7_75t_L g1921 ( 
.A(n_1781),
.B(n_1732),
.C(n_1731),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1797),
.B(n_1735),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1797),
.B(n_1745),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1806),
.B(n_1685),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1809),
.B(n_1813),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1782),
.B(n_1745),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1781),
.B(n_1730),
.C(n_1731),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1848),
.B(n_1791),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1878),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1897),
.B(n_1779),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1848),
.B(n_1791),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1886),
.B(n_1782),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1882),
.B(n_1830),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1844),
.B(n_1846),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1886),
.B(n_1784),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1889),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1844),
.B(n_1809),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1893),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1878),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1876),
.B(n_1784),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1878),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1857),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1893),
.B(n_1785),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1909),
.B(n_1830),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1861),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1862),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1881),
.B(n_1760),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1874),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1856),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1850),
.B(n_1813),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1854),
.B(n_1825),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1860),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1926),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1866),
.B(n_1825),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1906),
.B(n_1779),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1925),
.B(n_1806),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1925),
.B(n_1871),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1916),
.B(n_1810),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1920),
.B(n_1789),
.Y(n_1959)
);

INVx4_ASAP7_75t_L g1960 ( 
.A(n_1875),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1907),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1880),
.B(n_1697),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1908),
.B(n_1697),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1864),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1869),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1873),
.B(n_1787),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1911),
.B(n_1785),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1896),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1902),
.B(n_1788),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1898),
.B(n_1787),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1905),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1890),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1903),
.B(n_1910),
.Y(n_1973)
);

NAND2x1_ASAP7_75t_L g1974 ( 
.A(n_1924),
.B(n_1767),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1900),
.B(n_1788),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1917),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1922),
.B(n_1793),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1877),
.B(n_1793),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1904),
.B(n_1810),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1879),
.B(n_1799),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1915),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1921),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1890),
.B(n_1760),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1919),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1927),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1851),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1863),
.B(n_1815),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1845),
.Y(n_1988)
);

NOR2xp67_ASAP7_75t_L g1989 ( 
.A(n_1894),
.B(n_1767),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1923),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1891),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1913),
.B(n_1799),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1849),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1859),
.A2(n_1798),
.B1(n_1843),
.B2(n_1841),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1853),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1853),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1875),
.B(n_1865),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1858),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1988),
.A2(n_1852),
.B1(n_1859),
.B2(n_1872),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1964),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1986),
.B(n_1802),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1940),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1986),
.B(n_1802),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1934),
.B(n_1863),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1940),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1934),
.B(n_1899),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1964),
.B(n_1855),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1965),
.B(n_1803),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1934),
.B(n_1899),
.Y(n_2009)
);

AOI32xp33_ASAP7_75t_L g2010 ( 
.A1(n_1948),
.A2(n_1870),
.A3(n_1888),
.B1(n_1892),
.B2(n_1868),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1937),
.B(n_1831),
.Y(n_2011)
);

BUFx2_ASAP7_75t_L g2012 ( 
.A(n_1960),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1960),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_SL g2014 ( 
.A(n_1988),
.B(n_1888),
.C(n_1870),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1965),
.B(n_1803),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1960),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1977),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1949),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1977),
.Y(n_2019)
);

AND2x4_ASAP7_75t_L g2020 ( 
.A(n_1989),
.B(n_1811),
.Y(n_2020)
);

NAND2x1p5_ASAP7_75t_L g2021 ( 
.A(n_1960),
.B(n_1811),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1937),
.B(n_1836),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1985),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1975),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1975),
.Y(n_2025)
);

NAND5xp2_ASAP7_75t_L g2026 ( 
.A(n_1952),
.B(n_1847),
.C(n_1895),
.D(n_1892),
.E(n_1865),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1946),
.B(n_1952),
.Y(n_2027)
);

CKINVDCx16_ASAP7_75t_R g2028 ( 
.A(n_1987),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1979),
.B(n_1836),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1979),
.B(n_1987),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1961),
.B(n_1816),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1957),
.B(n_1815),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1942),
.Y(n_2033)
);

O2A1O1Ixp33_ASAP7_75t_SL g2034 ( 
.A1(n_1997),
.A2(n_1883),
.B(n_1858),
.C(n_1475),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1942),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1945),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1946),
.B(n_1816),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1961),
.B(n_1818),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1966),
.B(n_1949),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1985),
.B(n_1475),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1957),
.B(n_1885),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1945),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1992),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1928),
.B(n_1798),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1992),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1989),
.B(n_1884),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1928),
.B(n_1887),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1943),
.B(n_1818),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1968),
.B(n_1820),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1928),
.B(n_1918),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1944),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1992),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1931),
.B(n_1834),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1943),
.B(n_1820),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1968),
.B(n_1971),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_2016),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2008),
.Y(n_2057)
);

NOR2x1p5_ASAP7_75t_L g2058 ( 
.A(n_2016),
.B(n_1974),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2040),
.B(n_1993),
.Y(n_2059)
);

NAND4xp25_ASAP7_75t_L g2060 ( 
.A(n_2027),
.B(n_1971),
.C(n_1993),
.D(n_1948),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2028),
.B(n_1973),
.Y(n_2061)
);

INVx1_ASAP7_75t_SL g2062 ( 
.A(n_2012),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_2046),
.B(n_1947),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2000),
.B(n_1948),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_2023),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2014),
.A2(n_1991),
.B1(n_1981),
.B2(n_1984),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2053),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2023),
.Y(n_2068)
);

NAND2x1_ASAP7_75t_L g2069 ( 
.A(n_2051),
.B(n_1972),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_2013),
.B(n_1944),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2053),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2051),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2039),
.B(n_2007),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2055),
.B(n_1966),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2017),
.B(n_1982),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2013),
.B(n_2016),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2008),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2019),
.B(n_1982),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2024),
.B(n_2025),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2002),
.B(n_1980),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2015),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_2015),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2001),
.Y(n_2083)
);

NAND3xp33_ASAP7_75t_SL g2084 ( 
.A(n_2010),
.B(n_1981),
.C(n_1978),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2043),
.B(n_1930),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2045),
.B(n_2052),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_2004),
.B(n_1944),
.Y(n_2087)
);

O2A1O1Ixp33_ASAP7_75t_L g2088 ( 
.A1(n_1999),
.A2(n_1981),
.B(n_1978),
.C(n_1984),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2001),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2003),
.B(n_1930),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_2021),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2004),
.B(n_2030),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2003),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2037),
.Y(n_2094)
);

OAI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_2026),
.A2(n_1984),
.B1(n_1991),
.B2(n_1994),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2038),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2049),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2005),
.A2(n_1994),
.B1(n_1980),
.B2(n_1867),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2031),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2031),
.B(n_1990),
.Y(n_2100)
);

INVx5_ASAP7_75t_L g2101 ( 
.A(n_2051),
.Y(n_2101)
);

INVxp67_ASAP7_75t_SL g2102 ( 
.A(n_2018),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2033),
.B(n_1932),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_L g2104 ( 
.A(n_2021),
.B(n_1972),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2035),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2041),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2036),
.B(n_1932),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_2046),
.B(n_1947),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2042),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2048),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2057),
.Y(n_2111)
);

NAND2xp33_ASAP7_75t_L g2112 ( 
.A(n_2065),
.B(n_1972),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2077),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2081),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2083),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2061),
.B(n_2030),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2060),
.A2(n_2034),
.B(n_1935),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2089),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2082),
.B(n_2048),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2093),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2099),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2109),
.Y(n_2122)
);

AOI222xp33_ASAP7_75t_L g2123 ( 
.A1(n_2084),
.A2(n_1938),
.B1(n_1935),
.B2(n_1914),
.C1(n_1936),
.C2(n_1939),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2092),
.B(n_2006),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2079),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2082),
.B(n_2054),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2060),
.B(n_2054),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2087),
.B(n_2006),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2073),
.Y(n_2129)
);

OAI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2088),
.A2(n_1938),
.B1(n_1936),
.B2(n_1929),
.C(n_1941),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2087),
.B(n_2009),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2095),
.A2(n_1914),
.B1(n_1929),
.B2(n_1939),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2102),
.B(n_2009),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2068),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_2066),
.A2(n_1929),
.B1(n_1939),
.B2(n_1941),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2106),
.B(n_1976),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2091),
.B(n_2041),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2062),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2091),
.B(n_2070),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2064),
.B(n_1976),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2090),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2074),
.B(n_1953),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2101),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2110),
.Y(n_2144)
);

INVx4_ASAP7_75t_L g2145 ( 
.A(n_2101),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2086),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2064),
.B(n_1976),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_2059),
.A2(n_1941),
.B1(n_1962),
.B2(n_1739),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2075),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2070),
.B(n_2067),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2071),
.B(n_2050),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2101),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_2058),
.B(n_2020),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2138),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_SL g2155 ( 
.A1(n_2143),
.A2(n_2076),
.B(n_2072),
.C(n_2104),
.Y(n_2155)
);

NOR3xp33_ASAP7_75t_L g2156 ( 
.A(n_2130),
.B(n_2129),
.C(n_2127),
.Y(n_2156)
);

OAI32xp33_ASAP7_75t_L g2157 ( 
.A1(n_2127),
.A2(n_2078),
.A3(n_2063),
.B1(n_2108),
.B2(n_2080),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2141),
.B(n_2105),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2122),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2123),
.A2(n_2098),
.B1(n_2080),
.B2(n_2097),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2141),
.B(n_2105),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2125),
.B(n_2062),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2117),
.A2(n_2094),
.B(n_2096),
.C(n_2107),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2122),
.Y(n_2164)
);

INVxp67_ASAP7_75t_L g2165 ( 
.A(n_2134),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2125),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2146),
.Y(n_2167)
);

OAI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_2149),
.A2(n_2142),
.B1(n_2152),
.B2(n_2143),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_2135),
.A2(n_2107),
.B1(n_2103),
.B2(n_2100),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2146),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2128),
.B(n_2056),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2116),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2149),
.B(n_2085),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2111),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2111),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2116),
.B(n_2020),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2113),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_2153),
.B(n_2145),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_2153),
.B(n_2020),
.Y(n_2179)
);

OAI322xp33_ASAP7_75t_L g2180 ( 
.A1(n_2119),
.A2(n_2103),
.A3(n_2069),
.B1(n_1995),
.B2(n_1996),
.C1(n_1998),
.C2(n_1953),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2132),
.A2(n_2050),
.B1(n_2047),
.B2(n_1947),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2133),
.B(n_2119),
.Y(n_2182)
);

OAI32xp33_ASAP7_75t_L g2183 ( 
.A1(n_2145),
.A2(n_2047),
.A3(n_1996),
.B1(n_1998),
.B2(n_1995),
.Y(n_2183)
);

NAND2xp33_ASAP7_75t_R g2184 ( 
.A(n_2154),
.B(n_2143),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2172),
.B(n_2151),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2156),
.A2(n_2148),
.B1(n_2144),
.B2(n_2120),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2176),
.B(n_2128),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2173),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2165),
.B(n_2151),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2165),
.B(n_2124),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2158),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2176),
.B(n_2131),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2158),
.Y(n_2193)
);

NAND2x1_ASAP7_75t_L g2194 ( 
.A(n_2171),
.B(n_2145),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_2168),
.B(n_2153),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_2178),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2182),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2161),
.B(n_2156),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2161),
.B(n_2124),
.Y(n_2199)
);

AOI222xp33_ASAP7_75t_L g2200 ( 
.A1(n_2181),
.A2(n_2144),
.B1(n_2115),
.B2(n_2113),
.C1(n_2114),
.C2(n_2120),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2160),
.B(n_2114),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2166),
.B(n_2115),
.Y(n_2202)
);

INVxp67_ASAP7_75t_L g2203 ( 
.A(n_2162),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2167),
.B(n_2118),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_2170),
.B(n_2145),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2159),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2180),
.A2(n_2121),
.B1(n_2118),
.B2(n_2150),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2198),
.A2(n_2155),
.B(n_2157),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2194),
.B(n_2179),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_2163),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2184),
.B(n_2152),
.C(n_2164),
.Y(n_2211)
);

AOI221x1_ASAP7_75t_L g2212 ( 
.A1(n_2205),
.A2(n_2152),
.B1(n_2177),
.B2(n_2175),
.C(n_2174),
.Y(n_2212)
);

AOI221xp5_ASAP7_75t_L g2213 ( 
.A1(n_2186),
.A2(n_2183),
.B1(n_2169),
.B2(n_2121),
.C(n_2112),
.Y(n_2213)
);

NAND4xp25_ASAP7_75t_SL g2214 ( 
.A(n_2200),
.B(n_2150),
.C(n_2139),
.D(n_2137),
.Y(n_2214)
);

AOI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2186),
.A2(n_2147),
.B1(n_2140),
.B2(n_2126),
.C(n_2139),
.Y(n_2215)
);

NAND5xp2_ASAP7_75t_L g2216 ( 
.A(n_2188),
.B(n_2034),
.C(n_2131),
.D(n_2137),
.E(n_2136),
.Y(n_2216)
);

NAND3xp33_ASAP7_75t_L g2217 ( 
.A(n_2184),
.B(n_2126),
.C(n_2142),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2189),
.Y(n_2218)
);

A2O1A1Ixp33_ASAP7_75t_L g2219 ( 
.A1(n_2201),
.A2(n_2153),
.B(n_1947),
.C(n_1944),
.Y(n_2219)
);

NAND4xp25_ASAP7_75t_SL g2220 ( 
.A(n_2207),
.B(n_2199),
.C(n_2185),
.D(n_2187),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_2195),
.A2(n_2029),
.B(n_1974),
.Y(n_2221)
);

NOR4xp25_ASAP7_75t_L g2222 ( 
.A(n_2196),
.B(n_2029),
.C(n_1931),
.D(n_2011),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2213),
.B(n_2208),
.Y(n_2223)
);

AOI211x1_ASAP7_75t_L g2224 ( 
.A1(n_2220),
.A2(n_2190),
.B(n_2192),
.C(n_2191),
.Y(n_2224)
);

NOR3xp33_ASAP7_75t_L g2225 ( 
.A(n_2210),
.B(n_2203),
.C(n_2193),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2218),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_SL g2227 ( 
.A(n_2209),
.B(n_2205),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2217),
.Y(n_2228)
);

NOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2211),
.B(n_2206),
.Y(n_2229)
);

INVx1_ASAP7_75t_SL g2230 ( 
.A(n_2221),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2212),
.B(n_2207),
.Y(n_2231)
);

AOI211x1_ASAP7_75t_L g2232 ( 
.A1(n_2214),
.A2(n_2204),
.B(n_2202),
.C(n_2022),
.Y(n_2232)
);

NOR2x1_ASAP7_75t_L g2233 ( 
.A(n_2216),
.B(n_2044),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2219),
.A2(n_1884),
.B(n_2022),
.Y(n_2234)
);

AND4x1_ASAP7_75t_L g2235 ( 
.A(n_2222),
.B(n_1505),
.C(n_2044),
.D(n_1522),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_L g2236 ( 
.A(n_2215),
.B(n_1497),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2232),
.B(n_1963),
.Y(n_2237)
);

OAI211xp5_ASAP7_75t_SL g2238 ( 
.A1(n_2223),
.A2(n_2231),
.B(n_2228),
.C(n_2229),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2224),
.B(n_1963),
.Y(n_2239)
);

AND4x1_ASAP7_75t_L g2240 ( 
.A(n_2227),
.B(n_1497),
.C(n_1522),
.D(n_2011),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2230),
.B(n_1976),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2225),
.B(n_2226),
.Y(n_2242)
);

OAI211xp5_ASAP7_75t_L g2243 ( 
.A1(n_2231),
.A2(n_2032),
.B(n_1931),
.C(n_1950),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2233),
.B(n_2032),
.Y(n_2244)
);

AO221x1_ASAP7_75t_L g2245 ( 
.A1(n_2235),
.A2(n_1912),
.B1(n_1953),
.B2(n_1762),
.C(n_1765),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_L g2246 ( 
.A(n_2236),
.B(n_1962),
.C(n_1963),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2242),
.Y(n_2247)
);

INVxp67_ASAP7_75t_SL g2248 ( 
.A(n_2241),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2244),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2238),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2243),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2239),
.B(n_2237),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2246),
.A2(n_2234),
.B1(n_1933),
.B2(n_1990),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2240),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2245),
.A2(n_1962),
.B1(n_1933),
.B2(n_1983),
.Y(n_2255)
);

AND3x4_ASAP7_75t_L g2256 ( 
.A(n_2249),
.B(n_1983),
.C(n_1933),
.Y(n_2256)
);

OA21x2_ASAP7_75t_L g2257 ( 
.A1(n_2250),
.A2(n_1990),
.B(n_1973),
.Y(n_2257)
);

AND2x2_ASAP7_75t_SL g2258 ( 
.A(n_2247),
.B(n_1983),
.Y(n_2258)
);

NAND4xp25_ASAP7_75t_L g2259 ( 
.A(n_2251),
.B(n_1983),
.C(n_1933),
.D(n_1950),
.Y(n_2259)
);

OAI21xp33_ASAP7_75t_L g2260 ( 
.A1(n_2254),
.A2(n_1967),
.B(n_1969),
.Y(n_2260)
);

NAND4xp25_ASAP7_75t_L g2261 ( 
.A(n_2252),
.B(n_1951),
.C(n_1954),
.D(n_1956),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2248),
.B(n_1585),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2258),
.B(n_2253),
.Y(n_2263)
);

NOR3xp33_ASAP7_75t_L g2264 ( 
.A(n_2262),
.B(n_2259),
.C(n_2260),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2257),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2256),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2265),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2263),
.Y(n_2268)
);

NOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2267),
.B(n_2266),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2269),
.B(n_2268),
.Y(n_2270)
);

OAI22xp5_ASAP7_75t_SL g2271 ( 
.A1(n_2269),
.A2(n_2267),
.B1(n_2264),
.B2(n_2253),
.Y(n_2271)
);

OAI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2270),
.A2(n_2255),
.B1(n_2261),
.B2(n_1585),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_2271),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2273),
.A2(n_1973),
.B1(n_1955),
.B2(n_1970),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2272),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2275),
.A2(n_1955),
.B1(n_1970),
.B2(n_1969),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2276),
.A2(n_2274),
.B1(n_1959),
.B2(n_1827),
.Y(n_2277)
);

OAI221xp5_ASAP7_75t_R g2278 ( 
.A1(n_2277),
.A2(n_1951),
.B1(n_1954),
.B2(n_1956),
.C(n_1958),
.Y(n_2278)
);

AOI211xp5_ASAP7_75t_L g2279 ( 
.A1(n_2278),
.A2(n_1901),
.B(n_1762),
.C(n_1765),
.Y(n_2279)
);


endmodule