module fake_jpeg_26390_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_1),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_31),
.B1(n_17),
.B2(n_34),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_33),
.B1(n_30),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_38),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_63),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_73),
.B(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_69),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_40),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_76),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_48),
.B(n_38),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_37),
.B(n_2),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_35),
.B1(n_29),
.B2(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_88),
.Y(n_108)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_26),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_87),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_47),
.B1(n_57),
.B2(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_98),
.B1(n_102),
.B2(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_79),
.B1(n_90),
.B2(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_36),
.C(n_37),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_75),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_57),
.B1(n_41),
.B2(n_37),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_77),
.B(n_25),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_57),
.B1(n_24),
.B2(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_20),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_63),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_20),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_131),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_125),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_64),
.B1(n_74),
.B2(n_68),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_132),
.B1(n_143),
.B2(n_130),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_68),
.B1(n_78),
.B2(n_65),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_128),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_84),
.B(n_80),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_134),
.B(n_116),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_20),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_61),
.B1(n_67),
.B2(n_77),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_135),
.B(n_138),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_24),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_86),
.B1(n_44),
.B2(n_23),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_19),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_19),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_95),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_101),
.B(n_109),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_165),
.B(n_146),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_107),
.A3(n_111),
.B1(n_114),
.B2(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_118),
.B(n_114),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_164),
.B(n_3),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_158),
.B1(n_156),
.B2(n_159),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_118),
.B1(n_119),
.B2(n_112),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_121),
.B1(n_143),
.B2(n_124),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_97),
.B(n_109),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_100),
.A3(n_103),
.B1(n_82),
.B2(n_25),
.C1(n_104),
.C2(n_23),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_97),
.C(n_115),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_131),
.C(n_142),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_189),
.B(n_185),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_170),
.B1(n_148),
.B2(n_155),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_184),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_121),
.B1(n_132),
.B2(n_134),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_186),
.C(n_188),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_138),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_137),
.B1(n_100),
.B2(n_103),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_103),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_104),
.C(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_15),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_147),
.B1(n_169),
.B2(n_170),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_156),
.B1(n_148),
.B2(n_167),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_178),
.B1(n_191),
.B2(n_182),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_151),
.C(n_149),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.C(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_163),
.C(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_163),
.C(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_205),
.B(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_168),
.C(n_147),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_217),
.B(n_219),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_177),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_203),
.B1(n_193),
.B2(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_175),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_172),
.B(n_183),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_220),
.B1(n_190),
.B2(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_222),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_194),
.C(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_192),
.C(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_182),
.B1(n_180),
.B2(n_176),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.C(n_205),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_215),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_208),
.B(n_210),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_3),
.B(n_4),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_223),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_168),
.B1(n_153),
.B2(n_161),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_230),
.B1(n_153),
.B2(n_184),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_239),
.B(n_241),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_222),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_6),
.B(n_7),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_4),
.B(n_5),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_235),
.B(n_231),
.C(n_234),
.D(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_5),
.B(n_6),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_246),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_241),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_10),
.B(n_12),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_12),
.C(n_13),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_250),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_253),
.Y(n_254)
);


endmodule