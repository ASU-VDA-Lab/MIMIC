module fake_jpeg_29828_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_55),
.Y(n_95)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_51),
.Y(n_89)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_17),
.B(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_73),
.Y(n_110)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_66),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_14),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_26),
.B(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_36),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_40),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_25),
.B1(n_40),
.B2(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_100),
.B1(n_119),
.B2(n_121),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_25),
.B1(n_42),
.B2(n_18),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_99),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_39),
.B1(n_20),
.B2(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_125),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_103),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_123),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_56),
.B1(n_76),
.B2(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_34),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_130),
.B(n_136),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_59),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_146),
.Y(n_172)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_138),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_46),
.B1(n_81),
.B2(n_78),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_142),
.B1(n_143),
.B2(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_137),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_24),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_24),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_154),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_46),
.B1(n_75),
.B2(n_74),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_72),
.B1(n_80),
.B2(n_50),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_63),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_58),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g201 ( 
.A(n_148),
.B(n_42),
.C(n_18),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_31),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_104),
.B(n_31),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_SL g157 ( 
.A(n_88),
.B(n_61),
.C(n_53),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_124),
.B1(n_114),
.B2(n_112),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_23),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_48),
.C(n_68),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_91),
.C(n_97),
.Y(n_175)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_118),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_88),
.B1(n_113),
.B2(n_90),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_171),
.A2(n_158),
.B1(n_163),
.B2(n_139),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_175),
.B(n_188),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_134),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_202),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_20),
.B(n_91),
.C(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_132),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_103),
.B(n_82),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_191),
.B(n_137),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_109),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_207),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_82),
.B(n_97),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_193),
.B1(n_158),
.B2(n_149),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_126),
.A2(n_142),
.B1(n_135),
.B2(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_199),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_1),
.C(n_2),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_96),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_151),
.B1(n_145),
.B2(n_166),
.Y(n_218)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_129),
.A2(n_118),
.A3(n_124),
.B1(n_107),
.B2(n_109),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_147),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_96),
.Y(n_207)
);

AO22x2_ASAP7_75t_SL g208 ( 
.A1(n_126),
.A2(n_113),
.B1(n_112),
.B2(n_107),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_168),
.B(n_153),
.C(n_42),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_164),
.B(n_162),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_198),
.B(n_184),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_217),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_173),
.B1(n_192),
.B2(n_189),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_215),
.A2(n_228),
.B1(n_239),
.B2(n_242),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_13),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_199),
.B1(n_200),
.B2(n_195),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_167),
.C(n_155),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_172),
.C(n_169),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_169),
.B(n_127),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_225),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_133),
.C(n_156),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_197),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_198),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_173),
.B1(n_193),
.B2(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_229),
.B1(n_226),
.B2(n_237),
.Y(n_258)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_207),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_183),
.B1(n_195),
.B2(n_182),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_4),
.B(n_6),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_42),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_6),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_170),
.B(n_187),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_1),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_1),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_4),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_252),
.B1(n_257),
.B2(n_260),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_230),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_196),
.B1(n_202),
.B2(n_203),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_255),
.A2(n_259),
.B(n_240),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_229),
.B1(n_219),
.B2(n_216),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_200),
.B1(n_182),
.B2(n_205),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_265),
.B(n_231),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_179),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_279),
.C(n_224),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_275),
.B1(n_233),
.B2(n_225),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_210),
.A2(n_181),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_242),
.B1(n_239),
.B2(n_213),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_277),
.B1(n_223),
.B2(n_220),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_181),
.B1(n_7),
.B2(n_8),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_259),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_6),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_299),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_238),
.B(n_243),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_276),
.B1(n_266),
.B2(n_250),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_288),
.B1(n_298),
.B2(n_266),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_294),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_211),
.B(n_218),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_262),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_277),
.B1(n_268),
.B2(n_247),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_303),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_216),
.B(n_221),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_235),
.C(n_232),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_265),
.C(n_273),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_274),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_273),
.C(n_279),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_256),
.C(n_270),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_292),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_256),
.C(n_270),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_328),
.C(n_304),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_272),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_324),
.B(n_292),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_330),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_286),
.A2(n_248),
.B1(n_252),
.B2(n_260),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_271),
.B1(n_261),
.B2(n_217),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_278),
.C(n_271),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_227),
.B1(n_234),
.B2(n_249),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_332),
.A2(n_350),
.B1(n_312),
.B2(n_326),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_294),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_334),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_298),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_307),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_337),
.B(n_338),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_321),
.B(n_301),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_349),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_280),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_342),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_315),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_303),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_344),
.Y(n_357)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_322),
.Y(n_345)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_290),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_346),
.A2(n_351),
.B(n_319),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_302),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_320),
.C(n_309),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_296),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_324),
.A2(n_295),
.B1(n_287),
.B2(n_300),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_359),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_351),
.A2(n_316),
.B(n_328),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_361),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_350),
.A2(n_316),
.B1(n_319),
.B2(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_331),
.B1(n_323),
.B2(n_314),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_297),
.C(n_284),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.C(n_367),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_283),
.C(n_289),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_347),
.C(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_334),
.C(n_340),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_374),
.C(n_367),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_379),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_333),
.C(n_346),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_348),
.C(n_285),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_375),
.B(n_376),
.Y(n_381)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_291),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_357),
.A2(n_7),
.B(n_10),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_10),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_366),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_370),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_386),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_352),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_356),
.C(n_354),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_387),
.A2(n_370),
.B(n_358),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_352),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_391),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_398),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_SL g396 ( 
.A(n_388),
.B(n_368),
.C(n_363),
.Y(n_396)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_396),
.A2(n_390),
.B(n_383),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_387),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_361),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_400),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_406),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_397),
.C(n_400),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_392),
.A2(n_359),
.B(n_354),
.Y(n_404)
);

NOR3xp33_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_394),
.C(n_395),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g406 ( 
.A(n_396),
.B(n_381),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_408),
.B(n_409),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_405),
.C(n_402),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_411),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_412),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_410),
.C(n_11),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_11),
.Y(n_415)
);


endmodule