module fake_jpeg_24909_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_45),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_22),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_15),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_35),
.B1(n_22),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_30),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_16),
.C(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_25),
.B1(n_21),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_33),
.B1(n_20),
.B2(n_18),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_15),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_32),
.B(n_31),
.C(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_83),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_19),
.B(n_17),
.C(n_31),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_96),
.B(n_65),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_86),
.B1(n_99),
.B2(n_104),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_91),
.B1(n_98),
.B2(n_69),
.Y(n_142)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_94),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_97),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_56),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_32),
.B1(n_31),
.B2(n_28),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_112),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_108),
.Y(n_118)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_70),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_106),
.C(n_90),
.Y(n_131)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_129),
.B(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_53),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_31),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_141),
.C(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_69),
.B1(n_77),
.B2(n_51),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_97),
.B1(n_63),
.B2(n_32),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_78),
.C(n_71),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_145),
.B1(n_80),
.B2(n_92),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_96),
.A2(n_85),
.B1(n_100),
.B2(n_101),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_54),
.C(n_57),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_158),
.Y(n_191)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_153),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_100),
.B(n_107),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_150),
.A2(n_159),
.B(n_167),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_92),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_27),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_101),
.B1(n_92),
.B2(n_104),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_161),
.B1(n_144),
.B2(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_113),
.B(n_108),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_139),
.B(n_27),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_81),
.B1(n_116),
.B2(n_114),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_135),
.C(n_147),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_164),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_121),
.C(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_81),
.C(n_84),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_87),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_119),
.B(n_57),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_168),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_79),
.B(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_0),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_176),
.B(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_89),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_115),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_177),
.B1(n_139),
.B2(n_123),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_0),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_132),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_120),
.A2(n_28),
.B(n_27),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_118),
.A2(n_97),
.B1(n_63),
.B2(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_182),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_0),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_142),
.A3(n_146),
.B1(n_118),
.B2(n_124),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_167),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_128),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_160),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_201),
.B1(n_214),
.B2(n_172),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_0),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_206),
.B(n_209),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_210),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_202),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_197),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_144),
.B1(n_123),
.B2(n_126),
.Y(n_201)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_149),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_27),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_148),
.B(n_1),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_213),
.B(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_155),
.B(n_1),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_157),
.C(n_162),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_227),
.C(n_229),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_180),
.B1(n_184),
.B2(n_209),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_190),
.B(n_209),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_196),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_234),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_208),
.B(n_206),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_189),
.B1(n_215),
.B2(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_230),
.B1(n_237),
.B2(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_240),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_157),
.C(n_150),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_156),
.C(n_153),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_152),
.B1(n_169),
.B2(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_161),
.C(n_166),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_152),
.B1(n_177),
.B2(n_171),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_168),
.C(n_158),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_170),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_180),
.B(n_149),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_200),
.B(n_191),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_180),
.B1(n_174),
.B2(n_14),
.Y(n_242)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NOR4xp25_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_197),
.C(n_198),
.D(n_207),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_250),
.B(n_251),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_222),
.B1(n_239),
.B2(n_229),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_252),
.B1(n_262),
.B2(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_214),
.B1(n_200),
.B2(n_204),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_221),
.C(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_204),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_266),
.B(n_241),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_201),
.B1(n_188),
.B2(n_190),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_211),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_188),
.B1(n_193),
.B2(n_184),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_216),
.B1(n_231),
.B2(n_203),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_209),
.B1(n_185),
.B2(n_213),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_282),
.B(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_217),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_253),
.C(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_285),
.B1(n_266),
.B2(n_261),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_248),
.B(n_228),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_260),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_251),
.A2(n_242),
.B1(n_218),
.B2(n_231),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_283),
.B1(n_245),
.B2(n_263),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_216),
.B(n_185),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_290),
.C(n_296),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_249),
.B1(n_262),
.B2(n_257),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_301),
.B1(n_11),
.B2(n_4),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_291),
.B(n_272),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_259),
.C(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_254),
.C(n_258),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_245),
.C(n_247),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_282),
.C(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_247),
.B1(n_203),
.B2(n_5),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_267),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_273),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_277),
.B1(n_268),
.B2(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_311),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_314),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_281),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_298),
.B(n_296),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_287),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_11),
.Y(n_314)
);

AOI21x1_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_288),
.B(n_301),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_321),
.Y(n_325)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_307),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_3),
.C2(n_9),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_298),
.B1(n_294),
.B2(n_295),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_308),
.B(n_311),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_3),
.B(n_4),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_3),
.B(n_4),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_309),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_327),
.B(n_328),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_304),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_304),
.C(n_314),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_330),
.B(n_319),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_334),
.B(n_331),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_318),
.B(n_7),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_5),
.B(n_8),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_336),
.B(n_325),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_327),
.C(n_9),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);

HAxp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_10),
.CON(n_340),
.SN(n_340)
);


endmodule