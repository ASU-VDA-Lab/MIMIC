module fake_ariane_3159_n_21129 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_21129);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_21129;

wire n_9872;
wire n_9604;
wire n_12407;
wire n_12343;
wire n_20910;
wire n_3152;
wire n_12018;
wire n_6557;
wire n_20947;
wire n_10678;
wire n_2182;
wire n_11999;
wire n_13176;
wire n_12945;
wire n_20136;
wire n_17081;
wire n_9297;
wire n_4403;
wire n_10557;
wire n_19915;
wire n_14456;
wire n_7832;
wire n_8438;
wire n_12244;
wire n_11135;
wire n_1238;
wire n_19533;
wire n_3765;
wire n_19167;
wire n_17213;
wire n_18261;
wire n_15105;
wire n_1096;
wire n_17995;
wire n_12103;
wire n_7922;
wire n_17911;
wire n_2207;
wire n_16181;
wire n_9892;
wire n_6297;
wire n_14334;
wire n_16576;
wire n_16966;
wire n_9263;
wire n_5479;
wire n_6058;
wire n_9886;
wire n_17826;
wire n_10904;
wire n_9096;
wire n_6293;
wire n_13215;
wire n_9665;
wire n_17393;
wire n_14300;
wire n_12233;
wire n_17425;
wire n_10903;
wire n_11906;
wire n_14335;
wire n_13910;
wire n_15347;
wire n_6524;
wire n_146;
wire n_9592;
wire n_1909;
wire n_12260;
wire n_7464;
wire n_19439;
wire n_9683;
wire n_14979;
wire n_4260;
wire n_903;
wire n_7626;
wire n_15874;
wire n_11756;
wire n_7965;
wire n_13636;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_10276;
wire n_13196;
wire n_8460;
wire n_12085;
wire n_14960;
wire n_20861;
wire n_13980;
wire n_14861;
wire n_16646;
wire n_20372;
wire n_12089;
wire n_8734;
wire n_16798;
wire n_18224;
wire n_14592;
wire n_19300;
wire n_559;
wire n_12993;
wire n_16641;
wire n_4741;
wire n_7526;
wire n_21025;
wire n_561;
wire n_10634;
wire n_4273;
wire n_11444;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_786;
wire n_19109;
wire n_5833;
wire n_20492;
wire n_6887;
wire n_9119;
wire n_3552;
wire n_2301;
wire n_15423;
wire n_8504;
wire n_5744;
wire n_5691;
wire n_277;
wire n_7937;
wire n_18827;
wire n_3482;
wire n_18066;
wire n_7490;
wire n_13069;
wire n_5403;
wire n_17391;
wire n_20040;
wire n_20924;
wire n_4268;
wire n_6338;
wire n_587;
wire n_899;
wire n_11856;
wire n_13064;
wire n_334;
wire n_3325;
wire n_661;
wire n_19386;
wire n_11038;
wire n_13991;
wire n_1924;
wire n_17330;
wire n_21038;
wire n_9202;
wire n_11925;
wire n_19274;
wire n_1811;
wire n_6161;
wire n_20554;
wire n_18451;
wire n_12457;
wire n_19819;
wire n_5464;
wire n_10070;
wire n_4476;
wire n_6978;
wire n_579;
wire n_9677;
wire n_149;
wire n_15481;
wire n_20003;
wire n_4000;
wire n_9508;
wire n_13441;
wire n_18294;
wire n_13532;
wire n_2686;
wire n_570;
wire n_11597;
wire n_7874;
wire n_18683;
wire n_8533;
wire n_3511;
wire n_2077;
wire n_19765;
wire n_13912;
wire n_21093;
wire n_1947;
wire n_19473;
wire n_4529;
wire n_7695;
wire n_11611;
wire n_20292;
wire n_12663;
wire n_2800;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_5614;
wire n_5391;
wire n_21081;
wire n_5249;
wire n_3413;
wire n_15098;
wire n_12858;
wire n_19390;
wire n_19927;
wire n_9143;
wire n_5062;
wire n_20264;
wire n_4226;
wire n_10112;
wire n_14150;
wire n_4311;
wire n_5046;
wire n_7607;
wire n_16075;
wire n_13417;
wire n_8442;
wire n_3506;
wire n_1842;
wire n_7397;
wire n_7205;
wire n_555;
wire n_3212;
wire n_11022;
wire n_11025;
wire n_3529;
wire n_11251;
wire n_19364;
wire n_13787;
wire n_5586;
wire n_20095;
wire n_17115;
wire n_11091;
wire n_5056;
wire n_8556;
wire n_5204;
wire n_7307;
wire n_11208;
wire n_4959;
wire n_150;
wire n_7840;
wire n_11487;
wire n_2745;
wire n_8444;
wire n_18453;
wire n_16831;
wire n_19673;
wire n_11745;
wire n_12368;
wire n_19952;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_13054;
wire n_15923;
wire n_3747;
wire n_15957;
wire n_5897;
wire n_19196;
wire n_4894;
wire n_1812;
wire n_15215;
wire n_16402;
wire n_20431;
wire n_7256;
wire n_14458;
wire n_16211;
wire n_3891;
wire n_1623;
wire n_15779;
wire n_7021;
wire n_2435;
wire n_15700;
wire n_20811;
wire n_14375;
wire n_15085;
wire n_542;
wire n_17453;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_14705;
wire n_12944;
wire n_19348;
wire n_7690;
wire n_12973;
wire n_14053;
wire n_6044;
wire n_18530;
wire n_11292;
wire n_15016;
wire n_7966;
wire n_506;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_17645;
wire n_2467;
wire n_14626;
wire n_19495;
wire n_10240;
wire n_4195;
wire n_7007;
wire n_19097;
wire n_21013;
wire n_7230;
wire n_1220;
wire n_7900;
wire n_11203;
wire n_5708;
wire n_14228;
wire n_13801;
wire n_3010;
wire n_2160;
wire n_21096;
wire n_1209;
wire n_9309;
wire n_15480;
wire n_17096;
wire n_10427;
wire n_15527;
wire n_10626;
wire n_17143;
wire n_10138;
wire n_15556;
wire n_9063;
wire n_10532;
wire n_5983;
wire n_21105;
wire n_367;
wire n_15601;
wire n_2632;
wire n_18862;
wire n_12383;
wire n_4314;
wire n_4315;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_11427;
wire n_15739;
wire n_4857;
wire n_8927;
wire n_10398;
wire n_1651;
wire n_6009;
wire n_6382;
wire n_13869;
wire n_9028;
wire n_2677;
wire n_9654;
wire n_10249;
wire n_19135;
wire n_9810;
wire n_7294;
wire n_7414;
wire n_12852;
wire n_9701;
wire n_19632;
wire n_3589;
wire n_8996;
wire n_21051;
wire n_18773;
wire n_17522;
wire n_1943;
wire n_5138;
wire n_16151;
wire n_6048;
wire n_194;
wire n_1163;
wire n_4970;
wire n_16625;
wire n_11070;
wire n_14966;
wire n_8992;
wire n_2373;
wire n_12930;
wire n_20614;
wire n_17005;
wire n_15190;
wire n_12890;
wire n_20915;
wire n_18523;
wire n_6142;
wire n_6119;
wire n_12301;
wire n_17871;
wire n_19209;
wire n_2814;
wire n_11073;
wire n_1439;
wire n_6759;
wire n_3466;
wire n_7092;
wire n_14442;
wire n_4337;
wire n_13095;
wire n_16757;
wire n_15947;
wire n_17129;
wire n_5230;
wire n_17942;
wire n_4486;
wire n_3465;
wire n_12661;
wire n_18580;
wire n_2117;
wire n_20230;
wire n_1053;
wire n_13907;
wire n_9105;
wire n_13085;
wire n_11360;
wire n_5296;
wire n_20469;
wire n_18260;
wire n_16549;
wire n_18903;
wire n_8685;
wire n_1828;
wire n_10997;
wire n_9240;
wire n_19194;
wire n_9212;
wire n_17726;
wire n_17757;
wire n_10602;
wire n_15327;
wire n_17979;
wire n_12088;
wire n_9478;
wire n_19035;
wire n_9742;
wire n_3370;
wire n_21022;
wire n_3949;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_4583;
wire n_8555;
wire n_2118;
wire n_11702;
wire n_636;
wire n_18973;
wire n_1760;
wire n_13596;
wire n_3025;
wire n_14983;
wire n_3051;
wire n_2802;
wire n_13746;
wire n_14550;
wire n_9379;
wire n_18475;
wire n_16186;
wire n_20027;
wire n_2125;
wire n_18207;
wire n_13149;
wire n_4974;
wire n_8245;
wire n_7942;
wire n_4344;
wire n_12186;
wire n_1498;
wire n_16487;
wire n_21035;
wire n_9706;
wire n_957;
wire n_1242;
wire n_14139;
wire n_5596;
wire n_10118;
wire n_8106;
wire n_2217;
wire n_6335;
wire n_11355;
wire n_4460;
wire n_9434;
wire n_1119;
wire n_6229;
wire n_4798;
wire n_10350;
wire n_10654;
wire n_1500;
wire n_616;
wire n_13369;
wire n_5071;
wire n_13653;
wire n_19968;
wire n_3424;
wire n_11584;
wire n_7144;
wire n_3931;
wire n_12256;
wire n_10262;
wire n_11044;
wire n_7316;
wire n_7508;
wire n_19217;
wire n_13785;
wire n_15861;
wire n_1005;
wire n_16741;
wire n_3275;
wire n_5198;
wire n_15463;
wire n_16318;
wire n_2827;
wire n_13943;
wire n_10069;
wire n_16001;
wire n_3085;
wire n_15515;
wire n_12170;
wire n_10791;
wire n_19444;
wire n_12900;
wire n_10553;
wire n_20521;
wire n_20542;
wire n_1219;
wire n_710;
wire n_6631;
wire n_19353;
wire n_7151;
wire n_16736;
wire n_13836;
wire n_12855;
wire n_19967;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4662;
wire n_7075;
wire n_1540;
wire n_20344;
wire n_19855;
wire n_4440;
wire n_17715;
wire n_18105;
wire n_6770;
wire n_14317;
wire n_7611;
wire n_11437;
wire n_7796;
wire n_16663;
wire n_14682;
wire n_832;
wire n_13320;
wire n_12120;
wire n_21001;
wire n_2821;
wire n_10474;
wire n_20304;
wire n_10694;
wire n_20206;
wire n_20988;
wire n_19740;
wire n_20281;
wire n_3531;
wire n_5124;
wire n_655;
wire n_12568;
wire n_8800;
wire n_4652;
wire n_12278;
wire n_17778;
wire n_7655;
wire n_13318;
wire n_3135;
wire n_5719;
wire n_12231;
wire n_7546;
wire n_15343;
wire n_17128;
wire n_14876;
wire n_18259;
wire n_5318;
wire n_5108;
wire n_7407;
wire n_10463;
wire n_11731;
wire n_12097;
wire n_18326;
wire n_17736;
wire n_16579;
wire n_20668;
wire n_13427;
wire n_16339;
wire n_6929;
wire n_19077;
wire n_6012;
wire n_704;
wire n_18401;
wire n_1044;
wire n_4429;
wire n_5435;
wire n_5053;
wire n_16362;
wire n_1243;
wire n_17535;
wire n_16595;
wire n_3486;
wire n_608;
wire n_21066;
wire n_9890;
wire n_2457;
wire n_16272;
wire n_2992;
wire n_16130;
wire n_16164;
wire n_13201;
wire n_11234;
wire n_15375;
wire n_9949;
wire n_1878;
wire n_7076;
wire n_21068;
wire n_10888;
wire n_12714;
wire n_14759;
wire n_5829;
wire n_811;
wire n_20756;
wire n_14193;
wire n_791;
wire n_17172;
wire n_5881;
wire n_17041;
wire n_11895;
wire n_8192;
wire n_16972;
wire n_3450;
wire n_13770;
wire n_10807;
wire n_4050;
wire n_3173;
wire n_14048;
wire n_9546;
wire n_20222;
wire n_6735;
wire n_20723;
wire n_2726;
wire n_9602;
wire n_3266;
wire n_15846;
wire n_19964;
wire n_14816;
wire n_18101;
wire n_2691;
wire n_17611;
wire n_11868;
wire n_12189;
wire n_19506;
wire n_20736;
wire n_16571;
wire n_5419;
wire n_17192;
wire n_13668;
wire n_11571;
wire n_7346;
wire n_17007;
wire n_12069;
wire n_10780;
wire n_18331;
wire n_19616;
wire n_18959;
wire n_13587;
wire n_16559;
wire n_17738;
wire n_15271;
wire n_6904;
wire n_6329;
wire n_17919;
wire n_1488;
wire n_13365;
wire n_1330;
wire n_906;
wire n_6204;
wire n_16627;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_12157;
wire n_13938;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_19365;
wire n_17229;
wire n_15814;
wire n_18381;
wire n_20378;
wire n_11598;
wire n_19984;
wire n_14011;
wire n_21111;
wire n_8645;
wire n_8154;
wire n_5532;
wire n_7311;
wire n_19562;
wire n_6179;
wire n_5441;
wire n_14103;
wire n_7807;
wire n_19085;
wire n_12070;
wire n_3726;
wire n_8480;
wire n_11788;
wire n_14296;
wire n_17305;
wire n_18864;
wire n_20350;
wire n_3560;
wire n_5772;
wire n_6442;
wire n_8241;
wire n_140;
wire n_16249;
wire n_12161;
wire n_18659;
wire n_1009;
wire n_230;
wire n_3548;
wire n_15610;
wire n_6846;
wire n_10343;
wire n_142;
wire n_12238;
wire n_19715;
wire n_8138;
wire n_18027;
wire n_10652;
wire n_15735;
wire n_16479;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_20425;
wire n_15510;
wire n_8235;
wire n_13685;
wire n_1117;
wire n_3321;
wire n_10016;
wire n_6205;
wire n_8349;
wire n_9607;
wire n_7497;
wire n_16201;
wire n_10166;
wire n_2892;
wire n_6939;
wire n_16214;
wire n_2804;
wire n_11240;
wire n_9052;
wire n_426;
wire n_12154;
wire n_8140;
wire n_15276;
wire n_1367;
wire n_14477;
wire n_19424;
wire n_5679;
wire n_15143;
wire n_5141;
wire n_6627;
wire n_19011;
wire n_18623;
wire n_8129;
wire n_1291;
wire n_11156;
wire n_9535;
wire n_13511;
wire n_3987;
wire n_4249;
wire n_19142;
wire n_3160;
wire n_17266;
wire n_14608;
wire n_3223;
wire n_6551;
wire n_20359;
wire n_17591;
wire n_12350;
wire n_7505;
wire n_13993;
wire n_17073;
wire n_19154;
wire n_16545;
wire n_20530;
wire n_17242;
wire n_16668;
wire n_15763;
wire n_13931;
wire n_8934;
wire n_11020;
wire n_7318;
wire n_2613;
wire n_9977;
wire n_13378;
wire n_5667;
wire n_168;
wire n_9555;
wire n_15980;
wire n_17856;
wire n_13618;
wire n_10957;
wire n_3444;
wire n_14952;
wire n_20002;
wire n_1671;
wire n_2343;
wire n_869;
wire n_8221;
wire n_6798;
wire n_14646;
wire n_7895;
wire n_18955;
wire n_16655;
wire n_11339;
wire n_17002;
wire n_8225;
wire n_16721;
wire n_889;
wire n_4355;
wire n_20886;
wire n_17433;
wire n_9651;
wire n_10825;
wire n_2608;
wire n_18360;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_10040;
wire n_6395;
wire n_3243;
wire n_3865;
wire n_1194;
wire n_1647;
wire n_19465;
wire n_14864;
wire n_2459;
wire n_15000;
wire n_8689;
wire n_9629;
wire n_18627;
wire n_14985;
wire n_19166;
wire n_5426;
wire n_13426;
wire n_4093;
wire n_10524;
wire n_4123;
wire n_13799;
wire n_14207;
wire n_19379;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_6502;
wire n_6944;
wire n_18630;
wire n_18274;
wire n_3195;
wire n_13480;
wire n_9349;
wire n_15658;
wire n_11267;
wire n_20334;
wire n_13780;
wire n_10119;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_18569;
wire n_14227;
wire n_17569;
wire n_19231;
wire n_3168;
wire n_17549;
wire n_6075;
wire n_5125;
wire n_12547;
wire n_8928;
wire n_13967;
wire n_18956;
wire n_13014;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_12192;
wire n_16155;
wire n_20656;
wire n_7402;
wire n_6351;
wire n_2073;
wire n_7382;
wire n_10861;
wire n_14729;
wire n_5238;
wire n_750;
wire n_14992;
wire n_19051;
wire n_1612;
wire n_800;
wire n_18025;
wire n_19600;
wire n_5732;
wire n_18914;
wire n_10494;
wire n_724;
wire n_11653;
wire n_2931;
wire n_5556;
wire n_6006;
wire n_10078;
wire n_1589;
wire n_15475;
wire n_3786;
wire n_9995;
wire n_10629;
wire n_19336;
wire n_14165;
wire n_793;
wire n_14192;
wire n_6927;
wire n_13072;
wire n_19550;
wire n_9413;
wire n_4411;
wire n_18638;
wire n_17068;
wire n_4317;
wire n_15713;
wire n_494;
wire n_18549;
wire n_18018;
wire n_3550;
wire n_7956;
wire n_5510;
wire n_4785;
wire n_9775;
wire n_12922;
wire n_13033;
wire n_8580;
wire n_20237;
wire n_12193;
wire n_20383;
wire n_3610;
wire n_3279;
wire n_12243;
wire n_16855;
wire n_18016;
wire n_2923;
wire n_164;
wire n_9305;
wire n_16045;
wire n_5197;
wire n_18147;
wire n_14269;
wire n_7926;
wire n_2394;
wire n_11882;
wire n_14820;
wire n_17247;
wire n_8643;
wire n_15715;
wire n_19247;
wire n_7528;
wire n_20170;
wire n_16107;
wire n_8094;
wire n_2564;
wire n_11695;
wire n_14520;
wire n_13101;
wire n_13723;
wire n_783;
wire n_13556;
wire n_18478;
wire n_1127;
wire n_160;
wire n_15520;
wire n_12356;
wire n_18004;
wire n_5157;
wire n_14654;
wire n_9347;
wire n_5178;
wire n_13350;
wire n_9420;
wire n_12972;
wire n_3105;
wire n_16163;
wire n_1525;
wire n_8477;
wire n_1775;
wire n_12438;
wire n_18821;
wire n_15435;
wire n_14245;
wire n_14254;
wire n_4083;
wire n_12554;
wire n_1272;
wire n_18947;
wire n_18890;
wire n_7506;
wire n_9530;
wire n_10160;
wire n_6809;
wire n_13259;
wire n_6099;
wire n_10849;
wire n_3225;
wire n_244;
wire n_7561;
wire n_18413;
wire n_12860;
wire n_20322;
wire n_15616;
wire n_10282;
wire n_19020;
wire n_19044;
wire n_11393;
wire n_6407;
wire n_3040;
wire n_20204;
wire n_18179;
wire n_445;
wire n_1930;
wire n_1843;
wire n_9713;
wire n_19720;
wire n_2556;
wire n_19292;
wire n_9314;
wire n_12270;
wire n_15325;
wire n_3633;
wire n_857;
wire n_5701;
wire n_20618;
wire n_14949;
wire n_10522;
wire n_17484;
wire n_13348;
wire n_10244;
wire n_10914;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_7773;
wire n_20657;
wire n_1996;
wire n_10980;
wire n_7730;
wire n_20738;
wire n_13265;
wire n_8134;
wire n_18183;
wire n_4690;
wire n_18045;
wire n_9410;
wire n_16285;
wire n_4169;
wire n_8610;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_20553;
wire n_1344;
wire n_435;
wire n_9740;
wire n_9910;
wire n_2139;
wire n_7613;
wire n_15178;
wire n_20328;
wire n_9941;
wire n_9579;
wire n_2740;
wire n_14121;
wire n_15769;
wire n_18333;
wire n_17918;
wire n_20932;
wire n_10938;
wire n_6426;
wire n_4681;
wire n_11956;
wire n_18488;
wire n_9258;
wire n_20099;
wire n_11874;
wire n_5094;
wire n_16096;
wire n_3232;
wire n_3768;
wire n_21024;
wire n_4100;
wire n_20450;
wire n_11822;
wire n_12179;
wire n_19024;
wire n_1409;
wire n_14715;
wire n_5026;
wire n_18304;
wire n_2856;
wire n_18100;
wire n_7679;
wire n_18538;
wire n_20147;
wire n_10811;
wire n_1875;
wire n_10073;
wire n_18044;
wire n_20064;
wire n_5286;
wire n_14779;
wire n_13172;
wire n_19642;
wire n_20226;
wire n_16065;
wire n_15438;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_20913;
wire n_20126;
wire n_4407;
wire n_15080;
wire n_13650;
wire n_21075;
wire n_17696;
wire n_7100;
wire n_7243;
wire n_5243;
wire n_1915;
wire n_11034;
wire n_7415;
wire n_14747;
wire n_15462;
wire n_8795;
wire n_11560;
wire n_9186;
wire n_14054;
wire n_4918;
wire n_5110;
wire n_3659;
wire n_3928;
wire n_20191;
wire n_10500;
wire n_20801;
wire n_10359;
wire n_19999;
wire n_10548;
wire n_2513;
wire n_4408;
wire n_19884;
wire n_15638;
wire n_17505;
wire n_17801;
wire n_860;
wire n_6525;
wire n_5938;
wire n_14270;
wire n_7274;
wire n_17690;
wire n_14859;
wire n_10757;
wire n_8495;
wire n_17895;
wire n_19137;
wire n_17973;
wire n_6132;
wire n_11136;
wire n_18098;
wire n_3071;
wire n_11133;
wire n_14710;
wire n_14781;
wire n_17261;
wire n_6882;
wire n_4624;
wire n_16877;
wire n_4963;
wire n_4205;
wire n_1683;
wire n_15512;
wire n_8600;
wire n_8229;
wire n_415;
wire n_17419;
wire n_2384;
wire n_13579;
wire n_3895;
wire n_1091;
wire n_16079;
wire n_9369;
wire n_13634;
wire n_4338;
wire n_14804;
wire n_15732;
wire n_11804;
wire n_304;
wire n_9076;
wire n_17036;
wire n_5304;
wire n_16416;
wire n_20690;
wire n_2047;
wire n_17903;
wire n_1655;
wire n_3709;
wire n_1146;
wire n_11531;
wire n_12943;
wire n_20227;
wire n_3592;
wire n_15024;
wire n_20679;
wire n_16203;
wire n_14144;
wire n_7454;
wire n_12295;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_11883;
wire n_6931;
wire n_6521;
wire n_6379;
wire n_18431;
wire n_20092;
wire n_6306;
wire n_925;
wire n_12891;
wire n_17862;
wire n_6834;
wire n_2880;
wire n_1001;
wire n_4654;
wire n_13166;
wire n_15695;
wire n_1051;
wire n_10740;
wire n_19107;
wire n_3221;
wire n_17775;
wire n_10062;
wire n_2316;
wire n_8944;
wire n_15265;
wire n_5500;
wire n_9275;
wire n_15955;
wire n_11477;
wire n_5672;
wire n_4016;
wire n_5621;
wire n_9493;
wire n_20855;
wire n_548;
wire n_5966;
wire n_6589;
wire n_10721;
wire n_18468;
wire n_11742;
wire n_17761;
wire n_16452;
wire n_11312;
wire n_1931;
wire n_5559;
wire n_849;
wire n_4655;
wire n_7459;
wire n_7324;
wire n_8205;
wire n_11505;
wire n_20586;
wire n_8975;
wire n_6055;
wire n_1808;
wire n_6348;
wire n_9987;
wire n_20896;
wire n_1704;
wire n_8041;
wire n_20323;
wire n_14327;
wire n_1308;
wire n_11241;
wire n_6144;
wire n_10389;
wire n_1487;
wire n_17108;
wire n_12336;
wire n_9417;
wire n_15534;
wire n_2484;
wire n_20931;
wire n_8076;
wire n_12931;
wire n_1469;
wire n_11066;
wire n_8757;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_9386;
wire n_2500;
wire n_3181;
wire n_13915;
wire n_16645;
wire n_1713;
wire n_7816;
wire n_12119;
wire n_6748;
wire n_11275;
wire n_13589;
wire n_16618;
wire n_11329;
wire n_13189;
wire n_1566;
wire n_2837;
wire n_20018;
wire n_4116;
wire n_10501;
wire n_7269;
wire n_7047;
wire n_16348;
wire n_18839;
wire n_2702;
wire n_16113;
wire n_9176;
wire n_12405;
wire n_3561;
wire n_19056;
wire n_11809;
wire n_10777;
wire n_18900;
wire n_2529;
wire n_3154;
wire n_19784;
wire n_14685;
wire n_19625;
wire n_12780;
wire n_9465;
wire n_13277;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_12662;
wire n_10965;
wire n_11441;
wire n_13503;
wire n_20087;
wire n_4439;
wire n_3382;
wire n_3808;
wire n_17409;
wire n_4660;
wire n_8503;
wire n_15364;
wire n_13287;
wire n_15563;
wire n_2960;
wire n_6807;
wire n_17987;
wire n_13726;
wire n_20508;
wire n_11790;
wire n_402;
wire n_1979;
wire n_6616;
wire n_14621;
wire n_829;
wire n_12190;
wire n_15134;
wire n_11249;
wire n_8707;
wire n_6677;
wire n_5502;
wire n_8931;
wire n_8248;
wire n_14177;
wire n_1283;
wire n_20912;
wire n_13837;
wire n_7302;
wire n_13680;
wire n_9357;
wire n_11911;
wire n_19395;
wire n_8501;
wire n_5706;
wire n_11304;
wire n_2746;
wire n_242;
wire n_13146;
wire n_20621;
wire n_12128;
wire n_11776;
wire n_14544;
wire n_20247;
wire n_9289;
wire n_6443;
wire n_6072;
wire n_15656;
wire n_18454;
wire n_1528;
wire n_9797;
wire n_3315;
wire n_3523;
wire n_17804;
wire n_14440;
wire n_14765;
wire n_9793;
wire n_12017;
wire n_5213;
wire n_3474;
wire n_9514;
wire n_12139;
wire n_11078;
wire n_5620;
wire n_1542;
wire n_4831;
wire n_17831;
wire n_12592;
wire n_11218;
wire n_1851;
wire n_1415;
wire n_10258;
wire n_19378;
wire n_16765;
wire n_4597;
wire n_12791;
wire n_9501;
wire n_16279;
wire n_11775;
wire n_5187;
wire n_18980;
wire n_4147;
wire n_16066;
wire n_10042;
wire n_12162;
wire n_19545;
wire n_6531;
wire n_9481;
wire n_11768;
wire n_19248;
wire n_17633;
wire n_14330;
wire n_20305;
wire n_12960;
wire n_5148;
wire n_18673;
wire n_2867;
wire n_2899;
wire n_18116;
wire n_17765;
wire n_3877;
wire n_14380;
wire n_10754;
wire n_6386;
wire n_2722;
wire n_17246;
wire n_5107;
wire n_18736;
wire n_4680;
wire n_5067;
wire n_11932;
wire n_12485;
wire n_15183;
wire n_15904;
wire n_15113;
wire n_18746;
wire n_1012;
wire n_9748;
wire n_5987;
wire n_2512;
wire n_10851;
wire n_9005;
wire n_12090;
wire n_6642;
wire n_14081;
wire n_19979;
wire n_18920;
wire n_3084;
wire n_6781;
wire n_4593;
wire n_461;
wire n_6509;
wire n_8107;
wire n_6376;
wire n_16610;
wire n_10498;
wire n_18518;
wire n_9947;
wire n_14921;
wire n_10420;
wire n_4498;
wire n_772;
wire n_6741;
wire n_19302;
wire n_10520;
wire n_14839;
wire n_6434;
wire n_5741;
wire n_12583;
wire n_7827;
wire n_676;
wire n_7631;
wire n_8452;
wire n_6690;
wire n_2568;
wire n_2271;
wire n_3485;
wire n_3777;
wire n_9656;
wire n_1585;
wire n_18313;
wire n_12462;
wire n_212;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_11004;
wire n_19101;
wire n_2426;
wire n_6947;
wire n_16329;
wire n_20927;
wire n_9154;
wire n_10937;
wire n_10493;
wire n_21047;
wire n_5574;
wire n_13264;
wire n_18710;
wire n_5877;
wire n_14406;
wire n_912;
wire n_6375;
wire n_460;
wire n_17205;
wire n_17959;
wire n_13294;
wire n_20468;
wire n_10954;
wire n_9788;
wire n_9589;
wire n_17072;
wire n_7855;
wire n_15314;
wire n_8850;
wire n_794;
wire n_18794;
wire n_7886;
wire n_14740;
wire n_18784;
wire n_3306;
wire n_8993;
wire n_11159;
wire n_17906;
wire n_15450;
wire n_20960;
wire n_9946;
wire n_288;
wire n_1292;
wire n_8634;
wire n_11715;
wire n_13625;
wire n_8831;
wire n_14324;
wire n_9979;
wire n_6948;
wire n_13210;
wire n_1610;
wire n_19553;
wire n_11889;
wire n_306;
wire n_2952;
wire n_9007;
wire n_5066;
wire n_19281;
wire n_9260;
wire n_5200;
wire n_15203;
wire n_12365;
wire n_2836;
wire n_2864;
wire n_1717;
wire n_5992;
wire n_8646;
wire n_15782;
wire n_13573;
wire n_17796;
wire n_12518;
wire n_19285;
wire n_19377;
wire n_9752;
wire n_6632;
wire n_2333;
wire n_15041;
wire n_2147;
wire n_6623;
wire n_9395;
wire n_20340;
wire n_17477;
wire n_10294;
wire n_16578;
wire n_1240;
wire n_8031;
wire n_17461;
wire n_425;
wire n_8575;
wire n_20242;
wire n_5097;
wire n_11976;
wire n_3727;
wire n_17025;
wire n_6537;
wire n_17982;
wire n_10969;
wire n_13015;
wire n_15536;
wire n_20467;
wire n_7640;
wire n_3014;
wire n_7912;
wire n_2895;
wire n_4492;
wire n_15284;
wire n_10666;
wire n_19276;
wire n_16420;
wire n_5661;
wire n_17960;
wire n_4975;
wire n_11638;
wire n_16654;
wire n_5306;
wire n_13908;
wire n_11659;
wire n_20770;
wire n_2025;
wire n_8679;
wire n_11948;
wire n_11843;
wire n_16196;
wire n_19057;
wire n_10659;
wire n_11689;
wire n_19402;
wire n_16853;
wire n_9163;
wire n_2495;
wire n_5314;
wire n_14868;
wire n_9322;
wire n_14493;
wire n_10793;
wire n_14491;
wire n_5064;
wire n_6412;
wire n_11108;
wire n_7235;
wire n_16958;
wire n_19790;
wire n_14381;
wire n_13020;
wire n_18492;
wire n_19062;
wire n_15686;
wire n_17874;
wire n_9971;
wire n_2535;
wire n_345;
wire n_17747;
wire n_10976;
wire n_9624;
wire n_10045;
wire n_16761;
wire n_10232;
wire n_8525;
wire n_12166;
wire n_12507;
wire n_776;
wire n_15968;
wire n_6584;
wire n_18474;
wire n_21048;
wire n_6387;
wire n_16384;
wire n_15359;
wire n_19394;
wire n_6470;
wire n_15401;
wire n_14569;
wire n_7383;
wire n_12430;
wire n_4983;
wire n_3185;
wire n_10306;
wire n_12902;
wire n_17014;
wire n_17814;
wire n_17274;
wire n_11337;
wire n_2662;
wire n_18817;
wire n_1231;
wire n_5623;
wire n_19706;
wire n_19789;
wire n_9753;
wire n_5023;
wire n_10931;
wire n_9468;
wire n_7854;
wire n_16179;
wire n_9517;
wire n_7959;
wire n_16502;
wire n_6363;
wire n_15642;
wire n_20317;
wire n_19638;
wire n_15197;
wire n_6811;
wire n_6687;
wire n_18473;
wire n_6037;
wire n_4186;
wire n_19938;
wire n_19416;
wire n_4699;
wire n_17637;
wire n_4096;
wire n_19050;
wire n_12016;
wire n_1570;
wire n_20329;
wire n_10150;
wire n_6722;
wire n_9780;
wire n_18405;
wire n_19228;
wire n_5153;
wire n_18995;
wire n_17442;
wire n_4713;
wire n_17806;
wire n_19547;
wire n_16111;
wire n_18387;
wire n_18790;
wire n_10187;
wire n_17341;
wire n_7080;
wire n_8695;
wire n_7436;
wire n_8571;
wire n_7020;
wire n_5935;
wire n_13302;
wire n_5967;
wire n_5934;
wire n_1899;
wire n_16605;
wire n_17990;
wire n_3508;
wire n_18171;
wire n_17488;
wire n_4129;
wire n_18524;
wire n_11114;
wire n_16648;
wire n_10479;
wire n_7978;
wire n_5727;
wire n_3599;
wire n_20010;
wire n_5646;
wire n_16209;
wire n_7694;
wire n_5711;
wire n_8771;
wire n_6254;
wire n_20537;
wire n_3401;
wire n_10360;
wire n_14891;
wire n_16136;
wire n_9074;
wire n_12975;
wire n_19885;
wire n_11556;
wire n_7465;
wire n_19585;
wire n_5470;
wire n_1092;
wire n_2225;
wire n_16330;
wire n_1963;
wire n_16011;
wire n_9300;
wire n_14489;
wire n_13619;
wire n_18785;
wire n_2218;
wire n_8352;
wire n_7760;
wire n_21040;
wire n_12977;
wire n_19040;
wire n_2741;
wire n_2714;
wire n_21127;
wire n_13177;
wire n_17908;
wire n_10953;
wire n_15285;
wire n_6587;
wire n_6688;
wire n_19882;
wire n_8986;
wire n_17324;
wire n_20680;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_11342;
wire n_9114;
wire n_1055;
wire n_8396;
wire n_8514;
wire n_13482;
wire n_8151;
wire n_14688;
wire n_16242;
wire n_16862;
wire n_15579;
wire n_3568;
wire n_19433;
wire n_6220;
wire n_15439;
wire n_10598;
wire n_7882;
wire n_16818;
wire n_2470;
wire n_11750;
wire n_3551;
wire n_417;
wire n_13412;
wire n_1708;
wire n_11338;
wire n_18220;
wire n_5650;
wire n_5189;
wire n_15342;
wire n_8070;
wire n_15595;
wire n_10064;
wire n_14863;
wire n_3985;
wire n_15742;
wire n_6439;
wire n_148;
wire n_17983;
wire n_1741;
wire n_14247;
wire n_13075;
wire n_20874;
wire n_7902;
wire n_11408;
wire n_20364;
wire n_742;
wire n_5160;
wire n_12971;
wire n_769;
wire n_15193;
wire n_12674;
wire n_20085;
wire n_2366;
wire n_1753;
wire n_14419;
wire n_10800;
wire n_13038;
wire n_17708;
wire n_17789;
wire n_6478;
wire n_298;
wire n_5874;
wire n_19845;
wire n_19889;
wire n_3956;
wire n_17104;
wire n_4081;
wire n_20603;
wire n_606;
wire n_17101;
wire n_15490;
wire n_19073;
wire n_509;
wire n_1747;
wire n_18606;
wire n_14312;
wire n_12346;
wire n_5622;
wire n_14110;
wire n_20004;
wire n_8618;
wire n_18552;
wire n_16568;
wire n_4069;
wire n_3582;
wire n_15558;
wire n_3993;
wire n_4811;
wire n_2696;
wire n_17510;
wire n_4779;
wire n_5910;
wire n_9616;
wire n_10153;
wire n_1400;
wire n_7862;
wire n_17665;
wire n_18753;
wire n_7565;
wire n_7410;
wire n_1527;
wire n_7721;
wire n_9209;
wire n_16987;
wire n_2831;
wire n_10585;
wire n_5568;
wire n_14996;
wire n_5941;
wire n_11300;
wire n_14294;
wire n_13425;
wire n_17652;
wire n_15251;
wire n_17581;
wire n_6604;
wire n_19335;
wire n_3302;
wire n_18987;
wire n_2486;
wire n_9086;
wire n_1897;
wire n_6999;
wire n_7539;
wire n_17314;
wire n_6440;
wire n_4977;
wire n_14417;
wire n_11072;
wire n_7608;
wire n_15084;
wire n_16344;
wire n_2912;
wire n_14650;
wire n_18872;
wire n_595;
wire n_14789;
wire n_17975;
wire n_17392;
wire n_6784;
wire n_1757;
wire n_20652;
wire n_17860;
wire n_11421;
wire n_2090;
wire n_295;
wire n_10310;
wire n_4200;
wire n_5222;
wire n_6165;
wire n_10133;
wire n_12793;
wire n_11989;
wire n_21083;
wire n_1281;
wire n_2574;
wire n_1856;
wire n_18301;
wire n_13392;
wire n_12865;
wire n_4604;
wire n_20055;
wire n_1293;
wire n_18006;
wire n_961;
wire n_9261;
wire n_19346;
wire n_12285;
wire n_726;
wire n_7348;
wire n_14894;
wire n_12478;
wire n_3857;
wire n_19110;
wire n_9375;
wire n_13059;
wire n_19835;
wire n_18056;
wire n_2730;
wire n_9448;
wire n_13199;
wire n_806;
wire n_21041;
wire n_15654;
wire n_15531;
wire n_12369;
wire n_11118;
wire n_18073;
wire n_11844;
wire n_2064;
wire n_9271;
wire n_5663;
wire n_15332;
wire n_7933;
wire n_16704;
wire n_349;
wire n_16735;
wire n_12520;
wire n_4343;
wire n_15479;
wire n_5389;
wire n_2986;
wire n_19483;
wire n_15186;
wire n_15461;
wire n_3591;
wire n_20157;
wire n_13422;
wire n_3317;
wire n_19202;
wire n_13042;
wire n_11884;
wire n_15664;
wire n_14860;
wire n_4835;
wire n_554;
wire n_4420;
wire n_14513;
wire n_2244;
wire n_15011;
wire n_4742;
wire n_12605;
wire n_5038;
wire n_14830;
wire n_9850;
wire n_5766;
wire n_14223;
wire n_13234;
wire n_594;
wire n_10970;
wire n_12651;
wire n_13829;
wire n_2247;
wire n_1269;
wire n_16940;
wire n_14880;
wire n_12638;
wire n_21004;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_18686;
wire n_10148;
wire n_7939;
wire n_17286;
wire n_14040;
wire n_3982;
wire n_14361;
wire n_3647;
wire n_17872;
wire n_3973;
wire n_8052;
wire n_8733;
wire n_17507;
wire n_12815;
wire n_6700;
wire n_20361;
wire n_10830;
wire n_9196;
wire n_19490;
wire n_1103;
wire n_5594;
wire n_16530;
wire n_10086;
wire n_9029;
wire n_562;
wire n_7580;
wire n_19368;
wire n_7340;
wire n_8080;
wire n_10279;
wire n_7303;
wire n_914;
wire n_689;
wire n_6139;
wire n_7568;
wire n_20299;
wire n_20592;
wire n_7387;
wire n_13293;
wire n_17913;
wire n_4011;
wire n_21107;
wire n_19571;
wire n_3906;
wire n_3011;
wire n_17712;
wire n_497;
wire n_11645;
wire n_12199;
wire n_6333;
wire n_20642;
wire n_15538;
wire n_12584;
wire n_455;
wire n_18275;
wire n_4816;
wire n_4091;
wire n_10910;
wire n_1417;
wire n_9733;
wire n_3096;
wire n_7207;
wire n_8827;
wire n_4166;
wire n_16754;
wire n_18676;
wire n_15741;
wire n_16513;
wire n_685;
wire n_16864;
wire n_4061;
wire n_14203;
wire n_11504;
wire n_15146;
wire n_11587;
wire n_17993;
wire n_16543;
wire n_20059;
wire n_18398;
wire n_10865;
wire n_8171;
wire n_16812;
wire n_16932;
wire n_9877;
wire n_14578;
wire n_12969;
wire n_17463;
wire n_2396;
wire n_14222;
wire n_12607;
wire n_1559;
wire n_13695;
wire n_7633;
wire n_10246;
wire n_4684;
wire n_10439;
wire n_743;
wire n_1546;
wire n_5279;
wire n_18155;
wire n_962;
wire n_20608;
wire n_7768;
wire n_16947;
wire n_2196;
wire n_12475;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_14643;
wire n_12027;
wire n_14986;
wire n_5232;
wire n_16750;
wire n_1193;
wire n_11405;
wire n_11028;
wire n_6003;
wire n_8133;
wire n_18075;
wire n_2007;
wire n_17080;
wire n_6636;
wire n_9525;
wire n_1158;
wire n_11625;
wire n_12565;
wire n_18014;
wire n_3481;
wire n_7401;
wire n_10735;
wire n_20246;
wire n_6020;
wire n_18893;
wire n_14908;
wire n_14568;
wire n_12561;
wire n_20291;
wire n_9739;
wire n_6785;
wire n_17882;
wire n_17478;
wire n_14871;
wire n_2887;
wire n_4735;
wire n_18555;
wire n_5170;
wire n_5608;
wire n_11739;
wire n_9148;
wire n_10858;
wire n_10736;
wire n_9958;
wire n_2455;
wire n_827;
wire n_3437;
wire n_9323;
wire n_7522;
wire n_7188;
wire n_8088;
wire n_9155;
wire n_8662;
wire n_11291;
wire n_16286;
wire n_17762;
wire n_13566;
wire n_11425;
wire n_19623;
wire n_16470;
wire n_751;
wire n_11890;
wire n_13621;
wire n_5182;
wire n_1221;
wire n_8663;
wire n_10928;
wire n_16956;
wire n_19032;
wire n_6618;
wire n_16195;
wire n_1579;
wire n_18757;
wire n_2014;
wire n_20146;
wire n_2974;
wire n_12461;
wire n_923;
wire n_3969;
wire n_6873;
wire n_18122;
wire n_8118;
wire n_20669;
wire n_7101;
wire n_14191;
wire n_14841;
wire n_6063;
wire n_16245;
wire n_18854;
wire n_7578;
wire n_20856;
wire n_14146;
wire n_19561;
wire n_856;
wire n_8982;
wire n_16656;
wire n_6993;
wire n_9745;
wire n_14288;
wire n_17373;
wire n_508;
wire n_3706;
wire n_1858;
wire n_16351;
wire n_15733;
wire n_1361;
wire n_8381;
wire n_18661;
wire n_8835;
wire n_14553;
wire n_15258;
wire n_6558;
wire n_1411;
wire n_1359;
wire n_9108;
wire n_9907;
wire n_10959;
wire n_3536;
wire n_7263;
wire n_12067;
wire n_20730;
wire n_1317;
wire n_11040;
wire n_20439;
wire n_20124;
wire n_12870;
wire n_3594;
wire n_5383;
wire n_17824;
wire n_7245;
wire n_7310;
wire n_17415;
wire n_5690;
wire n_11332;
wire n_1980;
wire n_18650;
wire n_19151;
wire n_17223;
wire n_13279;
wire n_2604;
wire n_9852;
wire n_10881;
wire n_14049;
wire n_11943;
wire n_12933;
wire n_10544;
wire n_13895;
wire n_14403;
wire n_15899;
wire n_12131;
wire n_6082;
wire n_19581;
wire n_2817;
wire n_20954;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_19484;
wire n_15985;
wire n_16634;
wire n_12399;
wire n_19305;
wire n_7738;
wire n_14787;
wire n_2344;
wire n_8838;
wire n_7609;
wire n_3122;
wire n_6548;
wire n_8607;
wire n_20763;
wire n_14487;
wire n_14615;
wire n_2787;
wire n_10032;
wire n_7282;
wire n_8551;
wire n_16552;
wire n_20983;
wire n_2770;
wire n_18608;
wire n_9248;
wire n_19797;
wire n_5579;
wire n_4167;
wire n_7170;
wire n_11872;
wire n_6674;
wire n_13669;
wire n_12710;
wire n_7489;
wire n_9056;
wire n_9106;
wire n_18344;
wire n_17972;
wire n_14496;
wire n_7281;
wire n_12920;
wire n_4199;
wire n_18930;
wire n_16451;
wire n_11220;
wire n_20982;
wire n_16398;
wire n_7833;
wire n_20658;
wire n_3829;
wire n_5057;
wire n_6196;
wire n_5839;
wire n_2469;
wire n_11551;
wire n_20681;
wire n_3546;
wire n_17720;
wire n_10025;
wire n_16053;
wire n_3068;
wire n_17805;
wire n_19580;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_9786;
wire n_10833;
wire n_10685;
wire n_567;
wire n_20108;
wire n_13611;
wire n_13178;
wire n_20413;
wire n_5487;
wire n_5649;
wire n_16016;
wire n_831;
wire n_18940;
wire n_3970;
wire n_20454;
wire n_18226;
wire n_15617;
wire n_3218;
wire n_6954;
wire n_17677;
wire n_6450;
wire n_6995;
wire n_2447;
wire n_13009;
wire n_4193;
wire n_6347;
wire n_671;
wire n_8387;
wire n_17179;
wire n_11716;
wire n_8105;
wire n_13485;
wire n_6698;
wire n_18680;
wire n_4392;
wire n_17077;
wire n_498;
wire n_12415;
wire n_20489;
wire n_3966;
wire n_4397;
wire n_13273;
wire n_17898;
wire n_4803;
wire n_10155;
wire n_11367;
wire n_6743;
wire n_11418;
wire n_2852;
wire n_8597;
wire n_20128;
wire n_6330;
wire n_18368;
wire n_7045;
wire n_11576;
wire n_175;
wire n_8534;
wire n_21006;
wire n_15046;
wire n_9210;
wire n_17891;
wire n_8655;
wire n_4893;
wire n_13894;
wire n_2240;
wire n_4258;
wire n_14695;
wire n_14455;
wire n_2917;
wire n_20017;
wire n_5033;
wire n_11123;
wire n_14414;
wire n_10248;
wire n_17921;
wire n_11733;
wire n_12915;
wire n_1410;
wire n_20865;
wire n_9756;
wire n_1223;
wire n_572;
wire n_10877;
wire n_15954;
wire n_8879;
wire n_4767;
wire n_17542;
wire n_448;
wire n_9700;
wire n_11503;
wire n_6895;
wire n_8335;
wire n_16607;
wire n_4468;
wire n_3848;
wire n_7400;
wire n_17607;
wire n_16014;
wire n_19650;
wire n_20570;
wire n_4885;
wire n_7475;
wire n_3674;
wire n_716;
wire n_18470;
wire n_14001;
wire n_933;
wire n_5534;
wire n_1821;
wire n_16462;
wire n_12220;
wire n_3910;
wire n_492;
wire n_12375;
wire n_13333;
wire n_20745;
wire n_2995;
wire n_8462;
wire n_3228;
wire n_10651;
wire n_17669;
wire n_21074;
wire n_12809;
wire n_6869;
wire n_4761;
wire n_7672;
wire n_10770;
wire n_6137;
wire n_9467;
wire n_12043;
wire n_3088;
wire n_5254;
wire n_10393;
wire n_2761;
wire n_20946;
wire n_4520;
wire n_13355;
wire n_15639;
wire n_12504;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_6885;
wire n_8727;
wire n_8482;
wire n_6120;
wire n_3557;
wire n_20702;
wire n_1598;
wire n_15194;
wire n_12836;
wire n_17264;
wire n_18654;
wire n_15419;
wire n_10094;
wire n_19530;
wire n_11328;
wire n_17191;
wire n_5438;
wire n_9167;
wire n_15845;
wire n_7954;
wire n_6530;
wire n_4149;
wire n_1827;
wire n_6135;
wire n_246;
wire n_14359;
wire n_10623;
wire n_14786;
wire n_2361;
wire n_3505;
wire n_21029;
wire n_8365;
wire n_20357;
wire n_15973;
wire n_2239;
wire n_16466;
wire n_6942;
wire n_14108;
wire n_17236;
wire n_6892;
wire n_7357;
wire n_9290;
wire n_6782;
wire n_2464;
wire n_3697;
wire n_17514;
wire n_15319;
wire n_17597;
wire n_19917;
wire n_13340;
wire n_7229;
wire n_20928;
wire n_7336;
wire n_17540;
wire n_20511;
wire n_6598;
wire n_10105;
wire n_5919;
wire n_18414;
wire n_8346;
wire n_5012;
wire n_6614;
wire n_11781;
wire n_13310;
wire n_14548;
wire n_14169;
wire n_2517;
wire n_4696;
wire n_9113;
wire n_7493;
wire n_20256;
wire n_2590;
wire n_11140;
wire n_5823;
wire n_15174;
wire n_6989;
wire n_16836;
wire n_8237;
wire n_6299;
wire n_9813;
wire n_19622;
wire n_17592;
wire n_14527;
wire n_13833;
wire n_9394;
wire n_1069;
wire n_2037;
wire n_16213;
wire n_573;
wire n_11082;
wire n_9663;
wire n_7901;
wire n_20067;
wire n_10146;
wire n_913;
wire n_11949;
wire n_19574;
wire n_4834;
wire n_9994;
wire n_15095;
wire n_17739;
wire n_18563;
wire n_4692;
wire n_15153;
wire n_11693;
wire n_2559;
wire n_15717;
wire n_15670;
wire n_8946;
wire n_18447;
wire n_8055;
wire n_5870;
wire n_6233;
wire n_10918;
wire n_4299;
wire n_20301;
wire n_14879;
wire n_20174;
wire n_14597;
wire n_525;
wire n_19463;
wire n_2243;
wire n_13247;
wire n_16720;
wire n_2694;
wire n_6356;
wire n_13391;
wire n_8998;
wire n_4965;
wire n_7601;
wire n_17965;
wire n_11046;
wire n_15529;
wire n_15296;
wire n_11224;
wire n_2006;
wire n_17487;
wire n_12223;
wire n_16469;
wire n_7147;
wire n_8161;
wire n_11101;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_16041;
wire n_18561;
wire n_12378;
wire n_9211;
wire n_6032;
wire n_3435;
wire n_12794;
wire n_4897;
wire n_12436;
wire n_4674;
wire n_15724;
wire n_568;
wire n_4796;
wire n_10975;
wire n_2750;
wire n_11950;
wire n_17039;
wire n_17587;
wire n_8747;
wire n_7617;
wire n_19663;
wire n_16566;
wire n_14652;
wire n_7700;
wire n_20776;
wire n_11709;
wire n_18299;
wire n_20817;
wire n_16222;
wire n_20404;
wire n_10365;
wire n_10778;
wire n_4625;
wire n_7098;
wire n_14668;
wire n_20884;
wire n_16334;
wire n_5070;
wire n_13105;
wire n_4148;
wire n_5575;
wire n_7661;
wire n_16631;
wire n_17054;
wire n_13766;
wire n_13525;
wire n_4590;
wire n_13081;
wire n_10378;
wire n_1888;
wire n_11563;
wire n_19954;
wire n_1425;
wire n_19136;
wire n_18062;
wire n_557;
wire n_7323;
wire n_5048;
wire n_11565;
wire n_17325;
wire n_13257;
wire n_19389;
wire n_5363;
wire n_11164;
wire n_12633;
wire n_18228;
wire n_5665;
wire n_16806;
wire n_20326;
wire n_11414;
wire n_18288;
wire n_10330;
wire n_15136;
wire n_19443;
wire n_21058;
wire n_6394;
wire n_14370;
wire n_7929;
wire n_16456;
wire n_486;
wire n_18141;
wire n_11319;
wire n_9306;
wire n_4353;
wire n_2201;
wire n_10442;
wire n_13865;
wire n_10962;
wire n_10022;
wire n_13973;
wire n_4124;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_10127;
wire n_3596;
wire n_11128;
wire n_9332;
wire n_12262;
wire n_8043;
wire n_8159;
wire n_4608;
wire n_9294;
wire n_17769;
wire n_12235;
wire n_10375;
wire n_1977;
wire n_2650;
wire n_20011;
wire n_4184;
wire n_2391;
wire n_6343;
wire n_12406;
wire n_15213;
wire n_17543;
wire n_3883;
wire n_19792;
wire n_4032;
wire n_5736;
wire n_18161;
wire n_6029;
wire n_4117;
wire n_300;
wire n_12229;
wire n_19448;
wire n_14264;
wire n_3634;
wire n_6697;
wire n_11262;
wire n_16121;
wire n_11110;
wire n_13084;
wire n_14785;
wire n_5341;
wire n_2575;
wire n_13470;
wire n_12245;
wire n_2942;
wire n_15430;
wire n_1771;
wire n_14394;
wire n_6715;
wire n_3164;
wire n_17452;
wire n_2043;
wire n_6771;
wire n_12376;
wire n_4815;
wire n_5639;
wire n_10991;
wire n_11945;
wire n_11769;
wire n_17520;
wire n_12720;
wire n_209;
wire n_5503;
wire n_18264;
wire n_7718;
wire n_19724;
wire n_12708;
wire n_16934;
wire n_503;
wire n_12387;
wire n_13705;
wire n_9081;
wire n_8717;
wire n_9198;
wire n_10571;
wire n_4774;
wire n_4108;
wire n_20619;
wire n_17106;
wire n_17859;
wire n_14002;
wire n_19688;
wire n_9488;
wire n_18038;
wire n_4394;
wire n_15850;
wire n_6444;
wire n_8073;
wire n_17177;
wire n_20271;
wire n_9526;
wire n_4220;
wire n_577;
wire n_9962;
wire n_20593;
wire n_15869;
wire n_19980;
wire n_1468;
wire n_9667;
wire n_18503;
wire n_5166;
wire n_11256;
wire n_19237;
wire n_14018;
wire n_14935;
wire n_17287;
wire n_3624;
wire n_6725;
wire n_1182;
wire n_4594;
wire n_21099;
wire n_14877;
wire n_8447;
wire n_20683;
wire n_10897;
wire n_6913;
wire n_513;
wire n_15804;
wire n_15959;
wire n_10617;
wire n_14438;
wire n_7853;
wire n_9796;
wire n_5770;
wire n_8756;
wire n_2628;
wire n_16125;
wire n_20980;
wire n_1083;
wire n_12831;
wire n_8809;
wire n_16824;
wire n_11815;
wire n_17800;
wire n_18096;
wire n_15135;
wire n_18440;
wire n_16512;
wire n_5008;
wire n_9077;
wire n_12872;
wire n_15879;
wire n_3871;
wire n_19447;
wire n_15644;
wire n_17243;
wire n_6148;
wire n_8255;
wire n_990;
wire n_8216;
wire n_8693;
wire n_16509;
wire n_6522;
wire n_19250;
wire n_16570;
wire n_5582;
wire n_14348;
wire n_7880;
wire n_909;
wire n_8149;
wire n_10067;
wire n_18740;
wire n_10698;
wire n_964;
wire n_7342;
wire n_18835;
wire n_20851;
wire n_7810;
wire n_10260;
wire n_12370;
wire n_19934;
wire n_7114;
wire n_14813;
wire n_5862;
wire n_18443;
wire n_2253;
wire n_11550;
wire n_15965;
wire n_5886;
wire n_9451;
wire n_8479;
wire n_6783;
wire n_14524;
wire n_20774;
wire n_20274;
wire n_16990;
wire n_3673;
wire n_9710;
wire n_12634;
wire n_15896;
wire n_14287;
wire n_5285;
wire n_14052;
wire n_14216;
wire n_1234;
wire n_3936;
wire n_17526;
wire n_17766;
wire n_5162;
wire n_14925;
wire n_5442;
wire n_5802;
wire n_20015;
wire n_14475;
wire n_7858;
wire n_17109;
wire n_20327;
wire n_13699;
wire n_1095;
wire n_6078;
wire n_14122;
wire n_5630;
wire n_18534;
wire n_9452;
wire n_3869;
wire n_13675;
wire n_18428;
wire n_14977;
wire n_6815;
wire n_15275;
wire n_1387;
wire n_19491;
wire n_16981;
wire n_5054;
wire n_3171;
wire n_17998;
wire n_14080;
wire n_4751;
wire n_13814;
wire n_10381;
wire n_2490;
wire n_10554;
wire n_9057;
wire n_3300;
wire n_20188;
wire n_17295;
wire n_7174;
wire n_17751;
wire n_18432;
wire n_19418;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_15766;
wire n_4362;
wire n_15554;
wire n_3946;
wire n_2640;
wire n_4634;
wire n_4089;
wire n_1173;
wire n_18438;
wire n_11508;
wire n_20149;
wire n_7662;
wire n_11138;
wire n_19811;
wire n_14912;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_13585;
wire n_1648;
wire n_8137;
wire n_10841;
wire n_13142;
wire n_3863;
wire n_12642;
wire n_2327;
wire n_3882;
wire n_13974;
wire n_18508;
wire n_3916;
wire n_2437;
wire n_14070;
wire n_14909;
wire n_16004;
wire n_15294;
wire n_20671;
wire n_16660;
wire n_405;
wire n_10719;
wire n_17207;
wire n_12959;
wire n_7984;
wire n_15447;
wire n_481;
wire n_12919;
wire n_19603;
wire n_2308;
wire n_1939;
wire n_15379;
wire n_19427;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_12314;
wire n_20607;
wire n_8091;
wire n_1798;
wire n_19338;
wire n_1608;
wire n_5761;
wire n_18252;
wire n_547;
wire n_439;
wire n_20617;
wire n_3318;
wire n_7232;
wire n_13824;
wire n_9482;
wire n_15570;
wire n_6957;
wire n_20917;
wire n_5074;
wire n_21076;
wire n_3939;
wire n_590;
wire n_3569;
wire n_17910;
wire n_18130;
wire n_15226;
wire n_15927;
wire n_18579;
wire n_7422;
wire n_9785;
wire n_427;
wire n_21079;
wire n_9195;
wire n_8322;
wire n_15623;
wire n_6591;
wire n_8987;
wire n_13454;
wire n_3653;
wire n_9280;
wire n_19100;
wire n_7621;
wire n_13958;
wire n_18255;
wire n_163;
wire n_19692;
wire n_10373;
wire n_7158;
wire n_11173;
wire n_314;
wire n_21049;
wire n_7500;
wire n_1120;
wire n_4084;
wire n_9687;
wire n_7985;
wire n_8657;
wire n_11567;
wire n_6354;
wire n_10563;
wire n_5748;
wire n_17374;
wire n_321;
wire n_17152;
wire n_16250;
wire n_14050;
wire n_17094;
wire n_19732;
wire n_9569;
wire n_17836;
wire n_12463;
wire n_18232;
wire n_8071;
wire n_19432;
wire n_18822;
wire n_16355;
wire n_18169;
wire n_4615;
wire n_3044;
wire n_14088;
wire n_9227;
wire n_5657;
wire n_12510;
wire n_14364;
wire n_17750;
wire n_3579;
wire n_17663;
wire n_1667;
wire n_4067;
wire n_5114;
wire n_7587;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_10604;
wire n_18270;
wire n_18097;
wire n_2526;
wire n_19060;
wire n_1711;
wire n_10568;
wire n_20029;
wire n_18217;
wire n_451;
wire n_18132;
wire n_17680;
wire n_4464;
wire n_11317;
wire n_19850;
wire n_15854;
wire n_9147;
wire n_16394;
wire n_3180;
wire n_18319;
wire n_20377;
wire n_12132;
wire n_2119;
wire n_10803;
wire n_9658;
wire n_21080;
wire n_535;
wire n_17219;
wire n_17573;
wire n_3392;
wire n_11378;
wire n_10836;
wire n_5081;
wire n_2904;
wire n_12180;
wire n_20897;
wire n_12049;
wire n_14434;
wire n_19951;
wire n_9553;
wire n_4552;
wire n_12978;
wire n_19503;
wire n_19190;
wire n_10930;
wire n_9942;
wire n_13686;
wire n_837;
wire n_13842;
wire n_5406;
wire n_9213;
wire n_4328;
wire n_19707;
wire n_11391;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_18312;
wire n_20868;
wire n_18476;
wire n_4940;
wire n_15156;
wire n_9374;
wire n_19995;
wire n_14497;
wire n_1309;
wire n_8331;
wire n_8317;
wire n_20825;
wire n_14109;
wire n_5867;
wire n_17190;
wire n_17877;
wire n_3365;
wire n_12640;
wire n_7496;
wire n_3977;
wire n_10014;
wire n_10714;
wire n_14855;
wire n_4928;
wire n_18070;
wire n_12101;
wire n_16514;
wire n_11185;
wire n_7360;
wire n_6325;
wire n_12197;
wire n_2494;
wire n_1538;
wire n_17462;
wire n_8929;
wire n_14069;
wire n_4436;
wire n_5786;
wire n_15964;
wire n_18763;
wire n_9611;
wire n_1668;
wire n_9744;
wire n_16865;
wire n_1161;
wire n_8036;
wire n_4840;
wire n_20356;
wire n_4873;
wire n_9190;
wire n_15937;
wire n_1191;
wire n_7518;
wire n_10422;
wire n_7575;
wire n_8092;
wire n_16087;
wire n_10979;
wire n_6309;
wire n_9109;
wire n_10189;
wire n_20486;
wire n_18369;
wire n_408;
wire n_12702;
wire n_20078;
wire n_9741;
wire n_4766;
wire n_1632;
wire n_1929;
wire n_20097;
wire n_12211;
wire n_20270;
wire n_9021;
wire n_2929;
wire n_11145;
wire n_7579;
wire n_19153;
wire n_17795;
wire n_13982;
wire n_16979;
wire n_640;
wire n_6490;
wire n_10920;
wire n_11712;
wire n_19523;
wire n_13405;
wire n_16895;
wire n_16744;
wire n_1784;
wire n_17586;
wire n_3050;
wire n_13102;
wire n_8718;
wire n_18651;
wire n_16198;
wire n_19479;
wire n_15997;
wire n_15812;
wire n_3298;
wire n_5431;
wire n_12143;
wire n_5100;
wire n_1441;
wire n_1822;
wire n_9126;
wire n_2907;
wire n_2353;
wire n_10368;
wire n_686;
wire n_5746;
wire n_18781;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_20303;
wire n_19921;
wire n_1016;
wire n_8569;
wire n_10531;
wire n_4666;
wire n_18766;
wire n_12066;
wire n_8592;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_7952;
wire n_9998;
wire n_891;
wire n_13963;
wire n_885;
wire n_18298;
wire n_1864;
wire n_11121;
wire n_5414;
wire n_3086;
wire n_17667;
wire n_3165;
wire n_19771;
wire n_10035;
wire n_14523;
wire n_9045;
wire n_16233;
wire n_14883;
wire n_10107;
wire n_10283;
wire n_714;
wire n_17154;
wire n_8561;
wire n_6549;
wire n_9326;
wire n_18166;
wire n_5003;
wire n_20748;
wire n_6658;
wire n_6683;
wire n_154;
wire n_5745;
wire n_10050;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_15743;
wire n_5593;
wire n_6171;
wire n_5779;
wire n_20760;
wire n_7213;
wire n_20993;
wire n_5313;
wire n_2133;
wire n_14041;
wire n_12769;
wire n_8888;
wire n_1541;
wire n_9382;
wire n_11784;
wire n_20848;
wire n_7369;
wire n_15559;
wire n_14888;
wire n_9325;
wire n_9945;
wire n_9643;
wire n_13016;
wire n_7548;
wire n_12820;
wire n_18028;
wire n_7598;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_9771;
wire n_4715;
wire n_335;
wire n_19131;
wire n_344;
wire n_16031;
wire n_8794;
wire n_12689;
wire n_16827;
wire n_19025;
wire n_10095;
wire n_4078;
wire n_18612;
wire n_14812;
wire n_14000;
wire n_1624;
wire n_20250;
wire n_10488;
wire n_4418;
wire n_7924;
wire n_17946;
wire n_11103;
wire n_12420;
wire n_18363;
wire n_9232;
wire n_18187;
wire n_4125;
wire n_20408;
wire n_7012;
wire n_3043;
wire n_18160;
wire n_16599;
wire n_11837;
wire n_13501;
wire n_13533;
wire n_4527;
wire n_538;
wire n_2845;
wire n_9839;
wire n_7634;
wire n_1307;
wire n_7406;
wire n_19768;
wire n_19262;
wire n_2330;
wire n_13165;
wire n_5078;
wire n_7659;
wire n_3189;
wire n_16575;
wire n_4957;
wire n_15472;
wire n_9383;
wire n_1440;
wire n_11978;
wire n_11827;
wire n_19363;
wire n_7372;
wire n_6841;
wire n_11281;
wire n_16837;
wire n_361;
wire n_5624;
wire n_1065;
wire n_11772;
wire n_15837;
wire n_13448;
wire n_7371;
wire n_21017;
wire n_14752;
wire n_5447;
wire n_12153;
wire n_2692;
wire n_9621;
wire n_15966;
wire n_4102;
wire n_5755;
wire n_9158;
wire n_2553;
wire n_6889;
wire n_12586;
wire n_11993;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_11131;
wire n_12221;
wire n_17074;
wire n_8627;
wire n_1210;
wire n_14318;
wire n_18824;
wire n_19145;
wire n_8945;
wire n_9142;
wire n_9189;
wire n_18587;
wire n_1038;
wire n_4135;
wire n_6154;
wire n_19959;
wire n_14404;
wire n_12695;
wire n_11512;
wire n_20541;
wire n_14758;
wire n_20331;
wire n_20793;
wire n_10986;
wire n_15573;
wire n_10853;
wire n_13352;
wire n_20358;
wire n_11521;
wire n_10575;
wire n_8745;
wire n_5721;
wire n_7083;
wire n_18043;
wire n_316;
wire n_15889;
wire n_17473;
wire n_8260;
wire n_14153;
wire n_7143;
wire n_2303;
wire n_16939;
wire n_13484;
wire n_8688;
wire n_17661;
wire n_8279;
wire n_4639;
wire n_12864;
wire n_13478;
wire n_17989;
wire n_11042;
wire n_2154;
wire n_12570;
wire n_14124;
wire n_15932;
wire n_18407;
wire n_14344;
wire n_21015;
wire n_1986;
wire n_6818;
wire n_11761;
wire n_7209;
wire n_13374;
wire n_16906;
wire n_13182;
wire n_14867;
wire n_9871;
wire n_15632;
wire n_18923;
wire n_9698;
wire n_19566;
wire n_2881;
wire n_4270;
wire n_13690;
wire n_6255;
wire n_19891;
wire n_2305;
wire n_10026;
wire n_9731;
wire n_19589;
wire n_13577;
wire n_13098;
wire n_7237;
wire n_9642;
wire n_20808;
wire n_11189;
wire n_9050;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_12056;
wire n_15030;
wire n_8419;
wire n_10320;
wire n_975;
wire n_17875;
wire n_7304;
wire n_6266;
wire n_14905;
wire n_2503;
wire n_19988;
wire n_13362;
wire n_7754;
wire n_2989;
wire n_15631;
wire n_8826;
wire n_20493;
wire n_9732;
wire n_18742;
wire n_9685;
wire n_12529;
wire n_13983;
wire n_15856;
wire n_3389;
wire n_2126;
wire n_20233;
wire n_19942;
wire n_20627;
wire n_15058;
wire n_19869;
wire n_12473;
wire n_14295;
wire n_9378;
wire n_17112;
wire n_20678;
wire n_1445;
wire n_17268;
wire n_16859;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_14336;
wire n_11351;
wire n_8515;
wire n_18064;
wire n_11094;
wire n_332;
wire n_830;
wire n_5902;
wire n_3227;
wire n_11366;
wire n_8301;
wire n_18214;
wire n_9637;
wire n_5386;
wire n_4526;
wire n_4105;
wire n_10535;
wire n_969;
wire n_14655;
wire n_7180;
wire n_13778;
wire n_20420;
wire n_8972;
wire n_14709;
wire n_1630;
wire n_14606;
wire n_17672;
wire n_1720;
wire n_2409;
wire n_13913;
wire n_10313;
wire n_12983;
wire n_14003;
wire n_8891;
wire n_3897;
wire n_17733;
wire n_1735;
wire n_391;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_12313;
wire n_2597;
wire n_5980;
wire n_15114;
wire n_20244;
wire n_10445;
wire n_7771;
wire n_8810;
wire n_6469;
wire n_11119;
wire n_1271;
wire n_12696;
wire n_19559;
wire n_17644;
wire n_13730;
wire n_17627;
wire n_8932;
wire n_8264;
wire n_18034;
wire n_19256;
wire n_11954;
wire n_1323;
wire n_13438;
wire n_19731;
wire n_16813;
wire n_4142;
wire n_900;
wire n_5485;
wire n_10076;
wire n_5525;
wire n_17848;
wire n_14432;
wire n_1551;
wire n_13410;
wire n_9255;
wire n_12460;
wire n_8388;
wire n_15061;
wire n_5948;
wire n_8670;
wire n_20238;
wire n_7706;
wire n_15266;
wire n_13942;
wire n_2420;
wire n_7992;
wire n_7643;
wire n_9120;
wire n_19987;
wire n_16089;
wire n_20926;
wire n_15054;
wire n_9136;
wire n_1865;
wire n_18146;
wire n_7628;
wire n_19601;
wire n_15220;
wire n_16684;
wire n_483;
wire n_14013;
wire n_12065;
wire n_12275;
wire n_18745;
wire n_6035;
wire n_17301;
wire n_15669;
wire n_6405;
wire n_20557;
wire n_2235;
wire n_5850;
wire n_16751;
wire n_20747;
wire n_6786;
wire n_8299;
wire n_1848;
wire n_3776;
wire n_9060;
wire n_9792;
wire n_3778;
wire n_10801;
wire n_13013;
wire n_4322;
wire n_15744;
wire n_11217;
wire n_635;
wire n_12752;
wire n_19168;
wire n_1643;
wire n_4185;
wire n_3001;
wire n_19754;
wire n_18449;
wire n_2538;
wire n_14723;
wire n_19075;
wire n_4756;
wire n_11557;
wire n_18058;
wire n_2422;
wire n_19569;
wire n_654;
wire n_2933;
wire n_12715;
wire n_21077;
wire n_12787;
wire n_8636;
wire n_16345;
wire n_11442;
wire n_3584;
wire n_14102;
wire n_3446;
wire n_1059;
wire n_19481;
wire n_7592;
wire n_19824;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_17792;
wire n_2339;
wire n_392;
wire n_1866;
wire n_16243;
wire n_15052;
wire n_20429;
wire n_1558;
wire n_4107;
wire n_12722;
wire n_2519;
wire n_20819;
wire n_10821;
wire n_4361;
wire n_6219;
wire n_13590;
wire n_6445;
wire n_15778;
wire n_3137;
wire n_2544;
wire n_14887;
wire n_17394;
wire n_5612;
wire n_8493;
wire n_20187;
wire n_5172;
wire n_13670;
wire n_13148;
wire n_14962;
wire n_17992;
wire n_881;
wire n_1477;
wire n_6499;
wire n_1982;
wire n_20262;
wire n_5311;
wire n_19120;
wire n_290;
wire n_14506;
wire n_6842;
wire n_19834;
wire n_10079;
wire n_201;
wire n_2193;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_10361;
wire n_14154;
wire n_18644;
wire n_16454;
wire n_11635;
wire n_19181;
wire n_9571;
wire n_15703;
wire n_12323;
wire n_5379;
wire n_13387;
wire n_13068;
wire n_20601;
wire n_4329;
wire n_7696;
wire n_12015;
wire n_2562;
wire n_18103;
wire n_15992;
wire n_231;
wire n_11134;
wire n_8708;
wire n_10503;
wire n_5964;
wire n_6076;
wire n_10982;
wire n_12867;
wire n_13479;
wire n_13710;
wire n_1591;
wire n_14700;
wire n_15469;
wire n_8759;
wire n_18506;
wire n_6817;
wire n_5776;
wire n_2179;
wire n_14249;
wire n_9954;
wire n_18323;
wire n_7291;
wire n_13282;
wire n_17090;
wire n_3834;
wire n_8453;
wire n_18291;
wire n_583;
wire n_19892;
wire n_1000;
wire n_7017;
wire n_16649;
wire n_4072;
wire n_2792;
wire n_9640;
wire n_20402;
wire n_12411;
wire n_18052;
wire n_4026;
wire n_13295;
wire n_7889;
wire n_1702;
wire n_14349;
wire n_19152;
wire n_4852;
wire n_3202;
wire n_8968;
wire n_1082;
wire n_2318;
wire n_20430;
wire n_866;
wire n_21037;
wire n_2819;
wire n_11765;
wire n_18202;
wire n_7846;
wire n_3547;
wire n_2551;
wire n_3045;
wire n_9919;
wire n_20460;
wire n_15596;
wire n_11574;
wire n_2706;
wire n_13574;
wire n_17772;
wire n_14563;
wire n_12913;
wire n_1905;
wire n_13027;
wire n_1569;
wire n_5448;
wire n_17457;
wire n_19838;
wire n_15456;
wire n_6851;
wire n_4046;
wire n_17426;
wire n_7606;
wire n_9963;
wire n_18568;
wire n_3213;
wire n_1244;
wire n_14042;
wire n_19193;
wire n_13851;
wire n_19609;
wire n_4063;
wire n_19808;
wire n_13616;
wire n_12169;
wire n_893;
wire n_17175;
wire n_9426;
wire n_18767;
wire n_9293;
wire n_2824;
wire n_10065;
wire n_14500;
wire n_2089;
wire n_7896;
wire n_20564;
wire n_4688;
wire n_12657;
wire n_5900;
wire n_7319;
wire n_15721;
wire n_20697;
wire n_3619;
wire n_16977;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_2135;
wire n_4475;
wire n_6317;
wire n_17764;
wire n_10609;
wire n_13860;
wire n_6707;
wire n_13847;
wire n_18697;
wire n_12443;
wire n_17781;
wire n_4997;
wire n_19813;
wire n_7991;
wire n_781;
wire n_4090;
wire n_13610;
wire n_16021;
wire n_9302;
wire n_8258;
wire n_12781;
wire n_15991;
wire n_10506;
wire n_8416;
wire n_764;
wire n_12744;
wire n_1999;
wire n_11176;
wire n_4841;
wire n_11402;
wire n_17730;
wire n_8696;
wire n_9185;
wire n_18430;
wire n_2084;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_3905;
wire n_7163;
wire n_14845;
wire n_19367;
wire n_20675;
wire n_1836;
wire n_13164;
wire n_7027;
wire n_1453;
wire n_17679;
wire n_6964;
wire n_18193;
wire n_3145;
wire n_5749;
wire n_16716;
wire n_11711;
wire n_14541;
wire n_18774;
wire n_10941;
wire n_14689;
wire n_20740;
wire n_15667;
wire n_17701;
wire n_16797;
wire n_16190;
wire n_20823;
wire n_15588;
wire n_1746;
wire n_6610;
wire n_15919;
wire n_740;
wire n_16281;
wire n_13919;
wire n_6675;
wire n_9039;
wire n_12914;
wire n_12844;
wire n_7218;
wire n_5678;
wire n_16381;
wire n_7814;
wire n_8389;
wire n_2149;
wire n_12150;
wire n_16873;
wire n_18015;
wire n_16664;
wire n_13757;
wire n_15711;
wire n_19971;
wire n_21026;
wire n_7152;
wire n_2049;
wire n_7062;
wire n_2232;
wire n_5815;
wire n_15014;
wire n_1512;
wire n_5965;
wire n_16748;
wire n_4980;
wire n_18008;
wire n_17525;
wire n_20981;
wire n_2192;
wire n_19943;
wire n_7055;
wire n_693;
wire n_3207;
wire n_16160;
wire n_20461;
wire n_18988;
wire n_1637;
wire n_9864;
wire n_12144;
wire n_1751;
wire n_7056;
wire n_11486;
wire n_5310;
wire n_17640;
wire n_8680;
wire n_1548;
wire n_8394;
wire n_440;
wire n_14152;
wire n_20661;
wire n_7726;
wire n_2739;
wire n_11148;
wire n_6791;
wire n_13929;
wire n_6821;
wire n_2094;
wire n_13796;
wire n_3854;
wire n_13474;
wire n_10879;
wire n_12393;
wire n_2349;
wire n_17649;
wire n_18706;
wire n_19420;
wire n_3089;
wire n_9561;
wire n_20545;
wire n_17770;
wire n_16131;
wire n_19170;
wire n_942;
wire n_10705;
wire n_20721;
wire n_11032;
wire n_5234;
wire n_6890;
wire n_11454;
wire n_6988;
wire n_4747;
wire n_8000;
wire n_14686;
wire n_3472;
wire n_16542;
wire n_19643;
wire n_15179;
wire n_17062;
wire n_8709;
wire n_10504;
wire n_10687;
wire n_2806;
wire n_11045;
wire n_3191;
wire n_302;
wire n_2281;
wire n_8782;
wire n_10882;
wire n_5253;
wire n_10293;
wire n_355;
wire n_3280;
wire n_5418;
wire n_3095;
wire n_15584;
wire n_19219;
wire n_17495;
wire n_3698;
wire n_15493;
wire n_4513;
wire n_13152;
wire n_1442;
wire n_2620;
wire n_8716;
wire n_7264;
wire n_20168;
wire n_2549;
wire n_14829;
wire n_12631;
wire n_7492;
wire n_15331;
wire n_13546;
wire n_1656;
wire n_15791;
wire n_18050;
wire n_15687;
wire n_1562;
wire n_20341;
wire n_12455;
wire n_8266;
wire n_3407;
wire n_18354;
wire n_13601;
wire n_9214;
wire n_10090;
wire n_6512;
wire n_20613;
wire n_5342;
wire n_19764;
wire n_4843;
wire n_19355;
wire n_1418;
wire n_17926;
wire n_9991;
wire n_12880;
wire n_8457;
wire n_5795;
wire n_10763;
wire n_18322;
wire n_5715;
wire n_14997;
wire n_13918;
wire n_11180;
wire n_2155;
wire n_6231;
wire n_7503;
wire n_4795;
wire n_8124;
wire n_17976;
wire n_7997;
wire n_5659;
wire n_16510;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_18406;
wire n_13744;
wire n_18459;
wire n_3176;
wire n_20741;
wire n_3792;
wire n_8581;
wire n_10873;
wire n_19058;
wire n_5598;
wire n_17941;
wire n_2753;
wire n_13028;
wire n_19617;
wire n_3805;
wire n_3950;
wire n_9650;
wire n_11497;
wire n_20873;
wire n_17930;
wire n_6912;
wire n_3567;
wire n_5112;
wire n_5326;
wire n_14078;
wire n_20775;
wire n_5303;
wire n_3127;
wire n_6916;
wire n_9282;
wire n_18408;
wire n_8289;
wire n_19225;
wire n_10447;
wire n_20374;
wire n_13549;
wire n_11029;
wire n_6492;
wire n_17867;
wire n_1913;
wire n_13036;
wire n_15603;
wire n_9237;
wire n_18087;
wire n_6857;
wire n_20824;
wire n_16309;
wire n_10292;
wire n_20744;
wire n_7763;
wire n_13258;
wire n_16681;
wire n_16423;
wire n_20764;
wire n_13827;
wire n_12576;
wire n_14350;
wire n_3467;
wire n_5262;
wire n_18711;
wire n_16887;
wire n_18011;
wire n_20164;
wire n_20419;
wire n_927;
wire n_7469;
wire n_10163;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7856;
wire n_18314;
wire n_3816;
wire n_8099;
wire n_10876;
wire n_15092;
wire n_15397;
wire n_11449;
wire n_4725;
wire n_348;
wire n_10352;
wire n_9173;
wire n_2312;
wire n_13714;
wire n_1826;
wire n_14565;
wire n_20876;
wire n_2834;
wire n_18282;
wire n_4563;
wire n_637;
wire n_7128;
wire n_9849;
wire n_15454;
wire n_5335;
wire n_11096;
wire n_8459;
wire n_2801;
wire n_12288;
wire n_4334;
wire n_13025;
wire n_17449;
wire n_2718;
wire n_18389;
wire n_6950;
wire n_4923;
wire n_8540;
wire n_7057;
wire n_17695;
wire n_1802;
wire n_9823;
wire n_20918;
wire n_5168;
wire n_3200;
wire n_4274;
wire n_5583;
wire n_12629;
wire n_5433;
wire n_12893;
wire n_9281;
wire n_9103;
wire n_7088;
wire n_10883;
wire n_4007;
wire n_8433;
wire n_17957;
wire n_10429;
wire n_12732;
wire n_7048;
wire n_12569;
wire n_16673;
wire n_20684;
wire n_16629;
wire n_16885;
wire n_10859;
wire n_17745;
wire n_16756;
wire n_20098;
wire n_17059;
wire n_1134;
wire n_12980;
wire n_647;
wire n_18557;
wire n_2932;
wire n_8409;
wire n_16093;
wire n_11616;
wire n_14831;
wire n_9170;
wire n_17521;
wire n_3039;
wire n_5455;
wire n_2195;
wire n_6777;
wire n_16303;
wire n_6742;
wire n_16444;
wire n_20648;
wire n_6307;
wire n_14129;
wire n_16049;
wire n_4523;
wire n_13280;
wire n_8415;
wire n_3022;
wire n_6479;
wire n_11472;
wire n_13073;
wire n_3286;
wire n_5619;
wire n_2023;
wire n_13083;
wire n_5022;
wire n_9223;
wire n_19258;
wire n_2031;
wire n_5353;
wire n_9781;
wire n_3009;
wire n_7095;
wire n_6140;
wire n_18263;
wire n_20682;
wire n_20509;
wire n_18129;
wire n_16930;
wire n_9970;
wire n_5518;
wire n_14882;
wire n_17823;
wire n_15488;
wire n_7037;
wire n_17133;
wire n_18576;
wire n_1823;
wire n_20768;
wire n_5236;
wire n_10077;
wire n_3942;
wire n_3023;
wire n_17754;
wire n_10964;
wire n_14367;
wire n_9492;
wire n_10759;
wire n_9226;
wire n_19460;
wire n_1607;
wire n_221;
wire n_20842;
wire n_14363;
wire n_17932;
wire n_19518;
wire n_5814;
wire n_13526;
wire n_2256;
wire n_11488;
wire n_20438;
wire n_19106;
wire n_6069;
wire n_6515;
wire n_20001;
wire n_9513;
wire n_18180;
wire n_13267;
wire n_15249;
wire n_5671;
wire n_527;
wire n_20951;
wire n_10886;
wire n_20195;
wire n_10804;
wire n_7581;
wire n_343;
wire n_17968;
wire n_16875;
wire n_13834;
wire n_8935;
wire n_15081;
wire n_19372;
wire n_20112;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_19509;
wire n_13067;
wire n_2449;
wire n_16565;
wire n_12808;
wire n_20512;
wire n_12853;
wire n_8397;
wire n_17984;
wire n_18770;
wire n_17565;
wire n_6576;
wire n_9083;
wire n_17886;
wire n_1266;
wire n_14727;
wire n_13717;
wire n_6708;
wire n_10252;
wire n_16229;
wire n_9175;
wire n_15280;
wire n_6847;
wire n_8974;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_19659;
wire n_16952;
wire n_12965;
wire n_657;
wire n_14184;
wire n_15207;
wire n_7595;
wire n_2306;
wire n_7426;
wire n_2414;
wire n_17066;
wire n_5434;
wire n_6855;
wire n_14257;
wire n_8170;
wire n_1030;
wire n_13673;
wire n_20073;
wire n_19070;
wire n_2737;
wire n_12263;
wire n_9830;
wire n_14416;
wire n_9116;
wire n_8825;
wire n_4351;
wire n_8003;
wire n_1301;
wire n_8395;
wire n_13986;
wire n_18826;
wire n_14963;
wire n_20999;
wire n_5146;
wire n_7367;
wire n_11537;
wire n_8164;
wire n_11583;
wire n_4221;
wire n_8877;
wire n_16477;
wire n_1993;
wire n_134;
wire n_16385;
wire n_2540;
wire n_8476;
wire n_6218;
wire n_7685;
wire n_4009;
wire n_15237;
wire n_18848;
wire n_12299;
wire n_11929;
wire n_11340;
wire n_17091;
wire n_5577;
wire n_876;
wire n_9100;
wire n_15007;
wire n_15337;
wire n_13523;
wire n_17537;
wire n_10677;
wire n_18795;
wire n_2627;
wire n_1327;
wire n_10648;
wire n_19841;
wire n_5976;
wire n_9249;
wire n_4739;
wire n_19047;
wire n_17422;
wire n_8256;
wire n_4312;
wire n_14751;
wire n_10273;
wire n_12927;
wire n_1658;
wire n_1072;
wire n_18575;
wire n_1305;
wire n_1873;
wire n_13430;
wire n_10097;
wire n_2725;
wire n_19014;
wire n_19558;
wire n_13732;
wire n_20696;
wire n_18843;
wire n_12887;
wire n_15496;
wire n_16256;
wire n_5456;
wire n_4847;
wire n_3702;
wire n_10462;
wire n_20376;
wire n_1984;
wire n_12414;
wire n_12600;
wire n_7040;
wire n_2815;
wire n_4427;
wire n_7740;
wire n_4705;
wire n_15149;
wire n_6794;
wire n_819;
wire n_2945;
wire n_11205;
wire n_586;
wire n_10832;
wire n_9327;
wire n_2936;
wire n_18467;
wire n_16219;
wire n_10142;
wire n_10300;
wire n_18283;
wire n_1642;
wire n_14220;
wire n_12783;
wire n_20985;
wire n_12431;
wire n_8971;
wire n_3907;
wire n_4603;
wire n_4332;
wire n_17362;
wire n_9291;
wire n_19428;
wire n_20837;
wire n_3388;
wire n_15385;
wire n_8215;
wire n_5201;
wire n_20089;
wire n_5551;
wire n_16762;
wire n_2377;
wire n_14644;
wire n_17450;
wire n_5498;
wire n_16172;
wire n_7765;
wire n_14022;
wire n_20717;
wire n_12974;
wire n_1685;
wire n_2222;
wire n_17010;
wire n_13849;
wire n_12121;
wire n_12658;
wire n_13956;
wire n_19592;
wire n_10607;
wire n_2076;
wire n_19351;
wire n_19963;
wire n_19350;
wire n_14314;
wire n_15088;
wire n_5252;
wire n_11259;
wire n_5777;
wire n_19527;
wire n_8942;
wire n_7785;
wire n_18755;
wire n_5063;
wire n_14628;
wire n_18458;
wire n_4712;
wire n_7181;
wire n_11443;
wire n_19098;
wire n_858;
wire n_7355;
wire n_15449;
wire n_11161;
wire n_11770;
wire n_2136;
wire n_13509;
wire n_433;
wire n_7328;
wire n_17933;
wire n_18168;
wire n_2403;
wire n_5643;
wire n_9826;
wire n_11810;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_7916;
wire n_18853;
wire n_3055;
wire n_15862;
wire n_420;
wire n_5346;
wire n_7283;
wire n_18336;
wire n_20178;
wire n_1045;
wire n_14954;
wire n_14890;
wire n_16808;
wire n_10518;
wire n_11789;
wire n_1881;
wire n_2635;
wire n_20248;
wire n_20640;
wire n_4139;
wire n_6130;
wire n_16613;
wire n_6417;
wire n_368;
wire n_4867;
wire n_19873;
wire n_2713;
wire n_18786;
wire n_1965;
wire n_19826;
wire n_4450;
wire n_13725;
wire n_6979;
wire n_16876;
wire n_10971;
wire n_15757;
wire n_12341;
wire n_13297;
wire n_19540;
wire n_11854;
wire n_2210;
wire n_19928;
wire n_3141;
wire n_2053;
wire n_19354;
wire n_18250;
wire n_16593;
wire n_16097;
wire n_20428;
wire n_2450;
wire n_6831;
wire n_14302;
wire n_312;
wire n_20117;
wire n_728;
wire n_10340;
wire n_20488;
wire n_5722;
wire n_16043;
wire n_14170;
wire n_10681;
wire n_14303;
wire n_15077;
wire n_18318;
wire n_2478;
wire n_15202;
wire n_3509;
wire n_453;
wire n_6458;
wire n_12768;
wire n_19636;
wire n_6986;
wire n_15409;
wire n_601;
wire n_8313;
wire n_11382;
wire n_14298;
wire n_7775;
wire n_907;
wire n_5734;
wire n_15831;
wire n_20021;
wire n_747;
wire n_12543;
wire n_1135;
wire n_11254;
wire n_14797;
wire n_19370;
wire n_19857;
wire n_5774;
wire n_11388;
wire n_6546;
wire n_15548;
wire n_11043;
wire n_7186;
wire n_593;
wire n_1695;
wire n_4650;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_18120;
wire n_9340;
wire n_12774;
wire n_20687;
wire n_15892;
wire n_12653;
wire n_11824;
wire n_3478;
wire n_10226;
wire n_14515;
wire n_16052;
wire n_19582;
wire n_19721;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_12052;
wire n_3836;
wire n_19608;
wire n_9064;
wire n_14968;
wire n_14721;
wire n_11533;
wire n_4469;
wire n_16017;
wire n_19877;
wire n_8497;
wire n_18242;
wire n_5959;
wire n_16597;
wire n_8210;
wire n_8056;
wire n_3310;
wire n_7748;
wire n_13298;
wire n_540;
wire n_5668;
wire n_4703;
wire n_7686;
wire n_20632;
wire n_14391;
wire n_9817;
wire n_12505;
wire n_15546;
wire n_1587;
wire n_12875;
wire n_19127;
wire n_13794;
wire n_4804;
wire n_17414;
wire n_1014;
wire n_15126;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_13542;
wire n_10470;
wire n_12828;
wire n_18546;
wire n_9059;
wire n_11691;
wire n_9812;
wire n_2927;
wire n_3833;
wire n_9912;
wire n_11513;
wire n_9620;
wire n_15051;
wire n_7930;
wire n_13241;
wire n_580;
wire n_7077;
wire n_15037;
wire n_1183;
wire n_17359;
wire n_11111;
wire n_13270;
wire n_2889;
wire n_11938;
wire n_6043;
wire n_9497;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_14543;
wire n_7024;
wire n_17372;
wire n_15523;
wire n_12659;
wire n_13934;
wire n_5925;
wire n_5591;
wire n_18504;
wire n_18046;
wire n_20694;
wire n_15970;
wire n_19254;
wire n_15260;
wire n_3292;
wire n_16340;
wire n_13591;
wire n_8377;
wire n_10558;
wire n_16518;
wire n_20899;
wire n_1057;
wire n_18040;
wire n_978;
wire n_1509;
wire n_10044;
wire n_14919;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_13354;
wire n_8957;
wire n_5047;
wire n_20998;
wire n_6938;
wire n_2197;
wire n_12709;
wire n_4778;
wire n_18891;
wire n_556;
wire n_16428;
wire n_4667;
wire n_17838;
wire n_16772;
wire n_20643;
wire n_9381;
wire n_17928;
wire n_8904;
wire n_16725;
wire n_14683;
wire n_20535;
wire n_13887;
wire n_12968;
wire n_15107;
wire n_17686;
wire n_1620;
wire n_18377;
wire n_18648;
wire n_18589;
wire n_7110;
wire n_12111;
wire n_17079;
wire n_18818;
wire n_19627;
wire n_20214;
wire n_8527;
wire n_20672;
wire n_13419;
wire n_13383;
wire n_4578;
wire n_11424;
wire n_3644;
wire n_12178;
wire n_20496;
wire n_2176;
wire n_17951;
wire n_6138;
wire n_528;
wire n_16333;
wire n_9296;
wire n_10662;
wire n_2065;
wire n_19482;
wire n_7038;
wire n_4187;
wire n_13420;
wire n_16714;
wire n_8341;
wire n_16006;
wire n_10200;
wire n_18284;
wire n_14436;
wire n_5576;
wire n_8308;
wire n_18906;
wire n_17367;
wire n_14651;
wire n_10632;
wire n_16083;
wire n_9365;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_11166;
wire n_14881;
wire n_2967;
wire n_9869;
wire n_20273;
wire n_7757;
wire n_6242;
wire n_14143;
wire n_336;
wire n_6601;
wire n_12536;
wire n_2268;
wire n_10041;
wire n_12168;
wire n_19725;
wire n_19910;
wire n_12533;
wire n_20633;
wire n_20606;
wire n_18844;
wire n_2111;
wire n_18502;
wire n_17999;
wire n_9615;
wire n_11869;
wire n_5015;
wire n_5527;
wire n_9759;
wire n_9711;
wire n_13171;
wire n_4497;
wire n_6606;
wire n_8291;
wire n_9820;
wire n_7758;
wire n_19234;
wire n_11060;
wire n_9321;
wire n_11493;
wire n_19685;
wire n_1640;
wire n_8375;
wire n_13462;
wire n_10280;
wire n_9428;
wire n_11452;
wire n_15366;
wire n_7705;
wire n_18410;
wire n_2505;
wire n_17717;
wire n_369;
wire n_7333;
wire n_12246;
wire n_12297;
wire n_8006;
wire n_9565;
wire n_8491;
wire n_13089;
wire n_7337;
wire n_5726;
wire n_16336;
wire n_10483;
wire n_11864;
wire n_694;
wire n_6228;
wire n_16030;
wire n_15990;
wire n_4749;
wire n_14536;
wire n_5545;
wire n_16174;
wire n_8458;
wire n_1470;
wire n_3253;
wire n_16819;
wire n_17176;
wire n_19498;
wire n_6997;
wire n_6371;
wire n_904;
wire n_19595;
wire n_2005;
wire n_19253;
wire n_1696;
wire n_14642;
wire n_14809;
wire n_8013;
wire n_2108;
wire n_2246;
wire n_18713;
wire n_10250;
wire n_3846;
wire n_12682;
wire n_10831;
wire n_17180;
wire n_18221;
wire n_12621;
wire n_20255;
wire n_10172;
wire n_10333;
wire n_4668;
wire n_9868;
wire n_5782;
wire n_8119;
wire n_16460;
wire n_630;
wire n_1369;
wire n_20546;
wire n_7370;
wire n_7931;
wire n_12225;
wire n_15245;
wire n_18544;
wire n_19711;
wire n_16784;
wire n_19876;
wire n_15858;
wire n_12126;
wire n_15003;
wire n_10588;
wire n_5637;
wire n_7480;
wire n_12158;
wire n_8843;
wire n_13232;
wire n_16414;
wire n_13859;
wire n_5034;
wire n_8694;
wire n_10643;
wire n_8752;
wire n_3672;
wire n_14058;
wire n_2839;
wire n_16622;
wire n_10905;
wire n_11859;
wire n_17900;
wire n_15025;
wire n_5269;
wire n_16949;
wire n_1764;
wire n_19645;
wire n_11023;
wire n_8770;
wire n_18990;
wire n_5115;
wire n_7376;
wire n_16992;
wire n_902;
wire n_17016;
wire n_4915;
wire n_1946;
wire n_18868;
wire n_4383;
wire n_17093;
wire n_596;
wire n_8391;
wire n_20159;
wire n_4485;
wire n_6388;
wire n_5163;
wire n_16852;
wire n_4356;
wire n_9628;
wire n_10854;
wire n_14309;
wire n_13652;
wire n_1516;
wire n_13207;
wire n_4890;
wire n_15963;
wire n_11528;
wire n_8631;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_9730;
wire n_16556;
wire n_18245;
wire n_2209;
wire n_14423;
wire n_13128;
wire n_12177;
wire n_7586;
wire n_4244;
wire n_12141;
wire n_19994;
wire n_6738;
wire n_2081;
wire n_1474;
wire n_12795;
wire n_1794;
wire n_13370;
wire n_1375;
wire n_5014;
wire n_6346;
wire n_3772;
wire n_7026;
wire n_15286;
wire n_10560;
wire n_13103;
wire n_263;
wire n_360;
wire n_13720;
wire n_18142;
wire n_2798;
wire n_10773;
wire n_17458;
wire n_165;
wire n_15962;
wire n_16098;
wire n_20265;
wire n_1249;
wire n_16148;
wire n_5724;
wire n_340;
wire n_3201;
wire n_12622;
wire n_10391;
wire n_12857;
wire n_10630;
wire n_4467;
wire n_15785;
wire n_20399;
wire n_177;
wire n_18845;
wire n_17954;
wire n_10540;
wire n_17135;
wire n_21097;
wire n_15140;
wire n_3935;
wire n_1861;
wire n_12287;
wire n_12182;
wire n_8924;
wire n_4955;
wire n_16968;
wire n_18249;
wire n_447;
wire n_14258;
wire n_17742;
wire n_7025;
wire n_20869;
wire n_3798;
wire n_5241;
wire n_12492;
wire n_4248;
wire n_2228;
wire n_13231;
wire n_7478;
wire n_841;
wire n_3204;
wire n_7451;
wire n_15918;
wire n_20767;
wire n_5258;
wire n_18426;
wire n_16050;
wire n_14741;
wire n_18741;
wire n_19430;
wire n_6790;
wire n_8165;
wire n_12760;
wire n_11172;
wire n_17446;
wire n_17159;
wire n_15154;
wire n_6002;
wire n_11458;
wire n_18624;
wire n_1250;
wire n_5717;
wire n_10794;
wire n_18378;
wire n_13125;
wire n_16166;
wire n_2002;
wire n_14658;
wire n_12589;
wire n_5791;
wire n_20732;
wire n_20686;
wire n_21056;
wire n_10000;
wire n_11783;
wire n_17615;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_11799;
wire n_17873;
wire n_8699;
wire n_1131;
wire n_2653;
wire n_16300;
wire n_11377;
wire n_11246;
wire n_19284;
wire n_3115;
wire n_14066;
wire n_9985;
wire n_20048;
wire n_10169;
wire n_16759;
wire n_13755;
wire n_19267;
wire n_18633;
wire n_19038;
wire n_1985;
wire n_14226;
wire n_16188;
wire n_4853;
wire n_5229;
wire n_15921;
wire n_8449;
wire n_10968;
wire n_3348;
wire n_12315;
wire n_10688;
wire n_3261;
wire n_16157;
wire n_9466;
wire n_8953;
wire n_7368;
wire n_9787;
wire n_8598;
wire n_15671;
wire n_7562;
wire n_20346;
wire n_18163;
wire n_4512;
wire n_4132;
wire n_17430;
wire n_4500;
wire n_18915;
wire n_9318;
wire n_13715;
wire n_19203;
wire n_12671;
wire n_8720;
wire n_2663;
wire n_6539;
wire n_20746;
wire n_8422;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_16841;
wire n_17501;
wire n_7392;
wire n_9714;
wire n_16147;
wire n_1428;
wire n_1284;
wire n_10131;
wire n_11721;
wire n_14430;
wire n_4143;
wire n_19244;
wire n_11891;
wire n_14094;
wire n_11492;
wire n_2359;
wire n_9354;
wire n_12647;
wire n_6249;
wire n_18512;
wire n_9058;
wire n_6197;
wire n_19361;
wire n_3254;
wire n_2227;
wire n_15161;
wire n_5589;
wire n_18937;
wire n_16768;
wire n_12080;
wire n_1676;
wire n_6295;
wire n_11409;
wire n_823;
wire n_13138;
wire n_10644;
wire n_16369;
wire n_352;
wire n_19308;
wire n_18170;
wire n_9516;
wire n_365;
wire n_13996;
wire n_15788;
wire n_5158;
wire n_12185;
wire n_20280;
wire n_8939;
wire n_11652;
wire n_1917;
wire n_5092;
wire n_6542;
wire n_18338;
wire n_15930;
wire n_3612;
wire n_4505;
wire n_20482;
wire n_1840;
wire n_8715;
wire n_6740;
wire n_13458;
wire n_17244;
wire n_19991;
wire n_2956;
wire n_5292;
wire n_8991;
wire n_7438;
wire n_8855;
wire n_19525;
wire n_13762;
wire n_17482;
wire n_20765;
wire n_5086;
wire n_1949;
wire n_18927;
wire n_14236;
wire n_11309;
wire n_14156;
wire n_13118;
wire n_8630;
wire n_9308;
wire n_11233;
wire n_7108;
wire n_11047;
wire n_9638;
wire n_1121;
wire n_15057;
wire n_15429;
wire n_8435;
wire n_5060;
wire n_18643;
wire n_13290;
wire n_15828;
wire n_13379;
wire n_2263;
wire n_3518;
wire n_2116;
wire n_13838;
wire n_10715;
wire n_19471;
wire n_11381;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_11922;
wire n_249;
wire n_444;
wire n_18954;
wire n_7850;
wire n_5076;
wire n_6872;
wire n_15357;
wire n_17042;
wire n_18675;
wire n_16387;
wire n_4912;
wire n_14505;
wire n_8542;
wire n_14292;
wire n_19123;
wire n_8373;
wire n_9304;
wire n_6236;
wire n_11152;
wire n_13505;
wire n_17328;
wire n_366;
wire n_2791;
wire n_14951;
wire n_4871;
wire n_12517;
wire n_20072;
wire n_16228;
wire n_6563;
wire n_5968;
wire n_992;
wire n_966;
wire n_13821;
wire n_14065;
wire n_8519;
wire n_14958;
wire n_8075;
wire n_5468;
wire n_7638;
wire n_19778;
wire n_4233;
wire n_4791;
wire n_8642;
wire n_11713;
wire n_8648;
wire n_16666;
wire n_7224;
wire n_9934;
wire n_14639;
wire n_1178;
wire n_2015;
wire n_13186;
wire n_15101;
wire n_13463;
wire n_5984;
wire n_14039;
wire n_6705;
wire n_20050;
wire n_203;
wire n_8585;
wire n_3000;
wire n_2930;
wire n_17934;
wire n_16404;
wire n_19278;
wire n_9717;
wire n_16418;
wire n_16283;
wire n_18450;
wire n_14788;
wire n_10638;
wire n_14559;
wire n_2161;
wire n_13353;
wire n_6624;
wire n_7888;
wire n_17323;
wire n_11525;
wire n_6883;
wire n_9558;
wire n_16633;
wire n_15615;
wire n_17308;
wire n_428;
wire n_18148;
wire n_12967;
wire n_2257;
wire n_1343;
wire n_12907;
wire n_3116;
wire n_17664;
wire n_15368;
wire n_3784;
wire n_4422;
wire n_11087;
wire n_8814;
wire n_10394;
wire n_14368;
wire n_1780;
wire n_2825;
wire n_20466;
wire n_13394;
wire n_5974;
wire n_10917;
wire n_5723;
wire n_15815;
wire n_18613;
wire n_5922;
wire n_6378;
wire n_17970;
wire n_21070;
wire n_17556;
wire n_20921;
wire n_11483;
wire n_7488;
wire n_4307;
wire n_16567;
wire n_18200;
wire n_382;
wire n_20093;
wire n_4438;
wire n_19437;
wire n_11568;
wire n_3814;
wire n_11468;
wire n_7599;
wire n_7231;
wire n_6579;
wire n_12711;
wire n_16651;
wire n_1447;
wire n_19916;
wire n_12216;
wire n_9003;
wire n_18126;
wire n_12879;
wire n_20205;
wire n_16879;
wire n_17193;
wire n_20854;
wire n_5454;
wire n_19552;
wire n_17716;
wire n_4254;
wire n_11206;
wire n_18340;
wire n_12649;
wire n_8913;
wire n_404;
wire n_8355;
wire n_12447;
wire n_17224;
wire n_15910;
wire n_13822;
wire n_299;
wire n_7168;
wire n_15514;
wire n_11927;
wire n_11676;
wire n_19160;
wire n_2649;
wire n_6461;
wire n_2919;
wire n_3108;
wire n_15719;
wire n_18117;
wire n_5557;
wire n_20418;
wire n_6914;
wire n_8816;
wire n_15873;
wire n_8418;
wire n_14943;
wire n_16145;
wire n_15684;
wire n_3239;
wire n_19541;
wire n_10668;
wire n_8739;
wire n_12053;
wire n_13250;
wire n_1817;
wire n_13228;
wire n_7963;
wire n_17528;
wire n_15278;
wire n_20252;
wire n_21086;
wire n_14326;
wire n_15335;
wire n_4296;
wire n_138;
wire n_162;
wire n_13100;
wire n_16926;
wire n_2483;
wire n_18559;
wire n_7938;
wire n_20038;
wire n_18991;
wire n_17939;
wire n_2655;
wire n_9270;
wire n_11373;
wire n_17212;
wire n_20594;
wire n_19345;
wire n_13185;
wire n_9483;
wire n_720;
wire n_6263;
wire n_14593;
wire n_6731;
wire n_8156;
wire n_8845;
wire n_10229;
wire n_12268;
wire n_9256;
wire n_3054;
wire n_21043;
wire n_1868;
wire n_3601;
wire n_11107;
wire n_3881;
wire n_13195;
wire n_12298;
wire n_6224;
wire n_8510;
wire n_9854;
wire n_2099;
wire n_9737;
wire n_19324;
wire n_11154;
wire n_20563;
wire n_18233;
wire n_19295;
wire n_19635;
wire n_18195;
wire n_10358;
wire n_20075;
wire n_20076;
wire n_808;
wire n_4133;
wire n_2636;
wire n_17464;
wire n_6903;
wire n_15466;
wire n_2074;
wire n_6768;
wire n_19825;
wire n_12382;
wire n_9679;
wire n_15413;
wire n_17353;
wire n_17732;
wire n_8978;
wire n_14279;
wire n_6189;
wire n_15339;
wire n_9699;
wire n_16686;
wire n_20379;
wire n_9673;
wire n_15313;
wire n_19027;
wire n_11823;
wire n_18696;
wire n_17855;
wire n_1304;
wire n_14033;
wire n_3335;
wire n_5960;
wire n_16778;
wire n_478;
wire n_18931;
wire n_1349;
wire n_10261;
wire n_14045;
wire n_2102;
wire n_18238;
wire n_11806;
wire n_3477;
wire n_7868;
wire n_16999;
wire n_16238;
wire n_2286;
wire n_18971;
wire n_15034;
wire n_3036;
wire n_14305;
wire n_12421;
wire n_10730;
wire n_19977;
wire n_1162;
wire n_9146;
wire n_14835;
wire n_7176;
wire n_8565;
wire n_12133;
wire n_15167;
wire n_442;
wire n_11970;
wire n_3764;
wire n_13283;
wire n_4773;
wire n_5028;
wire n_9573;
wire n_986;
wire n_1104;
wire n_19211;
wire n_13327;
wire n_18712;
wire n_16921;
wire n_20042;
wire n_13534;
wire n_15356;
wire n_5123;
wire n_6689;
wire n_14846;
wire n_13992;
wire n_19118;
wire n_17178;
wire n_8753;
wire n_15230;
wire n_4856;
wire n_2707;
wire n_18809;
wire n_8325;
wire n_19539;
wire n_10875;
wire n_17590;
wire n_15018;
wire n_14071;
wire n_16825;
wire n_15256;
wire n_13097;
wire n_11261;
wire n_18964;
wire n_12579;
wire n_4229;
wire n_10564;
wire n_3337;
wire n_3750;
wire n_12342;
wire n_12877;
wire n_1523;
wire n_2516;
wire n_11893;
wire n_20472;
wire n_19375;
wire n_8677;
wire n_5818;
wire n_15525;
wire n_7869;
wire n_12468;
wire n_3710;
wire n_12426;
wire n_6943;
wire n_1957;
wire n_19270;
wire n_14555;
wire n_5889;
wire n_8602;
wire n_9609;
wire n_10284;
wire n_3944;
wire n_21101;
wire n_18761;
wire n_16343;
wire n_5632;
wire n_17060;
wire n_13569;
wire n_5613;
wire n_7472;
wire n_1373;
wire n_17270;
wire n_17551;
wire n_5450;
wire n_18646;
wire n_18870;
wire n_15622;
wire n_18928;
wire n_4781;
wire n_14328;
wire n_15457;
wire n_11722;
wire n_3333;
wire n_12149;
wire n_20885;
wire n_9557;
wire n_16991;
wire n_8039;
wire n_8193;
wire n_12116;
wire n_9073;
wire n_8432;
wire n_16088;
wire n_5374;
wire n_2424;
wire n_6456;
wire n_722;
wire n_17234;
wire n_13158;
wire n_12014;
wire n_9388;
wire n_14061;
wire n_11610;
wire n_16307;
wire n_2978;
wire n_6328;
wire n_11498;
wire n_11509;
wire n_15097;
wire n_14401;
wire n_14034;
wire n_15518;
wire n_15820;
wire n_2958;
wire n_1714;
wire n_11706;
wire n_7182;
wire n_11055;
wire n_8591;
wire n_5511;
wire n_13512;
wire n_8661;
wire n_10068;
wire n_9672;
wire n_9187;
wire n_9572;
wire n_12615;
wire n_20161;
wire n_16771;
wire n_19007;
wire n_7375;
wire n_8189;
wire n_13858;
wire n_266;
wire n_7736;
wire n_6435;
wire n_13949;
wire n_20110;
wire n_3646;
wire n_7419;
wire n_19941;
wire n_6600;
wire n_14087;
wire n_13681;
wire n_13700;
wire n_16095;
wire n_10277;
wire n_15242;
wire n_19081;
wire n_3864;
wire n_9251;
wire n_6201;
wire n_20053;
wire n_20103;
wire n_19415;
wire n_7918;
wire n_10331;
wire n_1406;
wire n_9181;
wire n_6803;
wire n_4288;
wire n_20864;
wire n_10981;
wire n_14063;
wire n_4511;
wire n_3422;
wire n_17594;
wire n_14521;
wire n_4675;
wire n_13701;
wire n_695;
wire n_17839;
wire n_11934;
wire n_13518;
wire n_2991;
wire n_16506;
wire n_14737;
wire n_386;
wire n_11969;
wire n_4289;
wire n_19648;
wire n_197;
wire n_8775;
wire n_678;
wire n_10158;
wire n_5077;
wire n_16173;
wire n_20193;
wire n_15852;
wire n_8804;
wire n_9577;
wire n_6573;
wire n_13805;
wire n_7385;
wire n_15425;
wire n_9802;
wire n_19467;
wire n_4846;
wire n_12381;
wire n_283;
wire n_9171;
wire n_18397;
wire n_13443;
wire n_374;
wire n_17046;
wire n_19914;
wire n_20491;
wire n_6756;
wire n_2606;
wire n_15268;
wire n_5826;
wire n_8697;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_14712;
wire n_9408;
wire n_7847;
wire n_18560;
wire n_16189;
wire n_2417;
wire n_6059;
wire n_14976;
wire n_17428;
wire n_8063;
wire n_3313;
wire n_13798;
wire n_15580;
wire n_2354;
wire n_14474;
wire n_3945;
wire n_14112;
wire n_18009;
wire n_10477;
wire n_11904;
wire n_10296;
wire n_19456;
wire n_17574;
wire n_13676;
wire n_1256;
wire n_5365;
wire n_9566;
wire n_15528;
wire n_6188;
wire n_10066;
wire n_11755;
wire n_19488;
wire n_16616;
wire n_4630;
wire n_18374;
wire n_20028;
wire n_16916;
wire n_4829;
wire n_12956;
wire n_7831;
wire n_18966;
wire n_5259;
wire n_15365;
wire n_18693;
wire n_18584;
wire n_11129;
wire n_20762;
wire n_4966;
wire n_18985;
wire n_6104;
wire n_15476;
wire n_20129;
wire n_15444;
wire n_1303;
wire n_2506;
wire n_9822;
wire n_1593;
wire n_2610;
wire n_10036;
wire n_15199;
wire n_19536;
wire n_2626;
wire n_10749;
wire n_7315;
wire n_21002;
wire n_16312;
wire n_5006;
wire n_14200;
wire n_3206;
wire n_4878;
wire n_6706;
wire n_4202;
wire n_6909;
wire n_13933;
wire n_6487;
wire n_12668;
wire n_10348;
wire n_13884;
wire n_1192;
wire n_20973;
wire n_3098;
wire n_4503;
wire n_15975;
wire n_17847;
wire n_12928;
wire n_5205;
wire n_16202;
wire n_19800;
wire n_13112;
wire n_17682;
wire n_7452;
wire n_15767;
wire n_7972;
wire n_13455;
wire n_8672;
wire n_20567;
wire n_3921;
wire n_282;
wire n_14280;
wire n_13946;
wire n_2766;
wire n_11270;
wire n_14961;
wire n_10722;
wire n_8847;
wire n_5508;
wire n_16659;
wire n_11344;
wire n_3851;
wire n_16624;
wire n_6500;
wire n_12847;
wire n_1048;
wire n_667;
wire n_7573;
wire n_2411;
wire n_8191;
wire n_13758;
wire n_18211;
wire n_11511;
wire n_20749;
wire n_6421;
wire n_10322;
wire n_5377;
wire n_6180;
wire n_20778;
wire n_20066;
wire n_7890;
wire n_17729;
wire n_19028;
wire n_16347;
wire n_9944;
wire n_13709;
wire n_9888;
wire n_10844;
wire n_4710;
wire n_17040;
wire n_19696;
wire n_19041;
wire n_15267;
wire n_4326;
wire n_15455;
wire n_2121;
wire n_10242;
wire n_16023;
wire n_20637;
wire n_4685;
wire n_9936;
wire n_19201;
wire n_2068;
wire n_17198;
wire n_10727;
wire n_6194;
wire n_1454;
wire n_11231;
wire n_3396;
wire n_17296;
wire n_15944;
wire n_11448;
wire n_12227;
wire n_10679;
wire n_12282;
wire n_452;
wire n_5693;
wire n_17439;
wire n_18866;
wire n_20952;
wire n_14365;
wire n_8304;
wire n_20519;
wire n_6318;
wire n_11940;
wire n_11348;
wire n_17408;
wire n_13613;
wire n_19470;
wire n_6805;
wire n_17846;
wire n_409;
wire n_19332;
wire n_5584;
wire n_3802;
wire n_13326;
wire n_6248;
wire n_6541;
wire n_848;
wire n_4733;
wire n_161;
wire n_18243;
wire n_1814;
wire n_19579;
wire n_10526;
wire n_11439;
wire n_4041;
wire n_4208;
wire n_4623;
wire n_11462;
wire n_19096;
wire n_9676;
wire n_4935;
wire n_4004;
wire n_8650;
wire n_11272;
wire n_12989;
wire n_16005;
wire n_7767;
wire n_19805;
wire n_21050;
wire n_4194;
wire n_11759;
wire n_17760;
wire n_2602;
wire n_17001;
wire n_11061;
wire n_8284;
wire n_6481;
wire n_11478;
wire n_5633;
wire n_18847;
wire n_12200;
wire n_6991;
wire n_13863;
wire n_7434;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_13926;
wire n_11748;
wire n_17110;
wire n_9135;
wire n_9776;
wire n_17364;
wire n_20919;
wire n_15673;
wire n_11867;
wire n_14678;
wire n_17290;
wire n_10286;
wire n_4996;
wire n_9107;
wire n_18188;
wire n_9548;
wire n_15117;
wire n_7651;
wire n_20866;
wire n_18899;
wire n_1494;
wire n_1893;
wire n_18198;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_15594;
wire n_17748;
wire n_3294;
wire n_2443;
wire n_185;
wire n_7536;
wire n_5513;
wire n_14671;
wire n_19863;
wire n_10441;
wire n_2843;
wire n_18574;
wire n_20498;
wire n_11764;
wire n_7671;
wire n_15924;
wire n_8033;
wire n_17333;
wire n_15021;
wire n_5834;
wire n_20863;
wire n_3109;
wire n_13418;
wire n_16358;
wire n_10628;
wire n_20499;
wire n_11787;
wire n_11539;
wire n_10134;
wire n_19761;
wire n_6209;
wire n_4672;
wire n_20034;
wire n_3558;
wire n_13489;
wire n_15225;
wire n_18941;
wire n_3034;
wire n_10317;
wire n_15238;
wire n_16713;
wire n_14821;
wire n_7413;
wire n_19045;
wire n_7821;
wire n_14238;
wire n_3963;
wire n_13032;
wire n_6274;
wire n_4496;
wire n_12269;
wire n_16962;
wire n_14556;
wire n_936;
wire n_19185;
wire n_13901;
wire n_17850;
wire n_6237;
wire n_13635;
wire n_6802;
wire n_18329;
wire n_19251;
wire n_8028;
wire n_2794;
wire n_3940;
wire n_14343;
wire n_14217;
wire n_10379;
wire n_15094;
wire n_3473;
wire n_20297;
wire n_13278;
wire n_11081;
wire n_20862;
wire n_6716;
wire n_15519;
wire n_5388;
wire n_11230;
wire n_7470;
wire n_12206;
wire n_6203;
wire n_14468;
wire n_20789;
wire n_6899;
wire n_7980;
wire n_19112;
wire n_3360;
wire n_17111;
wire n_3585;
wire n_9025;
wire n_19446;
wire n_2000;
wire n_4037;
wire n_14675;
wire n_4659;
wire n_13962;
wire n_5196;
wire n_20880;
wire n_10382;
wire n_19772;
wire n_14235;
wire n_19269;
wire n_17226;
wire n_9660;
wire n_5763;
wire n_19323;
wire n_13018;
wire n_12739;
wire n_1235;
wire n_2584;
wire n_15031;
wire n_1064;
wire n_633;
wire n_16758;
wire n_16436;
wire n_9902;
wire n_19477;
wire n_18934;
wire n_11397;
wire n_16601;
wire n_8726;
wire n_8977;
wire n_7018;
wire n_18047;
wire n_18840;
wire n_15248;
wire n_3258;
wire n_20006;
wire n_10691;
wire n_12650;
wire n_10764;
wire n_6174;
wire n_14690;
wire n_15116;
wire n_20559;
wire n_7297;
wire n_18539;
wire n_12279;
wire n_17027;
wire n_6013;
wire n_19207;
wire n_2987;
wire n_6279;
wire n_19173;
wire n_9588;
wire n_2651;
wire n_19851;
wire n_2733;
wire n_2103;
wire n_3316;
wire n_10071;
wire n_18553;
wire n_19459;
wire n_12588;
wire n_20731;
wire n_6131;
wire n_5384;
wire n_19730;
wire n_6477;
wire n_7486;
wire n_840;
wire n_6575;
wire n_11719;
wire n_20826;
wire n_19854;
wire n_5283;
wire n_17631;
wire n_15810;
wire n_8724;
wire n_12775;
wire n_17916;
wire n_6252;
wire n_14031;
wire n_12167;
wire n_8253;
wire n_15033;
wire n_4414;
wire n_14918;
wire n_9598;
wire n_10436;
wire n_228;
wire n_6668;
wire n_20123;
wire n_9311;
wire n_11982;
wire n_3445;
wire n_14448;
wire n_11522;
wire n_4087;
wire n_1684;
wire n_1148;
wire n_19149;
wire n_4619;
wire n_17043;
wire n_4398;
wire n_16316;
wire n_5350;
wire n_14906;
wire n_14187;
wire n_2429;
wire n_6779;
wire n_9608;
wire n_4449;
wire n_4607;
wire n_5949;
wire n_10515;
wire n_20427;
wire n_13713;
wire n_2971;
wire n_19802;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_20936;
wire n_19061;
wire n_20207;
wire n_8823;
wire n_8536;
wire n_17810;
wire n_20565;
wire n_5856;
wire n_7747;
wire n_14263;
wire n_12404;
wire n_4415;
wire n_18396;
wire n_1964;
wire n_14872;
wire n_7552;
wire n_18783;
wire n_9537;
wire n_19870;
wire n_9421;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_199;
wire n_14775;
wire n_4947;
wire n_2545;
wire n_15124;
wire n_8259;
wire n_12274;
wire n_4976;
wire n_11183;
wire n_9469;
wire n_17545;
wire n_4548;
wire n_7819;
wire n_15680;
wire n_3556;
wire n_4574;
wire n_8160;
wire n_20939;
wire n_2644;
wire n_10631;
wire n_10864;
wire n_1698;
wire n_18730;
wire n_5548;
wire n_13477;
wire n_1168;
wire n_10748;
wire n_5840;
wire n_3296;
wire n_9909;
wire n_15087;
wire n_3794;
wire n_19273;
wire n_656;
wire n_20267;
wire n_18517;
wire n_3293;
wire n_4902;
wire n_12002;
wire n_10751;
wire n_7794;
wire n_16311;
wire n_3934;
wire n_16846;
wire n_17377;
wire n_13987;
wire n_20106;
wire n_6965;
wire n_17670;
wire n_1846;
wire n_15607;
wire n_16731;
wire n_4161;
wire n_14673;
wire n_15943;
wire n_757;
wire n_6284;
wire n_17471;
wire n_14393;
wire n_5321;
wire n_18723;
wire n_9366;
wire n_5915;
wire n_9647;
wire n_17890;
wire n_20133;
wire n_7753;
wire n_12304;
wire n_1313;
wire n_4716;
wire n_14760;
wire n_8948;
wire n_13541;
wire n_18892;
wire n_13551;
wire n_15131;
wire n_20510;
wire n_11634;
wire n_19325;
wire n_2830;
wire n_4757;
wire n_6760;
wire n_4591;
wire n_9102;
wire n_7014;
wire n_2491;
wire n_13902;
wire n_5337;
wire n_1820;
wire n_10013;
wire n_17497;
wire n_7160;
wire n_18400;
wire n_16099;
wire n_20703;
wire n_19920;
wire n_15986;
wire n_6046;
wire n_16896;
wire n_21085;
wire n_8919;
wire n_20107;
wire n_6091;
wire n_1635;
wire n_8440;
wire n_18436;
wire n_15102;
wire n_4896;
wire n_17580;
wire n_4851;
wire n_9860;
wire n_17238;
wire n_9670;
wire n_13903;
wire n_15868;
wire n_5605;
wire n_15905;
wire n_1938;
wire n_13080;
wire n_17634;
wire n_16729;
wire n_5753;
wire n_15681;
wire n_4901;
wire n_16669;
wire n_13408;
wire n_6221;
wire n_12810;
wire n_8177;
wire n_13733;
wire n_2334;
wire n_14311;
wire n_14147;
wire n_610;
wire n_4602;
wire n_1436;
wire n_20922;
wire n_4900;
wire n_10110;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_16267;
wire n_17276;
wire n_8638;
wire n_20443;
wire n_9980;
wire n_19794;
wire n_16058;
wire n_12003;
wire n_10908;
wire n_6937;
wire n_16365;
wire n_19215;
wire n_5439;
wire n_8687;
wire n_137;
wire n_8721;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_16331;
wire n_14478;
wire n_19966;
wire n_5250;
wire n_12416;
wire n_14895;
wire n_9702;
wire n_520;
wire n_13056;
wire n_4985;
wire n_9000;
wire n_13087;
wire n_2248;
wire n_6446;
wire n_20945;
wire n_6071;
wire n_2579;
wire n_1535;
wire n_871;
wire n_8197;
wire n_18922;
wire n_12294;
wire n_15883;
wire n_14396;
wire n_339;
wire n_6178;
wire n_12786;
wire n_2221;
wire n_7550;
wire n_8554;
wire n_2442;
wire n_15756;
wire n_19246;
wire n_7292;
wire n_20705;
wire n_18787;
wire n_11471;
wire n_5098;
wire n_17402;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_8263;
wire n_5145;
wire n_13236;
wire n_2878;
wire n_11198;
wire n_14465;
wire n_3999;
wire n_17388;
wire n_13393;
wire n_7112;
wire n_868;
wire n_2458;
wire n_7971;
wire n_20925;
wire n_19298;
wire n_12802;
wire n_10633;
wire n_18010;
wire n_10573;
wire n_2859;
wire n_5216;
wire n_16983;
wire n_20504;
wire n_8474;
wire n_18271;
wire n_5703;
wire n_18965;
wire n_6886;
wire n_1636;
wire n_17648;
wire n_17617;
wire n_20283;
wire n_12296;
wire n_20867;
wire n_18418;
wire n_4546;
wire n_11288;
wire n_1254;
wire n_10570;
wire n_13151;
wire n_3073;
wire n_17558;
wire n_238;
wire n_4576;
wire n_5995;
wire n_17698;
wire n_11456;
wire n_19411;
wire n_8144;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_3136;
wire n_15320;
wire n_20475;
wire n_5330;
wire n_13935;
wire n_9351;
wire n_13930;
wire n_17076;
wire n_10106;
wire n_16338;
wire n_16811;
wire n_16747;
wire n_6345;
wire n_9242;
wire n_15303;
wire n_15598;
wire n_11821;
wire n_9522;
wire n_14560;
wire n_12488;
wire n_14028;
wire n_11395;
wire n_10387;
wire n_6291;
wire n_10615;
wire n_2595;
wire n_10790;
wire n_1465;
wire n_10555;
wire n_12896;
wire n_7123;
wire n_14670;
wire n_17145;
wire n_3860;
wire n_10222;
wire n_2909;
wire n_10671;
wire n_225;
wire n_15747;
wire n_19779;
wire n_546;
wire n_13292;
wire n_15250;
wire n_1159;
wire n_9662;
wire n_1669;
wire n_2969;
wire n_9768;
wire n_1675;
wire n_15934;
wire n_19381;
wire n_17868;
wire n_17870;
wire n_20477;
wire n_1935;
wire n_10255;
wire n_8742;
wire n_9835;
wire n_11643;
wire n_12618;
wire n_14604;
wire n_9475;
wire n_18721;
wire n_1351;
wire n_18800;
wire n_20712;
wire n_17455;
wire n_17232;
wire n_4850;
wire n_10007;
wire n_12127;
wire n_13651;
wire n_16614;
wire n_15773;
wire n_7157;
wire n_21073;
wire n_4937;
wire n_18072;
wire n_15012;
wire n_13678;
wire n_8310;
wire n_11212;
wire n_10552;
wire n_19414;
wire n_19654;
wire n_6042;
wire n_18902;
wire n_8238;
wire n_5203;
wire n_16443;
wire n_17418;
wire n_16408;
wire n_16359;
wire n_7091;
wire n_9833;
wire n_19330;
wire n_3159;
wire n_15560;
wire n_14590;
wire n_9861;
wire n_15526;
wire n_19678;
wire n_20638;
wire n_2848;
wire n_16534;
wire n_8943;
wire n_18570;
wire n_18434;
wire n_18841;
wire n_10376;
wire n_13617;
wire n_6970;
wire n_1026;
wire n_16476;
wire n_14956;
wire n_14509;
wire n_16299;
wire n_5408;
wire n_11278;
wire n_14692;
wire n_8758;
wire n_11671;
wire n_20165;
wire n_16882;
wire n_8544;
wire n_18877;
wire n_7087;
wire n_967;
wire n_10027;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_13597;
wire n_20719;
wire n_1079;
wire n_20651;
wire n_9235;
wire n_15822;
wire n_3393;
wire n_17743;
wire n_20792;
wire n_17436;
wire n_12423;
wire n_11372;
wire n_15219;
wire n_2172;
wire n_2601;
wire n_18437;
wire n_17083;
wire n_20959;
wire n_19904;
wire n_8999;
wire n_3629;
wire n_18957;
wire n_7713;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_21059;
wire n_15770;
wire n_11155;
wire n_3287;
wire n_11714;
wire n_12293;
wire n_13947;
wire n_16433;
wire n_3046;
wire n_2921;
wire n_3980;
wire n_3257;
wire n_18647;
wire n_21044;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_3979;
wire n_13648;
wire n_19180;
wire n_2695;
wire n_13274;
wire n_4003;
wire n_1832;
wire n_13472;
wire n_9397;
wire n_20201;
wire n_13870;
wire n_16278;
wire n_20249;
wire n_12000;
wire n_6799;
wire n_9767;
wire n_12903;
wire n_2274;
wire n_19846;
wire n_5640;
wire n_20044;
wire n_16007;
wire n_7298;
wire n_2768;
wire n_351;
wire n_17621;
wire n_12895;
wire n_7641;
wire n_19744;
wire n_5905;
wire n_2728;
wire n_5159;
wire n_19843;
wire n_9310;
wire n_16976;
wire n_8446;
wire n_1058;
wire n_20313;
wire n_7616;
wire n_5231;
wire n_19890;
wire n_15495;
wire n_564;
wire n_10837;
wire n_19759;
wire n_12664;
wire n_7271;
wire n_9055;
wire n_13311;
wire n_1689;
wire n_8605;
wire n_3031;
wire n_19343;
wire n_14766;
wire n_6930;
wire n_5482;
wire n_11098;
wire n_3215;
wire n_8312;
wire n_16035;
wire n_2041;
wire n_13786;
wire n_1933;
wire n_13645;
wire n_17920;
wire n_18352;
wire n_12044;
wire n_346;
wire n_15440;
wire n_5651;
wire n_264;
wire n_4074;
wire n_18700;
wire n_20739;
wire n_15252;
wire n_20342;
wire n_14664;
wire n_13299;
wire n_12257;
wire n_19998;
wire n_6374;
wire n_18611;
wire n_3917;
wire n_16255;
wire n_11778;
wire n_18952;
wire n_17866;
wire n_5735;
wire n_14338;
wire n_17555;
wire n_20398;
wire n_6588;
wire n_4243;
wire n_7897;
wire n_18982;
wire n_4225;
wire n_17883;
wire n_19049;
wire n_6865;
wire n_19087;
wire n_16194;
wire n_9586;
wire n_10670;
wire n_11177;
wire n_14900;
wire n_10004;
wire n_4907;
wire n_17037;
wire n_5787;
wire n_16573;
wire n_18668;
wire n_1611;
wire n_10171;
wire n_19076;
wire n_10406;
wire n_11236;
wire n_12562;
wire n_11600;
wire n_15517;
wire n_4916;
wire n_15334;
wire n_20023;
wire n_12217;
wire n_529;
wire n_17142;
wire n_17136;
wire n_17026;
wire n_6653;
wire n_6372;
wire n_7120;
wire n_15344;
wire n_11009;
wire n_16248;
wire n_6424;
wire n_11480;
wire n_20891;
wire n_19996;
wire n_983;
wire n_20024;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_1614;
wire n_5328;
wire n_20345;
wire n_6011;
wire n_15995;
wire n_18803;
wire n_3205;
wire n_11589;
wire n_729;
wire n_13110;
wire n_1122;
wire n_2593;
wire n_2184;
wire n_16430;
wire n_8360;
wire n_6505;
wire n_18869;
wire n_9837;
wire n_17758;
wire n_2754;
wire n_17787;
wire n_20035;
wire n_6762;
wire n_16795;
wire n_16632;
wire n_15191;
wire n_11011;
wire n_4514;
wire n_7629;
wire n_10787;
wire n_6987;
wire n_3908;
wire n_11812;
wire n_18852;
wire n_6308;
wire n_13074;
wire n_10896;
wire n_18511;
wire n_11959;
wire n_16774;
wire n_13927;
wire n_18566;
wire n_20458;
wire n_19676;
wire n_6187;
wire n_735;
wire n_15436;
wire n_19289;
wire n_13810;
wire n_14452;
wire n_1294;
wire n_20199;
wire n_7479;
wire n_13607;
wire n_7517;
wire n_11283;
wire n_18093;
wire n_15668;
wire n_18253;
wire n_6149;
wire n_11191;
wire n_10137;
wire n_19741;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_18218;
wire n_5648;
wire n_11644;
wire n_11354;
wire n_842;
wire n_13537;
wire n_18618;
wire n_6547;
wire n_9524;
wire n_7177;
wire n_20997;
wire n_18371;
wire n_12623;
wire n_20978;
wire n_2742;
wire n_5762;
wire n_20054;
wire n_5484;
wire n_18514;
wire n_16391;
wire n_10019;
wire n_14135;
wire n_1895;
wire n_21090;
wire n_16221;
wire n_16457;
wire n_19478;
wire n_2008;
wire n_454;
wire n_4989;
wire n_9084;
wire n_2127;
wire n_20307;
wire n_3151;
wire n_2460;
wire n_10995;
wire n_18573;
wire n_4528;
wire n_18782;
wire n_19958;
wire n_10597;
wire n_659;
wire n_12345;
wire n_15655;
wire n_7482;
wire n_13841;
wire n_16555;
wire n_20796;
wire n_18201;
wire n_8538;
wire n_13883;
wire n_9204;
wire n_17643;
wire n_19818;
wire n_4280;
wire n_20724;
wire n_17250;
wire n_5256;
wire n_17584;
wire n_2140;
wire n_14776;
wire n_2157;
wire n_17217;
wire n_12265;
wire n_18078;
wire n_3656;
wire n_8061;
wire n_10775;
wire n_8754;
wire n_12108;
wire n_19716;
wire n_8915;
wire n_11219;
wire n_5364;
wire n_19708;
wire n_15833;
wire n_11857;
wire n_5597;
wire n_11735;
wire n_19249;
wire n_11986;
wire n_8072;
wire n_15205;
wire n_9014;
wire n_19328;
wire n_20788;
wire n_5469;
wire n_3685;
wire n_17619;
wire n_13925;
wire n_8774;
wire n_16766;
wire n_2939;
wire n_3425;
wire n_16022;
wire n_16193;
wire n_5021;
wire n_19067;
wire n_20182;
wire n_17725;
wire n_19743;
wire n_19693;
wire n_14939;
wire n_1405;
wire n_3813;
wire n_13774;
wire n_19291;
wire n_9694;
wire n_13323;
wire n_10718;
wire n_10951;
wire n_2264;
wire n_805;
wire n_19832;
wire n_18286;
wire n_16427;
wire n_3811;
wire n_190;
wire n_5785;
wire n_3411;
wire n_10655;
wire n_10942;
wire n_4938;
wire n_6114;
wire n_463;
wire n_13192;
wire n_5505;
wire n_19875;
wire n_18636;
wire n_2905;
wire n_878;
wire n_6829;
wire n_9764;
wire n_20134;
wire n_19309;
wire n_18499;
wire n_6464;
wire n_8802;
wire n_2720;
wire n_8603;
wire n_15691;
wire n_17791;
wire n_10639;
wire n_5970;
wire n_11358;
wire n_6838;
wire n_6368;
wire n_20708;
wire n_16699;
wire n_1616;
wire n_19929;
wire n_5161;
wire n_14132;
wire n_12152;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_17660;
wire n_6166;
wire n_5378;
wire n_12511;
wire n_2022;
wire n_12705;
wire n_7743;
wire n_14934;
wire n_8584;
wire n_13017;
wire n_198;
wire n_15834;
wire n_1208;
wire n_12207;
wire n_20302;
wire n_17861;
wire n_15875;
wire n_20943;
wire n_19222;
wire n_18815;
wire n_15299;
wire n_7996;
wire n_12970;
wire n_2143;
wire n_5266;
wire n_20052;
wire n_18640;
wire n_16463;
wire n_17582;
wire n_8509;
wire n_12408;
wire n_17935;
wire n_4097;
wire n_18950;
wire n_17024;
wire n_11717;
wire n_5293;
wire n_19362;
wire n_8354;
wire n_16943;
wire n_16263;
wire n_422;
wire n_18332;
wire n_8277;
wire n_4727;
wire n_16448;
wire n_11473;
wire n_18944;
wire n_1047;
wire n_10055;
wire n_12698;
wire n_17071;
wire n_4008;
wire n_13878;
wire n_17434;
wire n_2285;
wire n_3184;
wire n_8644;
wire n_11534;
wire n_2173;
wire n_10465;
wire n_21012;
wire n_19188;
wire n_7314;
wire n_10610;
wire n_8609;
wire n_9758;
wire n_12078;
wire n_8082;
wire n_4534;
wire n_12502;
wire n_271;
wire n_19828;
wire n_15614;
wire n_5697;
wire n_13763;
wire n_17756;
wire n_15737;
wire n_11785;
wire n_6727;
wire n_5911;
wire n_20573;
wire n_256;
wire n_3600;
wire n_9967;
wire n_16078;
wire n_8819;
wire n_19241;
wire n_8487;
wire n_3027;
wire n_6454;
wire n_16183;
wire n_3800;
wire n_3462;
wire n_14579;
wire n_16390;
wire n_19208;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_7004;
wire n_16900;
wire n_588;
wire n_16139;
wire n_8517;
wire n_5356;
wire n_1341;
wire n_11853;
wire n_2431;
wire n_12988;
wire n_19584;
wire n_5841;
wire n_14542;
wire n_7030;
wire n_17089;
wire n_8203;
wire n_413;
wire n_19749;
wire n_9442;
wire n_1066;
wire n_20655;
wire n_13305;
wire n_12284;
wire n_11364;
wire n_20622;
wire n_11323;
wire n_13697;
wire n_3344;
wire n_12652;
wire n_1534;
wire n_16029;
wire n_21122;
wire n_12379;
wire n_10925;
wire n_16528;
wire n_9986;
wire n_18594;
wire n_16888;
wire n_3384;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_11902;
wire n_7280;
wire n_18435;
wire n_12701;
wire n_14008;
wire n_19340;
wire n_7597;
wire n_8884;
wire n_3113;
wire n_9225;
wire n_18182;
wire n_19763;
wire n_5645;
wire n_639;
wire n_5020;
wire n_6455;
wire n_13639;
wire n_16015;
wire n_16208;
wire n_8271;
wire n_8392;
wire n_15835;
wire n_19043;
wire n_20105;
wire n_10046;
wire n_9412;
wire n_17431;
wire n_11834;
wire n_8228;
wire n_16989;
wire n_11663;
wire n_16692;
wire n_4333;
wire n_15645;
wire n_8483;
wire n_18707;
wire n_5443;
wire n_15646;
wire n_12385;
wire n_1166;
wire n_3363;
wire n_1803;
wire n_872;
wire n_15075;
wire n_19417;
wire n_4455;
wire n_18295;
wire n_9575;
wire n_11566;
wire n_12164;
wire n_6994;
wire n_10456;
wire n_15383;
wire n_12224;
wire n_11649;
wire n_13061;
wire n_21119;
wire n_2236;
wire n_18641;
wire n_16012;
wire n_20991;
wire n_8936;
wire n_10822;
wire n_8738;
wire n_18832;
wire n_9727;
wire n_2648;
wire n_6870;
wire n_3810;
wire n_19514;
wire n_8226;
wire n_15272;
wire n_6501;
wire n_2204;
wire n_11308;
wire n_2040;
wire n_20526;
wire n_2151;
wire n_6467;
wire n_2231;
wire n_5702;
wire n_9545;
wire n_16706;
wire n_3574;
wire n_2289;
wire n_9046;
wire n_9430;
wire n_1027;
wire n_5806;
wire n_4110;
wire n_9625;
wire n_8783;
wire n_6507;
wire n_10842;
wire n_15865;
wire n_4048;
wire n_9485;
wire n_4949;
wire n_2181;
wire n_18873;
wire n_18372;
wire n_9129;
wire n_1124;
wire n_11832;
wire n_7872;
wire n_1326;
wire n_2282;
wire n_20734;
wire n_981;
wire n_8671;
wire n_19780;
wire n_12095;
wire n_11744;
wire n_15817;
wire n_10057;
wire n_20571;
wire n_2858;
wire n_15141;
wire n_15181;
wire n_3410;
wire n_13372;
wire n_5415;
wire n_10739;
wire n_12327;
wire n_4820;
wire n_11875;
wire n_10878;
wire n_1482;
wire n_8522;
wire n_1520;
wire n_12030;
wire n_9457;
wire n_16786;
wire n_16354;
wire n_16821;
wire n_17184;
wire n_6608;
wire n_11400;
wire n_16073;
wire n_12291;
wire n_2385;
wire n_20051;
wire n_7925;
wire n_6359;
wire n_20045;
wire n_10583;
wire n_7093;
wire n_4177;
wire n_19970;
wire n_8356;
wire n_1385;
wire n_16146;
wire n_17559;
wire n_16781;
wire n_5029;
wire n_2675;
wire n_3521;
wire n_16268;
wire n_16037;
wire n_20368;
wire n_3855;
wire n_6353;
wire n_5218;
wire n_16271;
wire n_18222;
wire n_8736;
wire n_919;
wire n_15625;
wire n_16465;
wire n_679;
wire n_10839;
wire n_18382;
wire n_220;
wire n_10603;
wire n_19974;
wire n_20847;
wire n_16854;
wire n_1550;
wire n_1200;
wire n_16149;
wire n_12762;
wire n_11518;
wire n_5512;
wire n_16928;
wire n_13580;
wire n_17518;
wire n_15336;
wire n_15473;
wire n_8213;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_13514;
wire n_9903;
wire n_15460;
wire n_20251;
wire n_17168;
wire n_372;
wire n_15524;
wire n_18762;
wire n_4550;
wire n_9238;
wire n_4347;
wire n_968;
wire n_12495;
wire n_19766;
wire n_5611;
wire n_3278;
wire n_12790;
wire n_3608;
wire n_14924;
wire n_12106;
wire n_11130;
wire n_18152;
wire n_11053;
wire n_19919;
wire n_15881;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_19722;
wire n_18724;
wire n_18720;
wire n_5308;
wire n_4434;
wire n_13303;
wire n_5739;
wire n_10596;
wire n_7820;
wire n_8437;
wire n_15437;
wire n_20556;
wire n_12991;
wire n_9071;
wire n_21010;
wire n_5425;
wire n_19758;
wire n_2358;
wire n_20540;
wire n_13368;
wire n_1390;
wire n_10708;
wire n_5887;
wire n_13948;
wire n_7808;
wire n_9519;
wire n_15960;
wire n_13598;
wire n_14341;
wire n_11153;
wire n_3038;
wire n_10513;
wire n_16516;
wire n_8613;
wire n_19990;
wire n_3693;
wire n_20355;
wire n_5880;
wire n_5002;
wire n_5531;
wire n_17424;
wire n_1619;
wire n_17820;
wire n_12025;
wire n_12669;
wire n_3188;
wire n_10410;
wire n_16917;
wire n_20987;
wire n_19756;
wire n_2101;
wire n_17114;
wire n_1236;
wire n_14885;
wire n_13748;
wire n_14878;
wire n_19544;
wire n_19474;
wire n_1334;
wire n_18138;
wire n_6745;
wire n_7943;
wire n_16848;
wire n_4471;
wire n_11967;
wire n_8900;
wire n_6064;
wire n_488;
wire n_17210;
wire n_9051;
wire n_16352;
wire n_7904;
wire n_16687;
wire n_684;
wire n_7296;
wire n_8323;
wire n_10459;
wire n_17445;
wire n_8711;
wire n_15787;
wire n_11628;
wire n_12704;
wire n_18317;
wire n_3874;
wire n_5730;
wire n_4165;
wire n_2056;
wire n_15289;
wire n_1144;
wire n_11026;
wire n_15672;
wire n_19195;
wire n_10915;
wire n_19830;
wire n_709;
wire n_16527;
wire n_14941;
wire n_1686;
wire n_20351;
wire n_4232;
wire n_662;
wire n_3461;
wire n_15903;
wire n_17125;
wire n_10624;
wire n_7682;
wire n_10152;
wire n_6861;
wire n_2297;
wire n_12888;
wire n_7300;
wire n_12034;
wire n_19023;
wire n_11188;
wire n_9166;
wire n_7798;
wire n_13906;
wire n_16615;
wire n_8969;
wire n_19612;
wire n_11209;
wire n_948;
wire n_6528;
wire n_8896;
wire n_5144;
wire n_3072;
wire n_6523;
wire n_5169;
wire n_14618;
wire n_11469;
wire n_9363;
wire n_11971;
wire n_19042;
wire n_4698;
wire n_18384;
wire n_18879;
wire n_18150;
wire n_853;
wire n_15497;
wire n_16519;
wire n_3763;
wire n_10823;
wire n_14623;
wire n_6389;
wire n_14635;
wire n_9307;
wire n_13922;
wire n_9876;
wire n_3947;
wire n_20518;
wire n_10814;
wire n_5183;
wire n_4533;
wire n_8286;
wire n_2164;
wire n_20114;
wire n_1186;
wire n_2052;
wire n_10549;
wire n_10370;
wire n_14171;
wire n_2205;
wire n_12513;
wire n_14988;
wire n_1724;
wire n_2080;
wire n_1126;
wire n_14975;
wire n_19271;
wire n_2357;
wire n_19108;
wire n_10543;
wire n_18023;
wire n_8639;
wire n_18739;
wire n_11301;
wire n_1302;
wire n_4444;
wire n_7681;
wire n_8566;
wire n_6613;
wire n_15492;
wire n_6404;
wire n_13905;
wire n_10259;
wire n_1583;
wire n_13936;
wire n_18759;
wire n_14386;
wire n_5997;
wire n_10302;
wire n_19116;
wire n_15243;
wire n_11276;
wire n_7150;
wire n_7974;
wire n_19922;
wire n_11326;
wire n_5563;
wire n_3030;
wire n_13144;
wire n_20352;
wire n_1296;
wire n_8112;
wire n_8489;
wire n_8060;
wire n_6230;
wire n_13134;
wire n_2514;
wire n_6977;
wire n_16832;
wire n_11732;
wire n_19549;
wire n_18351;
wire n_5932;
wire n_12321;
wire n_11855;
wire n_20949;
wire n_1299;
wire n_3489;
wire n_14306;
wire n_15765;
wire n_4967;
wire n_12104;
wire n_6001;
wire n_9682;
wire n_17347;
wire n_9278;
wire n_16719;
wire n_2797;
wire n_9222;
wire n_19320;
wire n_8562;
wire n_4376;
wire n_11350;
wire n_12799;
wire n_17443;
wire n_3712;
wire n_12202;
wire n_11057;
wire n_10170;
wire n_18529;
wire n_2823;
wire n_17381;
wire n_14371;
wire n_15759;
wire n_15378;
wire n_16060;
wire n_15287;
wire n_12055;
wire n_7116;
wire n_18861;
wire n_21104;
wire n_1353;
wire n_19419;
wire n_8537;
wire n_17116;
wire n_16763;
wire n_373;
wire n_7909;
wire n_12894;
wire n_6053;
wire n_11024;
wire n_18692;
wire n_17225;
wire n_13131;
wire n_5625;
wire n_9069;
wire n_20743;
wire n_8332;
wire n_3742;
wire n_14190;
wire n_16092;
wire n_16009;
wire n_11390;
wire n_14696;
wire n_18341;
wire n_4813;
wire n_3352;
wire n_12390;
wire n_20286;
wire n_15794;
wire n_2367;
wire n_9556;
wire n_14546;
wire n_11380;
wire n_5570;
wire n_6411;
wire n_5670;
wire n_20986;
wire n_13256;
wire n_11214;
wire n_2123;
wire n_10482;
wire n_1196;
wire n_410;
wire n_9243;
wire n_10733;
wire n_15127;
wire n_8812;
wire n_6401;
wire n_9928;
wire n_7976;
wire n_16647;
wire n_19172;
wire n_19560;
wire n_945;
wire n_10641;
wire n_11115;
wire n_3665;
wire n_8062;
wire n_3281;
wire n_16690;
wire n_3535;
wire n_5061;
wire n_4653;
wire n_15431;
wire n_15491;
wire n_5978;
wire n_6853;
wire n_14938;
wire n_14427;
wire n_500;
wire n_6181;
wire n_13964;
wire n_19662;
wire n_7801;
wire n_9975;
wire n_17638;
wire n_6907;
wire n_2342;
wire n_5177;
wire n_3856;
wire n_11371;
wire n_11939;
wire n_7876;
wire n_18231;
wire n_143;
wire n_2709;
wire n_3419;
wire n_10850;
wire n_13129;
wire n_19162;
wire n_18880;
wire n_6517;
wire n_17693;
wire n_6339;
wire n_20969;
wire n_14408;
wire n_14659;
wire n_14267;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_770;
wire n_5607;
wire n_14516;
wire n_2782;
wire n_15692;
wire n_3929;
wire n_971;
wire n_19522;
wire n_8212;
wire n_18392;
wire n_1650;
wire n_6504;
wire n_9891;
wire n_4176;
wire n_9078;
wire n_13553;
wire n_7556;
wire n_10972;
wire n_6814;
wire n_7216;
wire n_5278;
wire n_2779;
wire n_19512;
wire n_21112;
wire n_3756;
wire n_12391;
wire n_8223;
wire n_16941;
wire n_4077;
wire n_17798;
wire n_18660;
wire n_12731;
wire n_13623;
wire n_432;
wire n_18771;
wire n_13775;
wire n_17258;
wire n_4839;
wire n_9174;
wire n_5969;
wire n_20019;
wire n_15609;
wire n_611;
wire n_17440;
wire n_1013;
wire n_6686;
wire n_16217;
wire n_4929;
wire n_14067;
wire n_6536;
wire n_8434;
wire n_12508;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_14614;
wire n_10898;
wire n_3913;
wire n_8608;
wire n_13583;
wire n_1230;
wire n_376;
wire n_16481;
wire n_4541;
wire n_15872;
wire n_16110;
wire n_3861;
wire n_21007;
wire n_19392;
wire n_11287;
wire n_4171;
wire n_9117;
wire n_7022;
wire n_4665;
wire n_7476;
wire n_10590;
wire n_4884;
wire n_16185;
wire n_4276;
wire n_7208;
wire n_17163;
wire n_11277;
wire n_11919;
wire n_1112;
wire n_19933;
wire n_9001;
wire n_16910;
wire n_6868;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_18996;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_10159;
wire n_5174;
wire n_9024;
wire n_10178;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_14268;
wire n_20234;
wire n_13892;
wire n_14136;
wire n_12636;
wire n_20464;
wire n_3119;
wire n_6671;
wire n_18622;
wire n_4740;
wire n_10550;
wire n_16297;
wire n_257;
wire n_16112;
wire n_5544;
wire n_18280;
wire n_9725;
wire n_8842;
wire n_16473;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_12648;
wire n_20990;
wire n_4920;
wire n_5069;
wire n_10660;
wire n_17629;
wire n_15848;
wire n_14262;
wire n_8799;
wire n_4378;
wire n_6065;
wire n_12441;
wire n_19728;
wire n_4459;
wire n_11461;
wire n_5808;
wire n_13604;
wire n_18055;
wire n_8045;
wire n_7538;
wire n_14029;
wire n_13157;
wire n_11536;
wire n_20473;
wire n_9716;
wire n_15502;
wire n_7242;
wire n_20787;
wire n_11305;
wire n_15352;
wire n_179;
wire n_2925;
wire n_1435;
wire n_8022;
wire n_8227;
wire n_2072;
wire n_10309;
wire n_5381;
wire n_15569;
wire n_436;
wire n_19301;
wire n_10021;
wire n_324;
wire n_18752;
wire n_10053;
wire n_7389;
wire n_10765;
wire n_6265;
wire n_18799;
wire n_4914;
wire n_8604;
wire n_13092;
wire n_10907;
wire n_7834;
wire n_11299;
wire n_16085;
wire n_16116;
wire n_1139;
wire n_3688;
wire n_11273;
wire n_15416;
wire n_1312;
wire n_18637;
wire n_13147;
wire n_12871;
wire n_13212;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_8995;
wire n_20818;
wire n_3666;
wire n_16370;
wire n_17011;
wire n_867;
wire n_12785;
wire n_14808;
wire n_13661;
wire n_749;
wire n_19521;
wire n_3998;
wire n_16960;
wire n_17744;
wire n_7000;
wire n_2668;
wire n_10486;
wire n_2701;
wire n_2400;
wire n_15228;
wire n_10357;
wire n_650;
wire n_3741;
wire n_9177;
wire n_2557;
wire n_5109;
wire n_1071;
wire n_5281;
wire n_19712;
wire n_13874;
wire n_2220;
wire n_7044;
wire n_16490;
wire n_6108;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_18972;
wire n_18223;
wire n_14617;
wire n_7468;
wire n_7899;
wire n_8710;
wire n_21071;
wire n_4861;
wire n_16787;
wire n_8512;
wire n_13093;
wire n_2507;
wire n_16535;
wire n_13288;
wire n_9087;
wire n_4451;
wire n_7845;
wire n_2328;
wire n_347;
wire n_2434;
wire n_15044;
wire n_16913;
wire n_9956;
wire n_20203;
wire n_19809;
wire n_4784;
wire n_14206;
wire n_13606;
wire n_19374;
wire n_12901;
wire n_10589;
wire n_11019;
wire n_15829;
wire n_14837;
wire n_6513;
wire n_14978;
wire n_16055;
wire n_2262;
wire n_4613;
wire n_9197;
wire n_11076;
wire n_9140;
wire n_8401;
wire n_370;
wire n_9364;
wire n_9398;
wire n_17279;
wire n_20898;
wire n_17601;
wire n_14321;
wire n_9203;
wire n_6381;
wire n_20104;
wire n_12054;
wire n_8450;
wire n_12081;
wire n_14095;
wire n_20046;
wire n_5929;
wire n_20849;
wire n_19238;
wire n_4242;
wire n_16324;
wire n_11860;
wire n_8104;
wire n_4122;
wire n_16265;
wire n_10919;
wire n_4522;
wire n_15350;
wire n_14077;
wire n_17721;
wire n_5956;
wire n_3267;
wire n_6017;
wire n_13011;
wire n_12737;
wire n_6125;
wire n_4932;
wire n_19313;
wire n_1384;
wire n_12092;
wire n_21078;
wire n_2983;
wire n_15017;
wire n_20172;
wire n_11451;
wire n_11816;
wire n_9500;
wire n_3513;
wire n_9747;
wire n_20527;
wire n_9470;
wire n_6414;
wire n_1068;
wire n_11232;
wire n_10188;
wire n_6936;
wire n_14373;
wire n_20539;
wire n_487;
wire n_7003;
wire n_15587;
wire n_6302;
wire n_16912;
wire n_6922;
wire n_15185;
wire n_15772;
wire n_10582;
wire n_13494;
wire n_15210;
wire n_10934;
wire n_10747;
wire n_10711;
wire n_9409;
wire n_11088;
wire n_17188;
wire n_20131;
wire n_12899;
wire n_12616;
wire n_7366;
wire n_2242;
wire n_14953;
wire n_12010;
wire n_17331;
wire n_13751;
wire n_12394;
wire n_18277;
wire n_13465;
wire n_12797;
wire n_19611;
wire n_16231;
wire n_677;
wire n_8400;
wire n_11090;
wire n_9858;
wire n_7511;
wire n_10936;
wire n_12134;
wire n_19657;
wire n_12730;
wire n_17103;
wire n_3494;
wire n_17147;
wire n_727;
wire n_3837;
wire n_545;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_9965;
wire n_6449;
wire n_10862;
wire n_14333;
wire n_13357;
wire n_8889;
wire n_5681;
wire n_3801;
wire n_2338;
wire n_12427;
wire n_1080;
wire n_11353;
wire n_18936;
wire n_19005;
wire n_6342;
wire n_6195;
wire n_17753;
wire n_6441;
wire n_11116;
wire n_17283;
wire n_20083;
wire n_17052;
wire n_1371;
wire n_17438;
wire n_4240;
wire n_20032;
wire n_2774;
wire n_11881;
wire n_2799;
wire n_8311;
wire n_15786;
wire n_4393;
wire n_6662;
wire n_9088;
wire n_9580;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_20569;
wire n_17398;
wire n_6433;
wire n_1763;
wire n_2763;
wire n_3156;
wire n_10530;
wire n_1859;
wire n_18115;
wire n_3492;
wire n_6369;
wire n_9951;
wire n_9855;
wire n_2379;
wire n_10102;
wire n_888;
wire n_12537;
wire n_12076;
wire n_19000;
wire n_15836;
wire n_16289;
wire n_7865;
wire n_1097;
wire n_14447;
wire n_16039;
wire n_4387;
wire n_19637;
wire n_20589;
wire n_14745;
wire n_9584;
wire n_17307;
wire n_9287;
wire n_534;
wire n_3186;
wire n_9490;
wire n_2594;
wire n_19233;
wire n_8867;
wire n_890;
wire n_9846;
wire n_20090;
wire n_4598;
wire n_12072;
wire n_5106;
wire n_13339;
wire n_14672;
wire n_16988;
wire n_11903;
wire n_8641;
wire n_9578;
wire n_11813;
wire n_5080;
wire n_9396;
wire n_19935;
wire n_12745;
wire n_12841;
wire n_7198;
wire n_6921;
wire n_16743;
wire n_3353;
wire n_17722;
wire n_6106;
wire n_12603;
wire n_14964;
wire n_6172;
wire n_20957;
wire n_9805;
wire n_812;
wire n_12466;
wire n_16220;
wire n_4040;
wire n_19604;
wire n_18089;
wire n_12982;
wire n_14680;
wire n_13459;
wire n_11795;
wire n_5191;
wire n_17149;
wire n_17249;
wire n_11646;
wire n_17630;
wire n_13649;
wire n_3161;
wire n_2389;
wire n_7126;
wire n_11963;
wire n_1394;
wire n_15027;
wire n_17929;
wire n_4112;
wire n_20709;
wire n_2614;
wire n_5428;
wire n_12497;
wire n_19795;
wire n_6678;
wire n_10838;
wire n_6564;
wire n_7268;
wire n_8174;
wire n_15196;
wire n_8846;
wire n_9277;
wire n_14754;
wire n_6109;
wire n_17832;
wire n_21113;
wire n_10123;
wire n_5798;
wire n_19739;
wire n_8032;
wire n_14445;
wire n_11147;
wire n_10048;
wire n_11194;
wire n_4758;
wire n_12228;
wire n_11016;
wire n_19681;
wire n_3507;
wire n_8524;
wire n_11924;
wire n_4535;
wire n_8828;
wire n_9639;
wire n_15916;
wire n_12059;
wire n_9664;
wire n_16434;
wire n_4731;
wire n_7073;
wire n_21023;
wire n_1786;
wire n_16894;
wire n_13820;
wire n_14366;
wire n_18924;
wire n_5571;
wire n_592;
wire n_20167;
wire n_10686;
wire n_1318;
wire n_14197;
wire n_8764;
wire n_14454;
wire n_11411;
wire n_8502;
wire n_6585;
wire n_7786;
wire n_10913;
wire n_8454;
wire n_4358;
wire n_20218;
wire n_9122;
wire n_1526;
wire n_12335;
wire n_19174;
wire n_2656;
wire n_4904;
wire n_19886;
wire n_20490;
wire n_14068;
wire n_943;
wire n_14019;
wire n_17541;
wire n_7624;
wire n_18595;
wire n_14397;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_2857;
wire n_14319;
wire n_19016;
wire n_3919;
wire n_14910;
wire n_16252;
wire n_5475;
wire n_1352;
wire n_7778;
wire n_20113;
wire n_2764;
wire n_20970;
wire n_2633;
wire n_5752;
wire n_14362;
wire n_14026;
wire n_8441;
wire n_1429;
wire n_14114;
wire n_2528;
wire n_18086;
wire n_18394;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_18777;
wire n_14504;
wire n_3718;
wire n_6685;
wire n_756;
wire n_1149;
wire n_9574;
wire n_12032;
wire n_3140;
wire n_8865;
wire n_19862;
wire n_10031;
wire n_6016;
wire n_15948;
wire n_1659;
wire n_15568;
wire n_5366;
wire n_5322;
wire n_12176;
wire n_13266;
wire n_11805;
wire n_7791;
wire n_10847;
wire n_14242;
wire n_16295;
wire n_15660;
wire n_12740;
wire n_396;
wire n_19132;
wire n_9372;
wire n_9657;
wire n_7656;
wire n_21000;
wire n_3635;
wire n_11725;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_9904;
wire n_17568;
wire n_20176;
wire n_15486;
wire n_8410;
wire n_1577;
wire n_11694;
wire n_17711;
wire n_4921;
wire n_11540;
wire n_4377;
wire n_16156;
wire n_1877;
wire n_9301;
wire n_16964;
wire n_2497;
wire n_20758;
wire n_5446;
wire n_597;
wire n_7456;
wire n_15426;
wire n_152;
wire n_1185;
wire n_16154;
wire n_13435;
wire n_11074;
wire n_12750;
wire n_15936;
wire n_18391;
wire n_20151;
wire n_6676;
wire n_4304;
wire n_18216;
wire n_11102;
wire n_17869;
wire n_10088;
wire n_19894;
wire n_16251;
wire n_7525;
wire n_19396;
wire n_17570;
wire n_16924;
wire n_5351;
wire n_19557;
wire n_11852;
wire n_12500;
wire n_19093;
wire n_15958;
wire n_276;
wire n_19157;
wire n_11684;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_12112;
wire n_19957;
wire n_4291;
wire n_20216;
wire n_2036;
wire n_10887;
wire n_3358;
wire n_1128;
wire n_9346;
wire n_2419;
wire n_11041;
wire n_10742;
wire n_12614;
wire n_9968;
wire n_18760;
wire n_6162;
wire n_2309;
wire n_16315;
wire n_4855;
wire n_3289;
wire n_6127;
wire n_305;
wire n_10328;
wire n_10692;
wire n_15118;
wire n_6126;
wire n_1549;
wire n_15592;
wire n_10206;
wire n_7844;
wire n_16377;
wire n_20268;
wire n_1362;
wire n_9509;
wire n_20872;
wire n_3123;
wire n_18215;
wire n_14239;
wire n_2645;
wire n_2749;
wire n_15710;
wire n_20822;
wire n_18910;
wire n_1885;
wire n_3251;
wire n_6723;
wire n_3723;
wire n_13251;
wire n_12107;
wire n_13504;
wire n_13521;
wire n_16886;
wire n_3242;
wire n_13161;
wire n_7011;
wire n_14076;
wire n_6393;
wire n_12380;
wire n_8916;
wire n_18239;
wire n_613;
wire n_13309;
wire n_5465;
wire n_5154;
wire n_8018;
wire n_1767;
wire n_1973;
wire n_18616;
wire n_20494;
wire n_254;
wire n_7701;
wire n_16419;
wire n_4384;
wire n_16712;
wire n_1664;
wire n_4577;
wire n_7683;
wire n_532;
wire n_7669;
wire n_8298;
wire n_15802;
wire n_6438;
wire n_1857;
wire n_17047;
wire n_17878;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_621;
wire n_16969;
wire n_8053;
wire n_11407;
wire n_18032;
wire n_1311;
wire n_15840;
wire n_697;
wire n_9528;
wire n_17023;
wire n_4620;
wire n_14379;
wire n_4924;
wire n_4044;
wire n_15999;
wire n_3304;
wire n_10772;
wire n_7362;
wire n_17881;
wire n_14942;
wire n_7082;
wire n_8988;
wire n_3247;
wire n_10664;
wire n_17818;
wire n_16204;
wire n_13380;
wire n_8893;
wire n_20483;
wire n_5805;
wire n_11910;
wire n_3785;
wire n_5501;
wire n_13188;
wire n_14179;
wire n_7386;
wire n_15259;
wire n_11361;
wire n_11894;
wire n_3178;
wire n_19063;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_15521;
wire n_20568;
wire n_14995;
wire n_7404;
wire n_17113;
wire n_6147;
wire n_6765;
wire n_19946;
wire n_4792;
wire n_3537;
wire n_14252;
wire n_14851;
wire n_191;
wire n_19266;
wire n_11623;
wire n_15394;
wire n_8712;
wire n_6352;
wire n_11124;
wire n_2941;
wire n_10448;
wire n_15100;
wire n_10301;
wire n_11977;
wire n_15487;
wire n_17981;
wire n_10074;
wire n_5562;
wire n_6093;
wire n_10001;
wire n_14944;
wire n_17768;
wire n_7877;
wire n_7787;
wire n_15578;
wire n_13961;
wire n_13343;
wire n_12546;
wire n_987;
wire n_19806;
wire n_19613;
wire n_4673;
wire n_18951;
wire n_18750;
wire n_9387;
wire n_14512;
wire n_21027;
wire n_2639;
wire n_20797;
wire n_16835;
wire n_2603;
wire n_8892;
wire n_1167;
wire n_10674;
wire n_19412;
wire n_7563;
wire n_14850;
wire n_1926;
wire n_14531;
wire n_13740;
wire n_19146;
wire n_17420;
wire n_11549;
wire n_14437;
wire n_1738;
wire n_8941;
wire n_406;
wire n_7103;
wire n_10724;
wire n_14409;
wire n_18875;
wire n_2321;
wire n_1077;
wire n_6832;
wire n_12604;
wire n_9391;
wire n_16594;
wire n_765;
wire n_4092;
wire n_18541;
wire n_12558;
wire n_15503;
wire n_4255;
wire n_385;
wire n_12840;
wire n_20977;
wire n_10863;
wire n_10958;
wire n_2186;
wire n_16335;
wire n_10174;
wire n_4647;
wire n_13960;
wire n_12435;
wire n_7134;
wire n_18118;
wire n_3042;
wire n_8288;
wire n_15891;
wire n_14629;
wire n_14778;
wire n_14010;
wire n_10403;
wire n_11972;
wire n_9834;
wire n_9901;
wire n_7102;
wire n_10015;
wire n_5271;
wire n_17579;
wire n_17140;
wire n_733;
wire n_6651;
wire n_3838;
wire n_6289;
wire n_19307;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_19449;
wire n_20219;
wire n_4499;
wire n_17585;
wire n_4504;
wire n_20579;
wire n_10460;
wire n_14265;
wire n_3598;
wire n_835;
wire n_20725;
wire n_6186;
wire n_20179;
wire n_2641;
wire n_13490;
wire n_2580;
wire n_14836;
wire n_401;
wire n_13381;
wire n_9436;
wire n_20185;
wire n_11385;
wire n_1459;
wire n_13204;
wire n_18977;
wire n_9239;
wire n_4833;
wire n_3394;
wire n_18605;
wire n_11777;
wire n_18269;
wire n_8614;
wire n_8242;
wire n_4564;
wire n_15826;
wire n_3581;
wire n_8110;
wire n_14204;
wire n_19004;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_4080;
wire n_2206;
wire n_10327;
wire n_6766;
wire n_17714;
wire n_1320;
wire n_14157;
wire n_4981;
wire n_11651;
wire n_2347;
wire n_4676;
wire n_20436;
wire n_18617;
wire n_7519;
wire n_1934;
wire n_2577;
wire n_11196;
wire n_18281;
wire n_14933;
wire n_1576;
wire n_8468;
wire n_9031;
wire n_12910;
wire n_17639;
wire n_11084;
wire n_8933;
wire n_3952;
wire n_18074;
wire n_7884;
wire n_17785;
wire n_539;
wire n_10586;
wire n_8283;
wire n_977;
wire n_2532;
wire n_7344;
wire n_5859;
wire n_14104;
wire n_7892;
wire n_19548;
wire n_18500;
wire n_11918;
wire n_13460;
wire n_18769;
wire n_12712;
wire n_15494;
wire n_10961;
wire n_6175;
wire n_11077;
wire n_18501;
wire n_809;
wire n_3032;
wire n_16207;
wire n_12209;
wire n_14494;
wire n_14168;
wire n_910;
wire n_13452;
wire n_4964;
wire n_10180;
wire n_217;
wire n_18865;
wire n_20175;
wire n_11845;
wire n_1199;
wire n_13671;
wire n_1273;
wire n_15839;
wire n_19596;
wire n_5495;
wire n_17596;
wire n_4483;
wire n_3061;
wire n_15884;
wire n_15708;
wire n_5121;
wire n_8333;
wire n_9097;
wire n_4487;
wire n_20894;
wire n_11529;
wire n_9925;
wire n_15139;
wire n_4808;
wire n_13173;
wire n_3902;
wire n_12830;
wire n_3244;
wire n_11384;
wire n_14382;
wire n_10111;
wire n_5301;
wire n_13263;
wire n_17512;
wire n_3488;
wire n_14707;
wire n_2744;
wire n_14530;
wire n_599;
wire n_13848;
wire n_6982;
wire n_537;
wire n_991;
wire n_2275;
wire n_8832;
wire n_4606;
wire n_14999;
wire n_17503;
wire n_2029;
wire n_938;
wire n_14275;
wire n_5348;
wire n_16564;
wire n_13818;
wire n_313;
wire n_20877;
wire n_378;
wire n_12845;
wire n_4465;
wire n_20287;
wire n_15764;
wire n_5558;
wire n_12047;
wire n_3725;
wire n_10190;
wire n_20555;
wire n_17230;
wire n_9534;
wire n_15274;
wire n_17685;
wire n_5520;
wire n_19718;
wire n_17728;
wire n_16127;
wire n_7554;
wire n_16550;
wire n_18241;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_1725;
wire n_14819;
wire n_1722;
wire n_11017;
wire n_11307;
wire n_4014;
wire n_2255;
wire n_12811;
wire n_13346;
wire n_13331;
wire n_5135;
wire n_16071;
wire n_13307;
wire n_19119;
wire n_1662;
wire n_19829;
wire n_6621;
wire n_4701;
wire n_782;
wire n_11193;
wire n_4869;
wire n_13939;
wire n_5533;
wire n_1796;
wire n_14429;
wire n_14098;
wire n_13289;
wire n_10247;
wire n_2876;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_14490;
wire n_18532;
wire n_20285;
wire n_12801;
wire n_21052;
wire n_20524;
wire n_18857;
wire n_11762;
wire n_14030;
wire n_19383;
wire n_7156;
wire n_8629;
wire n_8186;
wire n_1486;
wire n_15082;
wire n_17746;
wire n_13366;
wire n_19124;
wire n_20082;
wire n_4013;
wire n_6122;
wire n_4085;
wire n_14814;
wire n_6570;
wire n_9445;
wire n_18591;
wire n_8282;
wire n_7516;
wire n_6928;
wire n_20726;
wire n_20013;
wire n_16569;
wire n_187;
wire n_11314;
wire n_18733;
wire n_19703;
wire n_12210;
wire n_18059;
wire n_10130;
wire n_8183;
wire n_5065;
wire n_13450;
wire n_15752;
wire n_10956;
wire n_15389;
wire n_11515;
wire n_2013;
wire n_2786;
wire n_11490;
wire n_4058;
wire n_4819;
wire n_6835;
wire n_2436;
wire n_15813;
wire n_6269;
wire n_7970;
wire n_1706;
wire n_2461;
wire n_7154;
wire n_17441;
wire n_634;
wire n_18748;
wire n_20815;
wire n_12573;
wire n_20393;
wire n_11374;
wire n_14519;
wire n_18144;
wire n_7194;
wire n_5173;
wire n_17958;
wire n_11771;
wire n_13431;
wire n_14507;
wire n_14020;
wire n_3797;
wire n_3416;
wire n_5861;
wire n_20522;
wire n_20716;
wire n_10855;
wire n_6320;
wire n_16680;
wire n_6316;
wire n_8619;
wire n_419;
wire n_7068;
wire n_13227;
wire n_2156;
wire n_8162;
wire n_20914;
wire n_18292;
wire n_9576;
wire n_20720;
wire n_12240;
wire n_13045;
wire n_13620;
wire n_4702;
wire n_16376;
wire n_10992;
wire n_4491;
wire n_6752;
wire n_19356;
wire n_9704;
wire n_18005;
wire n_17034;
wire n_7317;
wire n_18173;
wire n_11912;
wire n_13862;
wire n_15204;
wire n_1688;
wire n_5827;
wire n_16141;
wire n_16919;
wire n_19675;
wire n_7384;
wire n_11379;
wire n_7512;
wire n_1718;
wire n_12276;
wire n_200;
wire n_10029;
wire n_14271;
wire n_13595;
wire n_5555;
wire n_2078;
wire n_8886;
wire n_11899;
wire n_20448;
wire n_1195;
wire n_15705;
wire n_15574;
wire n_7090;
wire n_8202;
wire n_13633;
wire n_1847;
wire n_12118;
wire n_10599;
wire n_18484;
wire n_5084;
wire n_17956;
wire n_8668;
wire n_884;
wire n_18935;
wire n_13528;
wire n_6796;
wire n_8979;
wire n_14064;
wire n_15550;
wire n_13456;
wire n_10947;
wire n_18926;
wire n_10386;
wire n_3793;
wire n_8199;
wire n_16918;
wire n_10267;
wire n_17845;
wire n_929;
wire n_10401;
wire n_15666;
wire n_15511;
wire n_15933;
wire n_18477;
wire n_11127;
wire n_9688;
wire n_2427;
wire n_3613;
wire n_7388;
wire n_10428;
wire n_19606;
wire n_6489;
wire n_9023;
wire n_2769;
wire n_7849;
wire n_3013;
wire n_4572;
wire n_7417;
wire n_3962;
wire n_12312;
wire n_6038;
wire n_6245;
wire n_6030;
wire n_1544;
wire n_12580;
wire n_5588;
wire n_9993;
wire n_1354;
wire n_17480;
wire n_6583;
wire n_10545;
wire n_7859;
wire n_3449;
wire n_20782;
wire n_4854;
wire n_18620;
wire n_491;
wire n_1595;
wire n_8017;
wire n_5477;
wire n_17134;
wire n_2727;
wire n_17662;
wire n_9184;
wire n_16974;
wire n_7576;
wire n_10779;
wire n_11554;
wire n_14647;
wire n_16162;
wire n_11197;
wire n_14286;
wire n_15305;
wire n_9505;
wire n_19413;
wire n_12986;
wire n_17996;
wire n_17575;
wire n_6973;
wire n_19314;
wire n_20363;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_13691;
wire n_1838;
wire n_11341;
wire n_287;
wire n_1716;
wire n_12741;
wire n_3562;
wire n_17395;
wire n_7081;
wire n_7742;
wire n_6280;
wire n_20312;
wire n_15152;
wire n_13155;
wire n_14581;
wire n_1179;
wire n_18370;
wire n_6256;
wire n_12412;
wire n_12677;
wire n_7842;
wire n_9415;
wire n_10298;
wire n_18429;
wire n_13194;
wire n_8714;
wire n_19651;
wire n_14920;
wire n_9990;
wire n_3885;
wire n_19746;
wire n_17273;
wire n_19847;
wire n_13446;
wire n_10235;
wire n_3250;
wire n_14141;
wire n_3915;
wire n_5694;
wire n_3717;
wire n_17334;
wire n_11541;
wire n_4206;
wire n_4099;
wire n_11680;
wire n_12686;
wire n_2922;
wire n_20534;
wire n_2871;
wire n_12734;
wire n_5580;
wire n_15870;
wire n_337;
wire n_12331;
wire n_3937;
wire n_4763;
wire n_18088;
wire n_9339;
wire n_11596;
wire n_17320;
wire n_18315;
wire n_6243;
wire n_10266;
wire n_5561;
wire n_7051;
wire n_18348;
wire n_10290;
wire n_2439;
wire n_20284;
wire n_19240;
wire n_5430;
wire n_16890;
wire n_824;
wire n_11839;
wire n_9279;
wire n_18297;
wire n_15354;
wire n_18728;
wire n_19918;
wire n_11548;
wire n_13515;
wire n_15583;
wire n_470;
wire n_477;
wire n_15941;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_19924;
wire n_16504;
wire n_18024;
wire n_14574;
wire n_2682;
wire n_5854;
wire n_5585;
wire n_16693;
wire n_20828;
wire n_1627;
wire n_14014;
wire n_10220;
wire n_5783;
wire n_6837;
wire n_15696;
wire n_13467;
wire n_13245;
wire n_1731;
wire n_7894;
wire n_1147;
wire n_12892;
wire n_2213;
wire n_7121;
wire n_12448;
wire n_6410;
wire n_15180;
wire n_20907;
wire n_7961;
wire n_1674;
wire n_9920;
wire n_6574;
wire n_5299;
wire n_4484;
wire n_8863;
wire n_15551;
wire n_4517;
wire n_2069;
wire n_19487;
wire n_8705;
wire n_2287;
wire n_9815;
wire n_3415;
wire n_10820;
wire n_6646;
wire n_3414;
wire n_7928;
wire n_760;
wire n_10168;
wire n_11664;
wire n_20325;
wire n_598;
wire n_3889;
wire n_14782;
wire n_3262;
wire n_5319;
wire n_15358;
wire n_13940;
wire n_261;
wire n_19975;
wire n_6028;
wire n_11006;
wire n_8729;
wire n_6682;
wire n_12593;
wire n_20116;
wire n_13873;
wire n_13335;
wire n_15458;
wire n_7797;
wire n_9267;
wire n_6216;
wire n_3660;
wire n_11831;
wire n_16553;
wire n_16665;
wire n_8478;
wire n_19699;
wire n_4978;
wire n_14256;
wire n_9419;
wire n_3299;
wire n_905;
wire n_14922;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_3876;
wire n_8276;
wire n_16546;
wire n_14862;
wire n_15915;
wire n_8706;
wire n_18134;
wire n_6167;
wire n_12357;
wire n_3642;
wire n_10750;
wire n_8532;
wire n_18383;
wire n_16134;
wire n_17654;
wire n_5731;
wire n_20558;
wire n_14105;
wire n_15727;
wire n_18705;
wire n_1879;
wire n_20457;
wire n_17248;
wire n_20290;
wire n_20444;
wire n_17925;
wire n_7725;
wire n_18969;
wire n_3572;
wire n_3471;
wire n_1484;
wire n_11585;
wire n_6217;
wire n_3118;
wire n_9157;
wire n_5560;
wire n_20371;
wire n_16396;
wire n_4441;
wire n_16445;
wire n_20211;
wire n_11001;
wire n_16951;
wire n_10196;
wire n_4458;
wire n_14547;
wire n_3831;
wire n_13904;
wire n_13944;
wire n_15935;
wire n_13359;
wire n_18598;
wire n_11063;
wire n_5781;
wire n_9368;
wire n_3443;
wire n_14201;
wire n_8329;
wire n_6370;
wire n_1726;
wire n_10329;
wire n_19774;
wire n_3996;
wire n_16349;
wire n_4771;
wire n_21061;
wire n_1098;
wire n_13609;
wire n_13817;
wire n_9422;
wire n_18938;
wire n_12619;
wire n_12541;
wire n_3951;
wire n_13428;
wire n_19563;
wire n_9338;
wire n_8125;
wire n_4236;
wire n_3290;
wire n_6712;
wire n_19667;
wire n_11757;
wire n_20883;
wire n_18305;
wire n_17028;
wire n_6465;
wire n_5673;
wire n_861;
wire n_11519;
wire n_19588;
wire n_14571;
wire n_19639;
wire n_8615;
wire n_18395;
wire n_1666;
wire n_20971;
wire n_5103;
wire n_12191;
wire n_10207;
wire n_20009;
wire n_20909;
wire n_17138;
wire n_13998;
wire n_262;
wire n_11928;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9393;
wire n_6940;
wire n_14833;
wire n_17346;
wire n_14398;
wire n_19156;
wire n_12318;
wire n_14731;
wire n_4269;
wire n_7540;
wire n_13632;
wire n_15132;
wire n_10437;
wire n_19144;
wire n_16044;
wire n_13444;
wire n_21019;
wire n_12805;
wire n_2124;
wire n_8155;
wire n_9334;
wire n_14059;
wire n_6483;
wire n_7770;
wire n_16536;
wire n_10480;
wire n_5357;
wire n_10892;
wire n_10796;
wire n_15895;
wire n_3648;
wire n_16775;
wire n_9254;
wire n_7173;
wire n_20937;
wire n_1975;
wire n_5421;
wire n_11250;
wire n_16425;
wire n_16106;
wire n_19318;
wire n_8026;
wire n_11428;
wire n_18054;
wire n_10495;
wire n_1890;
wire n_12678;
wire n_10812;
wire n_4034;
wire n_14211;
wire n_11674;
wire n_11097;
wire n_14155;
wire n_12194;
wire n_16406;
wire n_3649;
wire n_16724;
wire n_7212;
wire n_12351;
wire n_7951;
wire n_14111;
wire n_10702;
wire n_10490;
wire n_862;
wire n_7444;
wire n_2637;
wire n_2071;
wire n_430;
wire n_13571;
wire n_2082;
wire n_10906;
wire n_1532;
wire n_10891;
wire n_15019;
wire n_20704;
wire n_12036;
wire n_9554;
wire n_16417;
wire n_16796;
wire n_9315;
wire n_16776;
wire n_11201;
wire n_1060;
wire n_9999;
wire n_4424;
wire n_6543;
wire n_3400;
wire n_20272;
wire n_18081;
wire n_8083;
wire n_14596;
wire n_8057;
wire n_19950;
wire n_1783;
wire n_19939;
wire n_17593;
wire n_17924;
wire n_4646;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_19493;
wire n_4035;
wire n_3670;
wire n_8366;
wire n_10342;
wire n_10435;
wire n_14584;
wire n_19261;
wire n_18780;
wire n_20691;
wire n_5013;
wire n_19937;
wire n_20639;
wire n_13208;
wire n_16010;
wire n_17222;
wire n_19993;
wire n_3524;
wire n_7560;
wire n_4717;
wire n_6888;
wire n_17369;
wire n_602;
wire n_5424;
wire n_15627;
wire n_20137;
wire n_4750;
wire n_10978;
wire n_13880;
wire n_2667;
wire n_19734;
wire n_3746;
wire n_7731;
wire n_13050;
wire n_1046;
wire n_10816;
wire n_13133;
wire n_18490;
wire n_6854;
wire n_7940;
wire n_6793;
wire n_11930;
wire n_421;
wire n_11269;
wire n_12539;
wire n_13358;
wire n_12758;
wire n_9438;
wire n_1556;
wire n_7537;
wire n_5345;
wire n_14875;
wire n_15920;
wire n_17061;
wire n_19573;
wire n_1971;
wire n_3448;
wire n_14057;
wire n_19583;
wire n_16500;
wire n_9313;
wire n_605;
wire n_4330;
wire n_4152;
wire n_6874;
wire n_14079;
wire n_18285;
wire n_15489;
wire n_15340;
wire n_5537;
wire n_17321;
wire n_17423;
wire n_4783;
wire n_3017;
wire n_10753;
wire n_5409;
wire n_15783;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_5142;
wire n_19304;
wire n_6039;
wire n_17834;
wire n_5010;
wire n_7226;
wire n_4052;
wire n_3357;
wire n_9882;
wire n_20881;
wire n_11873;
wire n_18077;
wire n_16959;
wire n_18968;
wire n_4404;
wire n_151;
wire n_7906;
wire n_2652;
wire n_1286;
wire n_6021;
wire n_11880;
wire n_19531;
wire n_4617;
wire n_20031;
wire n_3169;
wire n_18013;
wire n_18051;
wire n_12136;
wire n_6511;
wire n_2203;
wire n_18376;
wire n_1426;
wire n_17531;
wire n_17618;
wire n_11089;
wire n_17524;
wire n_11608;
wire n_13756;
wire n_4641;
wire n_15564;
wire n_20620;
wire n_12364;
wire n_19672;
wire n_7728;
wire n_17517;
wire n_19729;
wire n_7359;
wire n_10489;
wire n_253;
wire n_10347;
wire n_9937;
wire n_18929;
wire n_13168;
wire n_20840;
wire n_20200;
wire n_17774;
wire n_16170;
wire n_10952;
wire n_17022;
wire n_17700;
wire n_10758;
wire n_15798;
wire n_9453;
wire n_16128;
wire n_18603;
wire n_4769;
wire n_14164;
wire n_18842;
wire n_12358;
wire n_1958;
wire n_9178;
wire n_9689;
wire n_13999;
wire n_18884;
wire n_1422;
wire n_644;
wire n_5167;
wire n_18657;
wire n_12851;
wire n_12307;
wire n_5104;
wire n_16236;
wire n_13807;
wire n_17260;
wire n_511;
wire n_20577;
wire n_13395;
wire n_19186;
wire n_7720;
wire n_18609;
wire n_18702;
wire n_16152;
wire n_10404;
wire n_19836;
wire n_1049;
wire n_19690;
wire n_141;
wire n_19911;
wire n_5338;
wire n_7440;
wire n_9568;
wire n_1773;
wire n_18556;
wire n_5578;
wire n_12654;
wire n_19682;
wire n_12921;
wire n_2401;
wire n_19445;
wire n_16140;
wire n_3255;
wire n_2588;
wire n_935;
wire n_4961;
wire n_10221;
wire n_17120;
wire n_3770;
wire n_11465;
wire n_16935;
wire n_13221;
wire n_628;
wire n_5863;
wire n_18229;
wire n_7118;
wire n_9234;
wire n_9431;
wire n_10023;
wire n_8281;
wire n_12347;
wire n_12958;
wire n_3662;
wire n_6169;
wire n_7069;
wire n_5199;
wire n_13347;
wire n_17468;
wire n_4282;
wire n_10673;
wire n_10467;
wire n_8766;
wire n_13976;
wire n_16823;
wire n_4027;
wire n_4309;
wire n_20624;
wire n_609;
wire n_16350;
wire n_4944;
wire n_19333;
wire n_18960;
wire n_9380;
wire n_7666;
wire n_12353;
wire n_1774;
wire n_10818;
wire n_9976;
wire n_17697;
wire n_16474;
wire n_5977;
wire n_19735;
wire n_15311;
wire n_8239;
wire n_3583;
wire n_11905;
wire n_9746;
wire n_3540;
wire n_4930;
wire n_234;
wire n_13856;
wire n_5945;
wire n_4423;
wire n_10519;
wire n_18345;
wire n_3689;
wire n_7584;
wire n_16409;
wire n_6301;
wire n_15988;
wire n_2315;
wire n_14982;
wire n_21031;
wire n_14648;
wire n_15349;
wire n_15725;
wire n_6985;
wire n_10723;
wire n_17813;
wire n_2444;
wire n_9455;
wire n_2977;
wire n_10653;
wire n_6384;
wire n_15345;
wire n_15571;
wire n_15777;
wire n_585;
wire n_9916;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_12402;
wire n_14387;
wire n_19259;
wire n_5869;
wire n_9690;
wire n_11594;
wire n_9002;
wire n_10619;
wire n_14535;
wire n_13403;
wire n_11655;
wire n_3664;
wire n_19726;
wire n_434;
wire n_14060;
wire n_10871;
wire n_18012;
wire n_8518;
wire n_4720;
wire n_12670;
wire n_14923;
wire n_8350;
wire n_243;
wire n_11833;
wire n_17055;
wire n_5221;
wire n_8148;
wire n_1407;
wire n_8408;
wire n_6145;
wire n_8236;
wire n_14202;
wire n_16421;
wire n_14352;
wire n_9587;
wire n_1176;
wire n_13888;
wire n_15370;
wire n_13529;
wire n_12452;
wire n_13530;
wire n_3989;
wire n_4752;
wire n_5449;
wire n_8760;
wire n_15032;
wire n_17161;
wire n_16246;
wire n_4158;
wire n_10466;
wire n_6812;
wire n_3079;
wire n_558;
wire n_4231;
wire n_2591;
wire n_653;
wire n_6262;
wire n_2050;
wire n_4872;
wire n_10461;
wire n_15827;
wire n_18599;
wire n_170;
wire n_12721;
wire n_10113;
wire n_1471;
wire n_13023;
wire n_16150;
wire n_9194;
wire n_13268;
wire n_2816;
wire n_20432;
wire n_16809;
wire n_7678;
wire n_4837;
wire n_14848;
wire n_11248;
wire n_13660;
wire n_15712;
wire n_17053;
wire n_2169;
wire n_6953;
wire n_9652;
wire n_13143;
wire n_21125;
wire n_12966;
wire n_5305;
wire n_2175;
wire n_5689;
wire n_7891;
wire n_17494;
wire n_16904;
wire n_9137;
wire n_9390;
wire n_20030;
wire n_11995;
wire n_8038;
wire n_8190;
wire n_11701;
wire n_15803;
wire n_9080;
wire n_17141;
wire n_15878;
wire n_940;
wire n_13544;
wire n_1537;
wire n_15060;
wire n_19578;
wire n_20923;
wire n_17833;
wire n_17472;
wire n_7994;
wire n_9883;
wire n_8287;
wire n_18496;
wire n_13527;
wire n_13206;
wire n_13235;
wire n_4998;
wire n_13399;
wire n_20604;
wire n_18811;
wire n_19352;
wire n_7345;
wire n_1530;
wire n_13622;
wire n_5918;
wire n_631;
wire n_17598;
wire n_2724;
wire n_18442;
wire n_8965;
wire n_16635;
wire n_2258;
wire n_13564;
wire n_17085;
wire n_2012;
wire n_9600;
wire n_3182;
wire n_17460;
wire n_6871;
wire n_6672;
wire n_4021;
wire n_7028;
wire n_16373;
wire n_10645;
wire n_16544;
wire n_16505;
wire n_20506;
wire n_5835;
wire n_8579;
wire n_18289;
wire n_2948;
wire n_13792;
wire n_16319;
wire n_4812;
wire n_8973;
wire n_18140;
wire n_2583;
wire n_13764;
wire n_19441;
wire n_19204;
wire n_3155;
wire n_11264;
wire n_16018;
wire n_1770;
wire n_4472;
wire n_12516;
wire n_9819;
wire n_20362;
wire n_15722;
wire n_2699;
wire n_13698;
wire n_5819;
wire n_14959;
wire n_8612;
wire n_19898;
wire n_16978;
wire n_19615;
wire n_9292;
wire n_20513;
wire n_17513;
wire n_15977;
wire n_9018;
wire n_18417;
wire n_13741;
wire n_20065;
wire n_17429;
wire n_20293;
wire n_19021;
wire n_4197;
wire n_13440;
wire n_20989;
wire n_11495;
wire n_13325;
wire n_2721;
wire n_2615;
wire n_4787;
wire n_8218;
wire n_14006;
wire n_3933;
wire n_14757;
wire n_188;
wire n_16422;
wire n_5828;
wire n_7210;
wire n_16426;
wire n_15619;
wire n_14107;
wire n_7733;
wire n_13496;
wire n_921;
wire n_2104;
wire n_16678;
wire n_11293;
wire n_15122;
wire n_15341;
wire n_18519;
wire n_16805;
wire n_20625;
wire n_10700;
wire n_11961;
wire n_8306;
wire n_2088;
wire n_11981;
wire n_4238;
wire n_15391;
wire n_12172;
wire n_17447;
wire n_18571;
wire n_14897;
wire n_14476;
wire n_8342;
wire n_10502;
wire n_18137;
wire n_11239;
wire n_14221;
wire n_20742;
wire n_17544;
wire n_4189;
wire n_2705;
wire n_16254;
wire n_1316;
wire n_6264;
wire n_17659;
wire n_9264;
wire n_4168;
wire n_8582;
wire n_20612;
wire n_13181;
wire n_13004;
wire n_11067;
wire n_3143;
wire n_8044;
wire n_19844;
wire n_3229;
wire n_5864;
wire n_8921;
wire n_14072;
wire n_13397;
wire n_19903;
wire n_235;
wire n_10010;
wire n_12984;
wire n_2504;
wire n_17170;
wire n_16109;
wire n_9646;
wire n_18775;
wire n_18658;
wire n_8405;
wire n_13296;
wire n_13816;
wire n_6990;
wire n_2451;
wire n_17379;
wire n_2913;
wire n_13989;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_11228;
wire n_16583;
wire n_19860;
wire n_12725;
wire n_4036;
wire n_9671;
wire n_8430;
wire n_4807;
wire n_8426;
wire n_12474;
wire n_15056;
wire n_1723;
wire n_5324;
wire n_17233;
wire n_4830;
wire n_4391;
wire n_12484;
wire n_17371;
wire n_18945;
wire n_4095;
wire n_8507;
wire n_9188;
wire n_18080;
wire n_3327;
wire n_9231;
wire n_18102;
wire n_18999;
wire n_17673;
wire n_19776;
wire n_6679;
wire n_12862;
wire n_13442;
wire n_17008;
wire n_10201;
wire n_16144;
wire n_15128;
wire n_20485;
wire n_16008;
wire n_19554;
wire n_4573;
wire n_4943;
wire n_10676;
wire n_6599;
wire n_16609;
wire n_4042;
wire n_20660;
wire n_16554;
wire n_17122;
wire n_4708;
wire n_7052;
wire n_8428;
wire n_17671;
wire n_17199;
wire n_1634;
wire n_17057;
wire n_1203;
wire n_14634;
wire n_18989;
wire n_937;
wire n_11615;
wire n_11079;
wire n_14772;
wire n_9180;
wire n_9017;
wire n_9269;
wire n_5696;
wire n_19393;
wire n_20394;
wire n_20517;
wire n_16123;
wire n_2891;
wire n_16215;
wire n_13656;
wire n_11668;
wire n_13641;
wire n_12487;
wire n_7394;
wire n_9502;
wire n_4516;
wire n_18174;
wire n_7627;
wire n_6436;
wire n_9316;
wire n_18419;
wire n_14479;
wire n_14410;
wire n_7462;
wire n_18527;
wire n_19150;
wire n_6027;
wire n_13321;
wire n_10911;
wire n_11547;
wire n_11064;
wire n_9873;
wire n_1228;
wire n_10473;
wire n_15120;
wire n_19510;
wire n_7555;
wire n_12552;
wire n_6110;
wire n_14123;
wire n_17642;
wire n_12777;
wire n_19216;
wire n_9978;
wire n_16367;
wire n_15235;
wire n_5331;
wire n_10672;
wire n_9494;
wire n_4134;
wire n_5018;
wire n_19331;
wire n_19871;
wire n_4017;
wire n_12437;
wire n_1730;
wire n_13739;
wire n_2752;
wire n_3527;
wire n_4030;
wire n_19059;
wire n_11913;
wire n_20476;
wire n_17332;
wire n_3056;
wire n_18939;
wire n_2679;
wire n_16227;
wire n_6581;
wire n_5553;
wire n_7277;
wire n_16580;
wire n_19287;
wire n_17013;
wire n_4283;
wire n_11627;
wire n_8139;
wire n_4962;
wire n_19282;
wire n_11306;
wire n_15390;
wire n_17909;
wire n_15157;
wire n_17277;
wire n_13109;
wire n_14209;
wire n_5090;
wire n_864;
wire n_5302;
wire n_1379;
wire n_19738;
wire n_19125;
wire n_5712;
wire n_10704;
wire n_11431;
wire n_462;
wire n_9734;
wire n_2646;
wire n_8257;
wire n_737;
wire n_10213;
wire n_232;
wire n_4028;
wire n_5565;
wire n_6358;
wire n_8546;
wire n_2482;
wire n_15841;
wire n_17606;
wire n_17550;
wire n_958;
wire n_2554;
wire n_14473;
wire n_4321;
wire n_15801;
wire n_10468;
wire n_9241;
wire n_16032;
wire n_16284;
wire n_19992;
wire n_8744;
wire n_12574;
wire n_6313;
wire n_9939;
wire n_239;
wire n_19537;
wire n_6664;
wire n_11604;
wire n_9997;
wire n_7534;
wire n_17808;
wire n_17966;
wire n_6190;
wire n_1364;
wire n_7373;
wire n_10281;
wire n_16224;
wire n_2322;
wire n_331;
wire n_495;
wire n_4824;
wire n_12728;
wire n_7467;
wire n_20385;
wire n_350;
wire n_16657;
wire n_381;
wire n_18494;
wire n_14405;
wire n_14598;
wire n_10399;
wire n_8664;
wire n_18515;
wire n_17610;
wire n_901;
wire n_13058;
wire n_18151;
wire n_4136;
wire n_18311;
wire n_20495;
wire n_9295;
wire n_15363;
wire n_15602;
wire n_10595;
wire n_13180;
wire n_15577;
wire n_6253;
wire n_17000;
wire n_2950;
wire n_7200;
wire n_8326;
wire n_13090;
wire n_2847;
wire n_11819;
wire n_8920;
wire n_6808;
wire n_3749;
wire n_16257;
wire n_8985;
wire n_20181;
wire n_12599;
wire n_20096;
wire n_3960;
wire n_3975;
wire n_8035;
wire n_16652;
wire n_15063;
wire n_2004;
wire n_4018;
wire n_8660;
wire n_192;
wire n_15593;
wire n_9917;
wire n_5152;
wire n_20944;
wire n_16701;
wire n_20388;
wire n_13896;
wire n_20795;
wire n_16277;
wire n_16705;
wire n_20062;
wire n_273;
wire n_11974;
wire n_6452;
wire n_10426;
wire n_5247;
wire n_9512;
wire n_9923;
wire n_8469;
wire n_7306;
wire n_16368;
wire n_20223;
wire n_7507;
wire n_1267;
wire n_19972;
wire n_5210;
wire n_7379;
wire n_1213;
wire n_12556;
wire n_11200;
wire n_4443;
wire n_6136;
wire n_3458;
wire n_17912;
wire n_17811;
wire n_14587;
wire n_20125;
wire n_19296;
wire n_13830;
wire n_15665;
wire n_490;
wire n_575;
wire n_10245;
wire n_6156;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_12509;
wire n_4432;
wire n_10457;
wire n_11682;
wire n_19200;
wire n_9821;
wire n_2245;
wire n_16187;
wire n_5452;
wire n_14762;
wire n_12068;
wire n_20138;
wire n_3539;
wire n_5757;
wire n_19006;
wire n_6644;
wire n_2134;
wire n_18209;
wire n_20478;
wire n_12140;
wire n_9845;
wire n_3284;
wire n_17227;
wire n_13330;
wire n_7642;
wire n_14492;
wire n_1386;
wire n_7104;
wire n_15909;
wire n_4827;
wire n_6801;
wire n_1661;
wire n_16321;
wire n_4405;
wire n_15420;
wire n_10781;
wire n_13243;
wire n_3029;
wire n_2398;
wire n_5971;
wire n_19171;
wire n_18639;
wire n_16346;
wire n_13063;
wire n_15748;
wire n_7259;
wire n_12961;
wire n_20733;
wire n_11398;
wire n_12389;
wire n_2877;
wire n_4951;
wire n_12595;
wire n_11858;
wire n_14194;
wire n_13237;
wire n_619;
wire n_14255;
wire n_10239;
wire n_20653;
wire n_1357;
wire n_8560;
wire n_15360;
wire n_18039;
wire n_17674;
wire n_14990;
wire n_10464;
wire n_14166;
wire n_9715;
wire n_4905;
wire n_9016;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_6659;
wire n_9399;
wire n_7351;
wire n_959;
wire n_20701;
wire n_1101;
wire n_14353;
wire n_12020;
wire n_19748;
wire n_13272;
wire n_3372;
wire n_3559;
wire n_5778;
wire n_18460;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_16431;
wire n_10776;
wire n_14914;
wire n_13536;
wire n_632;
wire n_20423;
wire n_17624;
wire n_15212;
wire n_19255;
wire n_14093;
wire n_3493;
wire n_20442;
wire n_19782;
wire n_16101;
wire n_3700;
wire n_12706;
wire n_2795;
wire n_1680;
wire n_15825;
wire n_18162;
wire n_16807;
wire n_11031;
wire n_14929;
wire n_6538;
wire n_13815;
wire n_9648;
wire n_12470;
wire n_7717;
wire n_18385;
wire n_5091;
wire n_15483;
wire n_17313;
wire n_8675;
wire n_17817;
wire n_9095;
wire n_2019;
wire n_698;
wire n_9048;
wire n_1992;
wire n_10578;
wire n_646;
wire n_12093;
wire n_15247;
wire n_9932;
wire n_3438;
wire n_8220;
wire n_19344;
wire n_15170;
wire n_17327;
wire n_2625;
wire n_11779;
wire n_12724;
wire n_14557;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_18189;
wire n_3147;
wire n_3661;
wire n_18625;
wire n_4179;
wire n_20996;
wire n_11609;
wire n_16793;
wire n_133;
wire n_1029;
wire n_6860;
wire n_522;
wire n_1568;
wire n_7322;
wire n_5788;
wire n_12566;
wire n_20153;
wire n_19837;
wire n_5951;
wire n_5647;
wire n_18084;
wire n_12035;
wire n_2631;
wire n_12212;
wire n_9110;
wire n_3516;
wire n_4442;
wire n_424;
wire n_9969;
wire n_11375;
wire n_15749;
wire n_18003;
wire n_3087;
wire n_17641;
wire n_15004;
wire n_8243;
wire n_8798;
wire n_18128;
wire n_13893;
wire n_14699;
wire n_10683;
wire n_14232;
wire n_17132;
wire n_6615;
wire n_20595;
wire n_6192;
wire n_5773;
wire n_16907;
wire n_1032;
wire n_1592;
wire n_20812;
wire n_4714;
wire n_3074;
wire n_11878;
wire n_17405;
wire n_16738;
wire n_6418;
wire n_9437;
wire n_4588;
wire n_5149;
wire n_5280;
wire n_20870;
wire n_16046;
wire n_19227;
wire n_5052;
wire n_5137;
wire n_7141;
wire n_14116;
wire n_5775;
wire n_8961;
wire n_14551;
wire n_18662;
wire n_3323;
wire n_14940;
wire n_4643;
wire n_10826;
wire n_15086;
wire n_13886;
wire n_2476;
wire n_11973;
wire n_7416;
wire n_5031;
wire n_1665;
wire n_9669;
wire n_5082;
wire n_4788;
wire n_10835;
wire n_1414;
wire n_4555;
wire n_1901;
wire n_10416;
wire n_7191;
wire n_5796;
wire n_14411;
wire n_1906;
wire n_6761;
wire n_14304;
wire n_10860;
wire n_19461;
wire n_16672;
wire n_4780;
wire n_20523;
wire n_17752;
wire n_19660;
wire n_15162;
wire n_19464;
wire n_13889;
wire n_5985;
wire n_604;
wire n_1061;
wire n_4157;
wire n_10124;
wire n_20673;
wire n_874;
wire n_7654;
wire n_16604;
wire n_5336;
wire n_18629;
wire n_18789;
wire n_16742;
wire n_11321;
wire n_4292;
wire n_688;
wire n_14233;
wire n_8334;
wire n_1490;
wire n_1553;
wire n_1086;
wire n_15912;
wire n_8513;
wire n_887;
wire n_20809;
wire n_10948;
wire n_14056;
wire n_10927;
wire n_11496;
wire n_1156;
wire n_14151;
wire n_13727;
wire n_2861;
wire n_3130;
wire n_21030;
wire n_4216;
wire n_18402;
wire n_15002;
wire n_18933;
wire n_6482;
wire n_15585;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_15329;
wire n_14619;
wire n_4864;
wire n_19115;
wire n_2226;
wire n_5742;
wire n_10731;
wire n_15169;
wire n_5255;
wire n_15565;
wire n_13198;
wire n_5933;
wire n_9874;
wire n_4946;
wire n_4848;
wire n_4941;
wire n_21005;
wire n_1189;
wire n_14832;
wire n_14691;
wire n_9082;
wire n_16612;
wire n_17827;
wire n_11500;
wire n_20674;
wire n_9596;
wire n_16986;
wire n_11109;
wire n_12909;
wire n_10729;
wire n_10973;
wire n_4182;
wire n_12822;
wire n_3214;
wire n_14948;
wire n_3373;
wire n_5539;
wire n_12267;
wire n_1844;
wire n_15876;
wire n_1953;
wire n_20585;
wire n_17336;
wire n_19656;
wire n_17897;
wire n_13469;
wire n_16970;
wire n_4729;
wire n_16260;
wire n_14229;
wire n_14425;
wire n_4800;
wire n_15324;
wire n_13076;
wire n_14917;
wire n_5427;
wire n_6508;
wire n_16598;
wire n_7989;
wire n_13082;
wire n_8047;
wire n_15064;
wire n_3696;
wire n_9233;
wire n_19691;
wire n_10529;
wire n_16863;
wire n_20878;
wire n_20012;
wire n_1529;
wire n_8751;
wire n_20319;
wire n_18022;
wire n_14444;
wire n_1007;
wire n_9435;
wire n_18119;
wire n_4925;
wire n_7254;
wire n_951;
wire n_13677;
wire n_18520;
wire n_14422;
wire n_11997;
wire n_6628;
wire n_10270;
wire n_8684;
wire n_4765;
wire n_9721;
wire n_4863;
wire n_18585;
wire n_12363;
wire n_13115;
wire n_15599;
wire n_1766;
wire n_1338;
wire n_16499;
wire n_12008;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_14498;
wire n_10689;
wire n_9507;
wire n_5476;
wire n_18820;
wire n_19620;
wire n_19494;
wire n_8090;
wire n_7605;
wire n_15513;
wire n_15330;
wire n_12748;
wire n_12272;
wire n_20710;
wire n_10363;
wire n_6124;
wire n_317;
wire n_3197;
wire n_19435;
wire n_13388;
wire n_14484;
wire n_7423;
wire n_13674;
wire n_16308;
wire n_6344;
wire n_8811;
wire n_14486;
wire n_14580;
wire n_18522;
wire n_14421;
wire n_4694;
wire n_4664;
wire n_14703;
wire n_14653;
wire n_8573;
wire n_4633;
wire n_2026;
wire n_20845;
wire n_642;
wire n_5073;
wire n_6360;
wire n_19113;
wire n_2684;
wire n_17931;
wire n_17557;
wire n_13377;
wire n_11455;
wire n_17257;
wire n_3452;
wire n_474;
wire n_17479;
wire n_21033;
wire n_18578;
wire n_18083;
wire n_5894;
wire n_13750;
wire n_12639;
wire n_8339;
wire n_1596;
wire n_2723;
wire n_2016;
wire n_19480;
wire n_12428;
wire n_14384;
wire n_4689;
wire n_5165;
wire n_6102;
wire n_1874;
wire n_16948;
wire n_14276;
wire n_3780;
wire n_1657;
wire n_13488;
wire n_6650;
wire n_10024;
wire n_12214;
wire n_3753;
wire n_6244;
wire n_9250;
wire n_10191;
wire n_20471;
wire n_4076;
wire n_7148;
wire n_7169;
wire n_15297;
wire n_9350;
wire n_11257;
wire n_12330;
wire n_9441;
wire n_7600;
wire n_9124;
wire n_18684;
wire n_20243;
wire n_14645;
wire n_12926;
wire n_18510;
wire n_1829;
wire n_13094;
wire n_6804;
wire n_1493;
wire n_2911;
wire n_515;
wire n_6427;
wire n_17100;
wire n_14459;
wire n_4281;
wire n_14811;
wire n_16696;
wire n_4419;
wire n_17063;
wire n_5405;
wire n_9750;
wire n_18834;
wire n_7660;
wire n_13735;
wire n_9529;
wire n_20409;
wire n_10339;
wire n_16357;
wire n_17448;
wire n_10606;
wire n_3421;
wire n_1448;
wire n_19086;
wire n_10054;
wire n_8261;
wire n_6645;
wire n_15020;
wire n_13985;
wire n_6749;
wire n_19034;
wire n_13342;
wire n_2612;
wire n_20375;
wire n_8702;
wire n_11601;
wire n_14250;
wire n_10944;
wire n_6247;
wire n_5921;
wire n_1849;
wire n_11710;
wire n_2250;
wire n_9940;
wire n_20853;
wire n_12476;
wire n_4188;
wire n_21060;
wire n_2001;
wire n_15273;
wire n_11010;
wire n_15901;
wire n_4825;
wire n_3715;
wire n_20497;
wire n_9443;
wire n_17092;
wire n_8429;
wire n_10419;
wire n_15726;
wire n_15470;
wire n_8486;
wire n_18550;
wire n_2070;
wire n_13123;
wire n_7431;
wire n_398;
wire n_17214;
wire n_3842;
wire n_17759;
wire n_166;
wire n_8117;
wire n_18035;
wire n_17239;
wire n_825;
wire n_2619;
wire n_19528;
wire n_10058;
wire n_10355;
wire n_7253;
wire n_5208;
wire n_17215;
wire n_5113;
wire n_10304;
wire n_19079;
wire n_11955;
wire n_12538;
wire n_12151;
wire n_1160;
wire n_1976;
wire n_2711;
wire n_12409;
wire n_3386;
wire n_400;
wire n_15411;
wire n_10060;
wire n_16600;
wire n_20843;
wire n_1517;
wire n_2647;
wire n_16891;
wire n_3380;
wire n_2826;
wire n_5825;
wire n_846;
wire n_1398;
wire n_1921;
wire n_14886;
wire n_17319;
wire n_5629;
wire n_13167;
wire n_1504;
wire n_9590;
wire n_7498;
wire n_11829;
wire n_20321;
wire n_12680;
wire n_11581;
wire n_19339;
wire n_7453;
wire n_16184;
wire n_12163;
wire n_19821;
wire n_3818;
wire n_14131;
wire n_18547;
wire n_7932;
wire n_5599;
wire n_3587;
wire n_19236;
wire n_6004;
wire n_9763;
wire n_21108;
wire n_810;
wire n_4278;
wire n_12738;
wire n_1959;
wire n_6275;
wire n_3497;
wire n_14622;
wire n_4542;
wire n_9966;
wire n_6350;
wire n_16115;
wire n_565;
wire n_7189;
wire n_19880;
wire n_4060;
wire n_9341;
wire n_14984;
wire n_20150;
wire n_5807;
wire n_18819;
wire n_6475;
wire n_12525;
wire n_11132;
wire n_12932;
wire n_14849;
wire n_19010;
wire n_17267;
wire n_16064;
wire n_16407;
wire n_1521;
wire n_12037;
wire n_15147;
wire n_10030;
wire n_16288;
wire n_20373;
wire n_4722;
wire n_16929;
wire n_16726;
wire n_18749;
wire n_8163;
wire n_11947;
wire n_16914;
wire n_4126;
wire n_20208;
wire n_2561;
wire n_1056;
wire n_12424;
wire n_5320;
wire n_12942;
wire n_9038;
wire n_17703;
wire n_8698;
wire n_10709;
wire n_3911;
wire n_1584;
wire n_11436;
wire n_11909;
wire n_9034;
wire n_4922;
wire n_6066;
wire n_629;
wire n_13150;
wire n_12747;
wire n_20507;
wire n_14564;
wire n_216;
wire n_6638;
wire n_7063;
wire n_4509;
wire n_8384;
wire n_834;
wire n_3630;
wire n_14044;
wire n_16415;
wire n_5906;
wire n_2189;
wire n_14431;
wire n_20016;
wire n_16908;
wire n_16258;
wire n_20276;
wire n_10478;
wire n_10534;
wire n_8374;
wire n_16702;
wire n_6474;
wire n_13662;
wire n_16677;
wire n_4111;
wire n_7510;
wire n_9041;
wire n_875;
wire n_1626;
wire n_19358;
wire n_14240;
wire n_1715;
wire n_9011;
wire n_4204;
wire n_20440;
wire n_3553;
wire n_5323;
wire n_6744;
wire n_15055;
wire n_12660;
wire n_14708;
wire n_10695;
wire n_21103;
wire n_1485;
wire n_2883;
wire n_15823;
wire n_7735;
wire n_8531;
wire n_8074;
wire n_14246;
wire n_7495;
wire n_17567;
wire n_2870;
wire n_16143;
wire n_13857;
wire n_19757;
wire n_9288;
wire n_5011;
wire n_18744;
wire n_1554;
wire n_15047;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_13696;
wire n_10043;
wire n_4832;
wire n_2010;
wire n_13041;
wire n_1952;
wire n_5784;
wire n_15806;
wire n_5128;
wire n_13498;
wire n_14290;
wire n_2356;
wire n_12403;
wire n_17840;
wire n_15099;
wire n_10440;
wire n_15618;
wire n_18610;
wire n_13000;
wire n_4053;
wire n_18918;
wire n_11980;
wire n_7620;
wire n_20470;
wire n_12837;
wire n_3091;
wire n_13937;
wire n_16442;
wire n_1024;
wire n_176;
wire n_12764;
wire n_17271;
wire n_2518;
wire n_14687;
wire n_13508;
wire n_10706;
wire n_4596;
wire n_18007;
wire n_13224;
wire n_17354;
wire n_908;
wire n_19030;
wire n_1036;
wire n_14993;
wire n_15608;
wire n_20007;
wire n_10297;
wire n_19973;
wire n_11296;
wire n_10605;
wire n_9446;
wire n_16234;
wire n_3680;
wire n_3565;
wire n_7885;
wire n_14100;
wire n_15410;
wire n_6905;
wire n_17437;
wire n_9865;
wire n_8456;
wire n_7722;
wire n_5824;
wire n_19773;
wire n_2453;
wire n_3331;
wire n_13179;
wire n_10458;
wire n_12947;
wire n_2138;
wire n_4230;
wire n_19440;
wire n_11892;
wire n_7817;
wire n_6413;
wire n_1809;
wire n_11105;
wire n_8293;
wire n_7299;
wire n_917;
wire n_18350;
wire n_8029;
wire n_18109;
wire n_20888;
wire n_3847;
wire n_6960;
wire n_1261;
wire n_7249;
wire n_16715;
wire n_15062;
wire n_363;
wire n_6061;
wire n_17385;
wire n_9769;
wire n_1462;
wire n_7002;
wire n_1446;
wire n_15688;
wire n_19551;
wire n_19369;
wire n_1701;
wire n_7396;
wire n_19384;
wire n_731;
wire n_20315;
wire n_2997;
wire n_16783;
wire n_18178;
wire n_6746;
wire n_6545;
wire n_6763;
wire n_13415;
wire n_1106;
wire n_2009;
wire n_1473;
wire n_5895;
wire n_753;
wire n_4024;
wire n_19303;
wire n_17797;
wire n_485;
wire n_4064;
wire n_3351;
wire n_16703;
wire n_14767;
wire n_19179;
wire n_17636;
wire n_2324;
wire n_17337;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_14794;
wire n_8113;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_14446;
wire n_15877;
wire n_7140;
wire n_20033;
wire n_20963;
wire n_4066;
wire n_19122;
wire n_15091;
wire n_9228;
wire n_3303;
wire n_13461;
wire n_7910;
wire n_10214;
wire n_13979;
wire n_10354;
wire n_248;
wire n_12060;
wire n_7741;
wire n_18205;
wire n_4295;
wire n_11450;
wire n_11723;
wire n_18466;
wire n_1265;
wire n_14062;
wire n_8232;
wire n_12842;
wire n_1588;
wire n_12499;
wire n_21118;
wire n_21121;
wire n_3235;
wire n_18551;
wire n_3265;
wire n_18480;
wire n_12693;
wire n_20333;
wire n_19822;
wire n_7698;
wire n_14873;
wire n_16927;
wire n_18911;
wire n_10164;
wire n_3285;
wire n_10205;
wire n_1039;
wire n_5676;
wire n_12326;
wire n_6336;
wire n_1628;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_16276;
wire n_9818;
wire n_17291;
wire n_4777;
wire n_3941;
wire n_16563;
wire n_5399;
wire n_14004;
wire n_11698;
wire n_2846;
wire n_3371;
wire n_10338;
wire n_9599;
wire n_8674;
wire n_8016;
wire n_5760;
wire n_12483;
wire n_18802;
wire n_9935;
wire n_17107;
wire n_12258;
wire n_11871;
wire n_8966;
wire n_16291;
wire n_14826;
wire n_19833;
wire n_10018;
wire n_3366;
wire n_15537;
wire n_6998;
wire n_16537;
wire n_13209;
wire n_7650;
wire n_3020;
wire n_12823;
wire n_20649;
wire n_7535;
wire n_19084;
wire n_708;
wire n_17699;
wire n_17349;
wire n_12905;
wire n_10291;
wire n_17731;
wire n_2017;
wire n_1810;
wire n_12849;
wire n_11167;
wire n_11297;
wire n_9473;
wire n_10208;
wire n_3555;
wire n_19598;
wire n_11285;
wire n_11740;
wire n_15428;
wire n_19083;
wire n_14679;
wire n_6494;
wire n_17865;
wire n_8980;
wire n_11434;
wire n_16480;
wire n_8336;
wire n_21084;
wire n_13711;
wire n_774;
wire n_16261;
wire n_6974;
wire n_14783;
wire n_219;
wire n_18411;
wire n_3762;
wire n_6498;
wire n_6562;
wire n_12442;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_14649;
wire n_17131;
wire n_768;
wire n_3707;
wire n_10434;
wire n_5917;
wire n_15853;
wire n_12419;
wire n_16399;
wire n_2058;
wire n_3231;
wire n_14210;
wire n_13262;
wire n_6168;
wire n_20257;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_946;
wire n_9729;
wire n_3398;
wire n_13543;
wire n_19286;
wire n_20791;
wire n_2536;
wire n_10263;
wire n_18082;
wire n_8473;
wire n_8351;
wire n_7276;
wire n_174;
wire n_19653;
wire n_17552;
wire n_12410;
wire n_963;
wire n_7085;
wire n_12938;
wire n_4120;
wire n_13493;
wire n_1115;
wire n_12572;
wire n_10318;
wire n_3158;
wire n_11039;
wire n_10128;
wire n_8020;
wire n_7946;
wire n_10717;
wire n_1010;
wire n_19404;
wire n_4622;
wire n_803;
wire n_1871;
wire n_9520;
wire n_19787;
wire n_6471;
wire n_6949;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_14128;
wire n_11818;
wire n_4570;
wire n_10945;
wire n_7920;
wire n_7841;
wire n_18287;
wire n_12469;
wire n_15387;
wire n_18251;
wire n_7054;
wire n_19230;
wire n_11555;
wire n_13917;
wire n_16388;
wire n_10565;
wire n_7837;
wire n_359;
wire n_6788;
wire n_15730;
wire n_20966;
wire n_1451;
wire n_5528;
wire n_2163;
wire n_6896;
wire n_18582;
wire n_5358;
wire n_12248;
wire n_10020;
wire n_12713;
wire n_8897;
wire n_5493;
wire n_6285;
wire n_14149;
wire n_3578;
wire n_1109;
wire n_7430;
wire n_19905;
wire n_2011;
wire n_18970;
wire n_20958;
wire n_5901;
wire n_17309;
wire n_11923;
wire n_717;
wire n_952;
wire n_16310;
wire n_2446;
wire n_6582;
wire n_20516;
wire n_7724;
wire n_5360;
wire n_15160;
wire n_19816;
wire n_17410;
wire n_12292;
wire n_4363;
wire n_1839;
wire n_1138;
wire n_214;
wire n_18722;
wire n_2374;
wire n_6115;
wire n_1225;
wire n_9866;
wire n_13808;
wire n_11975;
wire n_17947;
wire n_7879;
wire n_8730;
wire n_6607;
wire n_12854;
wire n_870;
wire n_7117;
wire n_813;
wire n_10082;
wire n_12796;
wire n_10870;
wire n_11914;
wire n_995;
wire n_12028;
wire n_8315;
wire n_16531;
wire n_11175;
wire n_10411;
wire n_6849;
wire n_2844;
wire n_11753;
wire n_9407;
wire n_6719;
wire n_10423;
wire n_8019;
wire n_11791;
wire n_7875;
wire n_13665;
wire n_8962;
wire n_14533;
wire n_2317;
wire n_2838;
wire n_13242;
wire n_1736;
wire n_15269;
wire n_20449;
wire n_2200;
wire n_2781;
wire n_6191;
wire n_13121;
wire n_9477;
wire n_16274;
wire n_13734;
wire n_14591;
wire n_7238;
wire n_3657;
wire n_2634;
wire n_13047;
wire n_21054;
wire n_21069;
wire n_18701;
wire n_7804;
wire n_20198;
wire n_15780;
wire n_14904;
wire n_17986;
wire n_13475;
wire n_20584;
wire n_11794;
wire n_16478;
wire n_9828;
wire n_19679;
wire n_7248;
wire n_3830;
wire n_13336;
wire n_5466;
wire n_15015;
wire n_6552;
wire n_10665;
wire n_6094;
wire n_14482;
wire n_12113;
wire n_16380;
wire n_518;
wire n_14214;
wire n_13202;
wire n_8196;
wire n_3420;
wire n_8822;
wire n_14483;
wire n_5738;
wire n_8885;
wire n_17678;
wire n_11564;
wire n_4782;
wire n_1539;
wire n_3412;
wire n_2162;
wire n_5953;
wire n_15799;
wire n_16439;
wire n_13811;
wire n_17356;
wire n_19713;
wire n_8152;
wire n_12491;
wire n_17166;
wire n_18111;
wire n_5119;
wire n_19981;
wire n_21021;
wire n_1703;
wire n_12454;
wire n_12992;
wire n_20955;
wire n_3297;
wire n_11708;
wire n_15407;
wire n_10098;
wire n_19001;
wire n_6935;
wire n_1560;
wire n_6984;
wire n_12046;
wire n_17340;
wire n_8058;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_12749;
wire n_3728;
wire n_6596;
wire n_14630;
wire n_512;
wire n_15302;
wire n_18714;
wire n_14464;
wire n_15188;
wire n_18108;
wire n_1790;
wire n_19610;
wire n_17218;
wire n_2788;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_14281;
wire n_18801;
wire n_705;
wire n_17821;
wire n_17616;
wire n_7667;
wire n_8024;
wire n_4562;
wire n_3554;
wire n_15233;
wire n_2717;
wire n_18234;
wire n_2981;
wire n_13959;
wire n_9930;
wire n_2743;
wire n_17078;
wire n_2466;
wire n_6593;
wire n_8748;
wire n_14420;
wire n_20972;
wire n_5423;
wire n_17657;
wire n_1594;
wire n_8393;
wire n_11117;
wire n_14613;
wire n_3767;
wire n_20502;
wire n_6056;
wire n_5866;
wire n_3692;
wire n_11475;
wire n_21016;
wire n_8912;
wire n_10612;
wire n_15613;
wire n_19666;
wire n_15676;
wire n_1260;
wire n_19770;
wire n_19909;
wire n_11223;
wire n_16667;
wire n_8740;
wire n_3391;
wire n_10104;
wire n_18487;
wire n_4786;
wire n_20154;
wire n_7908;
wire n_20759;
wire n_4354;
wire n_6315;
wire n_16133;
wire n_19327;
wire n_2855;
wire n_19511;
wire n_7675;
wire n_16328;
wire n_18979;
wire n_12329;
wire n_17835;
wire n_11631;
wire n_7774;
wire n_12611;
wire n_13034;
wire n_13122;
wire n_3460;
wire n_5155;
wire n_14337;
wire n_19360;
wire n_2202;
wire n_17454;
wire n_16746;
wire n_19053;
wire n_3530;
wire n_10087;
wire n_5540;
wire n_11782;
wire n_7381;
wire n_7999;
wire n_931;
wire n_4992;
wire n_5130;
wire n_14392;
wire n_14973;
wire n_9112;
wire n_7873;
wire n_16401;
wire n_12861;
wire n_19191;
wire n_1880;
wire n_5684;
wire n_13708;
wire n_7228;
wire n_14987;
wire n_19322;
wire n_1855;
wire n_19555;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2167;
wire n_2293;
wire n_15908;
wire n_18184;
wire n_4984;
wire n_4410;
wire n_9804;
wire n_12450;
wire n_3730;
wire n_16640;
wire n_18309;
wire n_18386;
wire n_7084;
wire n_2598;
wire n_976;
wire n_6390;
wire n_2302;
wire n_10806;
wire n_2294;
wire n_12309;
wire n_13401;
wire n_13891;
wire n_8557;
wire n_9384;
wire n_15894;
wire n_21046;
wire n_3625;
wire n_397;
wire n_3760;
wire n_3515;
wire n_12023;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_16287;
wire n_9906;
wire n_15942;
wire n_3744;
wire n_5457;
wire n_4022;
wire n_7764;
wire n_17021;
wire n_4336;
wire n_8128;
wire n_12719;
wire n_8359;
wire n_2223;
wire n_18071;
wire n_6271;
wire n_6572;
wire n_10211;
wire n_3981;
wire n_13749;
wire n_2681;
wire n_13945;
wire n_14172;
wire n_16501;
wire n_15177;
wire n_8443;
wire n_19092;
wire n_19064;
wire n_3138;
wire n_10819;
wire n_2860;
wire n_466;
wire n_9373;
wire n_4201;
wire n_14374;
wire n_20574;
wire n_16019;
wire n_11279;
wire n_9770;
wire n_11514;
wire n_5287;
wire n_4719;
wire n_19499;
wire n_3994;
wire n_11606;
wire n_1217;
wire n_10103;
wire n_17348;
wire n_12839;
wire n_17609;
wire n_16963;
wire n_12925;
wire n_11658;
wire n_10710;
wire n_4275;
wire n_3774;
wire n_17208;
wire n_15821;
wire n_17914;
wire n_9544;
wire n_2296;
wire n_14728;
wire n_15009;
wire n_11369;
wire n_19786;
wire n_14865;
wire n_11720;
wire n_18813;
wire n_20145;
wire n_4658;
wire n_13500;
wire n_14815;
wire n_7135;
wire n_8488;
wire n_1501;
wire n_17599;
wire n_11284;
wire n_19888;
wire n_20779;
wire n_12553;
wire n_7211;
wire n_5139;
wire n_20263;
wire n_7132;
wire n_12496;
wire n_18175;
wire n_16042;
wire n_7533;
wire n_13655;
wire n_6420;
wire n_16638;
wire n_3961;
wire n_7766;
wire n_11221;
wire n_1287;
wire n_11095;
wire n_16353;
wire n_11211;
wire n_7129;
wire n_4870;
wire n_6981;
wire n_4818;
wire n_12230;
wire n_8767;
wire n_15925;
wire n_14588;
wire n_6696;
wire n_8472;
wire n_21120;
wire n_6045;
wire n_14261;
wire n_15581;
wire n_17171;
wire n_6300;
wire n_18669;
wire n_13969;
wire n_10033;
wire n_6900;
wire n_15137;
wire n_6660;
wire n_5988;
wire n_17459;
wire n_17945;
wire n_10696;
wire n_3734;
wire n_9245;
wire n_15142;
wire n_5832;
wire n_15418;
wire n_13269;
wire n_7460;
wire n_7142;
wire n_16866;
wire n_6526;
wire n_16794;
wire n_2523;
wire n_1945;
wire n_11423;
wire n_12691;
wire n_3819;
wire n_16378;
wire n_4616;
wire n_5016;
wire n_9330;
wire n_14231;
wire n_8917;
wire n_12587;
wire n_17508;
wire n_14663;
wire n_3868;
wire n_11667;
wire n_18994;
wire n_8230;
wire n_10414;
wire n_6222;
wire n_19263;
wire n_12422;
wire n_9918;
wire n_390;
wire n_20115;
wire n_13853;
wire n_8465;
wire n_19901;
wire n_15421;
wire n_14701;
wire n_17723;
wire n_11633;
wire n_15697;
wire n_4826;
wire n_6453;
wire n_11142;
wire n_1395;
wire n_3892;
wire n_13773;
wire n_15582;
wire n_21039;
wire n_1346;
wire n_12196;
wire n_1089;
wire n_1478;
wire n_2555;
wire n_12493;
wire n_2708;
wire n_6597;
wire n_12440;
wire n_13800;
wire n_4049;
wire n_845;
wire n_19423;
wire n_20525;
wire n_17927;
wire n_16002;
wire n_5037;
wire n_7305;
wire n_17841;
wire n_5581;
wire n_14896;
wire n_8866;
wire n_13329;
wire n_11661;
wire n_3766;
wire n_9376;
wire n_12515;
wire n_17937;
wire n_16135;
wire n_278;
wire n_2266;
wire n_12249;
wire n_4324;
wire n_15298;
wire n_1907;
wire n_14462;
wire n_16574;
wire n_19783;
wire n_1719;
wire n_13051;
wire n_15206;
wire n_19450;
wire n_1372;
wire n_14514;
wire n_13812;
wire n_14733;
wire n_10762;
wire n_7353;
wire n_11935;
wire n_8054;
wire n_3791;
wire n_915;
wire n_11037;
wire n_8841;
wire n_14681;
wire n_14453;
wire n_19777;
wire n_6906;
wire n_18380;
wire n_19564;
wire n_15657;
wire n_15720;
wire n_3367;
wire n_4898;
wire n_21003;
wire n_2292;
wire n_2772;
wire n_14036;
wire n_20984;
wire n_19387;
wire n_14994;
wire n_10561;
wire n_16789;
wire n_7818;
wire n_7645;
wire n_18316;
wire n_17936;
wire n_3990;
wire n_11726;
wire n_14522;
wire n_15647;
wire n_1171;
wire n_10243;
wire n_5635;
wire n_8590;
wire n_17536;
wire n_14945;
wire n_7907;
wire n_16492;
wire n_8970;
wire n_17117;
wire n_2576;
wire n_8791;
wire n_5595;
wire n_521;
wire n_10165;
wire n_5380;
wire n_17842;
wire n_3735;
wire n_8703;
wire n_6422;
wire n_12147;
wire n_3069;
wire n_17734;
wire n_15755;
wire n_8864;
wire n_21109;
wire n_10985;
wire n_4891;
wire n_13791;
wire n_1257;
wire n_10587;
wire n_6611;
wire n_12102;
wire n_2137;
wire n_6019;
wire n_18085;
wire n_14611;
wire n_16100;
wire n_16760;
wire n_16878;
wire n_16508;
wire n_6976;
wire n_7234;
wire n_15860;
wire n_1449;
wire n_13538;
wire n_797;
wire n_9044;
wire n_14176;
wire n_5936;
wire n_20210;
wire n_17504;
wire n_5312;
wire n_20424;
wire n_16237;
wire n_8470;
wire n_15216;
wire n_2032;
wire n_19737;
wire n_8050;
wire n_3124;
wire n_20718;
wire n_14980;
wire n_9633;
wire n_2364;
wire n_15189;
wire n_2928;
wire n_13433;
wire n_14662;
wire n_1118;
wire n_2884;
wire n_3408;
wire n_11331;
wire n_19684;
wire n_11953;
wire n_4118;
wire n_3110;
wire n_9472;
wire n_16294;
wire n_3157;
wire n_12522;
wire n_13451;
wire n_20860;
wire n_1180;
wire n_1697;
wire n_5129;
wire n_649;
wire n_1561;
wire n_2405;
wire n_16102;
wire n_13191;
wire n_2700;
wire n_14133;
wire n_10690;
wire n_12681;
wire n_8143;
wire n_3640;
wire n_18604;
wire n_12084;
wire n_19864;
wire n_20581;
wire n_4744;
wire n_5626;
wire n_1505;
wire n_11861;
wire n_14443;
wire n_9101;
wire n_2454;
wire n_18856;
wire n_17241;
wire n_6550;
wire n_8574;
wire n_12832;
wire n_21114;
wire n_7043;
wire n_7986;
wire n_9927;
wire n_12782;
wire n_17489;
wire n_10621;
wire n_5653;
wire n_15507;
wire n_19867;
wire n_10789;
wire n_10496;
wire n_12384;
wire n_354;
wire n_18194;
wire n_4559;
wire n_15683;
wire n_14724;
wire n_15679;
wire n_15871;
wire n_10319;
wire n_16936;
wire n_14021;
wire n_1133;
wire n_883;
wire n_16223;
wire n_4372;
wire n_5396;
wire n_4162;
wire n_10499;
wire n_10224;
wire n_779;
wire n_4790;
wire n_7035;
wire n_20417;
wire n_19129;
wire n_15059;
wire n_6047;
wire n_9432;
wire n_3573;
wire n_2943;
wire n_11464;
wire n_3319;
wire n_11243;
wire n_17755;
wire n_10827;
wire n_16472;
wire n_3654;
wire n_5627;
wire n_18958;
wire n_19380;
wire n_10783;
wire n_2158;
wire n_8583;
wire n_7715;
wire n_19634;
wire n_11749;
wire n_7350;
wire n_16383;
wire n_13955;
wire n_20026;
wire n_9144;
wire n_18268;
wire n_12481;
wire n_4799;
wire n_16395;
wire n_5882;
wire n_12129;
wire n_5636;
wire n_9931;
wire n_7699;
wire n_16126;
wire n_15530;
wire n_465;
wire n_5707;
wire n_15474;
wire n_19614;
wire n_3738;
wire n_21091;
wire n_21008;
wire n_510;
wire n_12697;
wire n_17483;
wire n_19868;
wire n_13437;
wire n_11440;
wire n_15849;
wire n_12908;
wire n_7870;
wire n_7399;
wire n_5382;
wire n_11545;
wire n_13487;
wire n_15591;
wire n_13239;
wire n_18321;
wire n_3395;
wire n_9881;
wire n_11263;
wire n_19912;
wire n_13854;
wire n_13361;
wire n_20666;
wire n_8382;
wire n_20220;
wire n_11324;
wire n_18373;
wire n_13803;
wire n_19624;
wire n_2234;
wire n_20552;
wire n_17492;
wire n_14537;
wire n_3322;
wire n_10109;
wire n_20942;
wire n_10857;
wire n_15096;
wire n_715;
wire n_13244;
wire n_2331;
wire n_11359;
wire n_9630;
wire n_19486;
wire n_9898;
wire n_15926;
wire n_1712;
wire n_11620;
wire n_8340;
wire n_4754;
wire n_18859;
wire n_12850;
wire n_10179;
wire n_9636;
wire n_18296;
wire n_8369;
wire n_5043;
wire n_17383;
wire n_7339;
wire n_16581;
wire n_12898;
wire n_4241;
wire n_4183;
wire n_918;
wire n_19587;
wire n_2371;
wire n_19567;
wire n_19755;
wire n_13772;
wire n_19820;
wire n_6107;
wire n_12218;
wire n_10795;
wire n_13602;
wire n_6476;
wire n_16197;
wire n_2560;
wire n_4256;
wire n_20689;
wire n_1345;
wire n_3037;
wire n_1033;
wire n_7612;
wire n_14407;
wire n_15882;
wire n_15321;
wire n_20228;
wire n_11071;
wire n_15626;
wire n_11187;
wire n_12882;
wire n_3522;
wire n_17948;
wire n_8172;
wire n_18177;
wire n_13341;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_13400;
wire n_11271;
wire n_19940;
wire n_19310;
wire n_5101;
wire n_9738;
wire n_9252;
wire n_12800;
wire n_14259;
wire n_7594;
wire n_7321;
wire n_223;
wire n_1816;
wire n_2803;
wire n_10508;
wire n_3305;
wire n_15323;
wire n_13281;
wire n_7574;
wire n_2093;
wire n_14874;
wire n_7529;
wire n_3354;
wire n_20212;
wire n_19068;
wire n_6466;
wire n_11828;
wire n_19852;
wire n_14138;
wire n_4212;
wire n_622;
wire n_9779;
wire n_14244;
wire n_8930;
wire n_17901;
wire n_13114;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_12398;
wire n_4217;
wire n_14015;
wire n_12941;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_8364;
wire n_16306;
wire n_20784;
wire n_8981;
wire n_8490;
wire n_3873;
wire n_4649;
wire n_8785;
wire n_10210;
wire n_1204;
wire n_7843;
wire n_12998;
wire n_15952;
wire n_20433;
wire n_9047;
wire n_18909;
wire n_1360;
wire n_11641;
wire n_15464;
wire n_3076;
wire n_7261;
wire n_4592;
wire n_18482;
wire n_20382;
wire n_1564;
wire n_12038;
wire n_10533;
wire n_3701;
wire n_16585;
wire n_13978;
wire n_8100;
wire n_17784;
wire n_13563;
wire n_13141;
wire n_10993;
wire n_18324;
wire n_18528;
wire n_9320;
wire n_16777;
wire n_20515;
wire n_17884;
wire n_6767;
wire n_4656;
wire n_4862;
wire n_15001;
wire n_13517;
wire n_6755;
wire n_16602;
wire n_1721;
wire n_20785;
wire n_11062;
wire n_10940;
wire n_13783;
wire n_6780;
wire n_14038;
wire n_6635;
wire n_16899;
wire n_294;
wire n_14385;
wire n_19517;
wire n_14027;
wire n_7585;
wire n_17427;
wire n_1998;
wire n_13007;
wire n_16317;
wire n_12395;
wire n_7418;
wire n_2985;
wire n_21095;
wire n_2630;
wire n_6577;
wire n_13213;
wire n_10491;
wire n_17069;
wire n_17481;
wire n_2092;
wire n_13507;
wire n_3622;
wire n_8918;
wire n_11766;
wire n_1458;
wire n_12766;
wire n_18356;
wire n_13790;
wire n_19357;
wire n_19373;
wire n_13510;
wire n_1358;
wire n_8616;
wire n_6105;
wire n_826;
wire n_14346;
wire n_3520;
wire n_11960;
wire n_19091;
wire n_11274;
wire n_15699;
wire n_5923;
wire n_3687;
wire n_13806;
wire n_2676;
wire n_9831;
wire n_8436;
wire n_13261;
wire n_14717;
wire n_14167;
wire n_12137;
wire n_11624;
wire n_10580;
wire n_7921;
wire n_5193;
wire n_10512;
wire n_5514;
wire n_11917;
wire n_20572;
wire n_20875;
wire n_1282;
wire n_16745;
wire n_5143;
wire n_12434;
wire n_19026;
wire n_5049;
wire n_2212;
wire n_16403;
wire n_18191;
wire n_12881;
wire n_20166;
wire n_21094;
wire n_7863;
wire n_6493;
wire n_17763;
wire n_4019;
wire n_7968;
wire n_18986;
wire n_10507;
wire n_6023;
wire n_816;
wire n_1322;
wire n_19556;
wire n_7750;
wire n_20831;
wire n_16247;
wire n_12995;
wire n_10967;
wire n_1125;
wire n_14339;
wire n_14971;
wire n_16996;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_14180;
wire n_18846;
wire n_8984;
wire n_19192;
wire n_5248;
wire n_17786;
wire n_11030;
wire n_20908;
wire n_13495;
wire n_8012;
wire n_12012;
wire n_13777;
wire n_5666;
wire n_18663;
wire n_11368;
wire n_12098;
wire n_19944;
wire n_7988;
wire n_15468;
wire n_13205;
wire n_4448;
wire n_6824;
wire n_8763;
wire n_9370;
wire n_17625;
wire n_20074;
wire n_15553;
wire n_20426;
wire n_16175;
wire n_17737;
wire n_16438;
wire n_13747;
wire n_4776;
wire n_14972;
wire n_10984;
wire n_10144;
wire n_19229;
wire n_3103;
wire n_14439;
wire n_505;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_5682;
wire n_5461;
wire n_12951;
wire n_6164;
wire n_11426;
wire n_3616;
wire n_9484;
wire n_8731;
wire n_2191;
wire n_20830;
wire n_19524;
wire n_7178;
wire n_20043;
wire n_1017;
wire n_12884;
wire n_16056;
wire n_734;
wire n_13414;
wire n_10949;
wire n_310;
wire n_12911;
wire n_8496;
wire n_17280;
wire n_20332;
wire n_2432;
wire n_10156;
wire n_5075;
wire n_14449;
wire n_16273;
wire n_8078;
wire n_19088;
wire n_17523;
wire n_939;
wire n_17705;
wire n_19630;
wire n_1325;
wire n_20893;
wire n_18513;
wire n_1983;
wire n_9141;
wire n_4569;
wire n_10316;
wire n_17281;
wire n_15192;
wire n_10385;
wire n_15775;
wire n_2961;
wire n_15917;
wire n_1923;
wire n_18213;
wire n_13145;
wire n_3631;
wire n_12549;
wire n_1031;
wire n_16003;
wire n_1571;
wire n_12237;
wire n_14586;
wire n_20790;
wire n_252;
wire n_4287;
wire n_9959;
wire n_17499;
wire n_18704;
wire n_14495;
wire n_20155;
wire n_13872;
wire n_8964;
wire n_10611;
wire n_4627;
wire n_15635;
wire n_3590;
wire n_12337;
wire n_19853;
wire n_8247;
wire n_17876;
wire n_14182;
wire n_895;
wire n_15246;
wire n_1639;
wire n_19989;
wire n_20920;
wire n_3295;
wire n_12489;
wire n_12886;
wire n_10321;
wire n_15173;
wire n_5039;
wire n_4265;
wire n_19147;
wire n_15956;
wire n_14884;
wire n_11018;
wire n_19572;
wire n_2269;
wire n_7491;
wire n_14243;
wire n_10909;
wire n_4612;
wire n_17228;
wire n_17782;
wire n_15796;
wire n_6602;
wire n_4958;
wire n_15969;
wire n_8839;
wire n_13627;
wire n_1752;
wire n_4538;
wire n_17378;
wire n_7860;
wire n_4730;
wire n_13364;
wire n_8859;
wire n_4421;
wire n_882;
wire n_2304;
wire n_19710;
wire n_10485;
wire n_8096;
wire n_11946;
wire n_19341;
wire n_289;
wire n_16850;
wire n_19104;
wire n_20685;
wire n_6506;
wire n_2079;
wire n_9705;
wire n_2152;
wire n_14676;
wire n_20213;
wire n_2095;
wire n_15967;
wire n_14355;
wire n_14025;
wire n_8658;
wire n_5944;
wire n_2208;
wire n_15939;
wire n_18554;
wire n_12643;
wire n_11445;
wire n_10592;
wire n_5246;
wire n_19458;
wire n_15022;
wire n_12694;
wire n_20061;
wire n_4305;
wire n_20903;
wire n_2953;
wire n_17187;
wire n_19700;
wire n_18545;
wire n_7273;
wire n_5725;
wire n_5404;
wire n_1507;
wire n_9723;
wire n_16791;
wire n_17923;
wire n_16270;
wire n_2346;
wire n_12506;
wire n_19401;
wire n_3268;
wire n_5616;
wire n_16621;
wire n_10848;
wire n_20289;
wire n_4259;
wire n_2030;
wire n_850;
wire n_12333;
wire n_13502;
wire n_17530;
wire n_6758;
wire n_14801;
wire n_2407;
wire n_17272;
wire n_5288;
wire n_5601;
wire n_15561;
wire n_17181;
wire n_7033;
wire n_17245;
wire n_4178;
wire n_6010;
wire n_12551;
wire n_17355;
wire n_15604;
wire n_8157;
wire n_10990;
wire n_18632;
wire n_8484;
wire n_17400;
wire n_12627;
wire n_12226;
wire n_5294;
wire n_17879;
wire n_9337;
wire n_5955;
wire n_10278;
wire n_2238;
wire n_4793;
wire n_14174;
wire n_10996;
wire n_8692;
wire n_2380;
wire n_16341;
wire n_16244;
wire n_1745;
wire n_14158;
wire n_14218;
wire n_11033;
wire n_19037;
wire n_1088;
wire n_7138;
wire n_766;
wire n_19055;
wire n_7279;
wire n_5184;
wire n_377;
wire n_17651;
wire n_16437;
wire n_10484;
wire n_2547;
wire n_19405;
wire n_4575;
wire n_7137;
wire n_20022;
wire n_3858;
wire n_4589;
wire n_10584;
wire n_8667;
wire n_3220;
wire n_14466;
wire n_11542;
wire n_19823;
wire n_4845;
wire n_9134;
wire n_6654;
wire n_11491;
wire n_4968;
wire n_8807;
wire n_9765;
wire n_20245;
wire n_4038;
wire n_5316;
wire n_953;
wire n_13057;
wire n_1224;
wire n_10324;
wire n_2109;
wire n_20735;
wire n_17727;
wire n_15395;
wire n_795;
wire n_20544;
wire n_1936;
wire n_821;
wire n_1514;
wire n_19455;
wire n_17749;
wire n_569;
wire n_19842;
wire n_11415;
wire n_222;
wire n_4431;
wire n_3347;
wire n_13248;
wire n_17050;
wire n_18888;
wire n_14278;
wire n_19421;
wire n_17978;
wire n_10824;
wire n_3209;
wire n_5220;
wire n_21128;
wire n_6691;
wire n_3948;
wire n_1074;
wire n_1765;
wire n_9132;
wire n_17278;
wire n_206;
wire n_9547;
wire n_2060;
wire n_18444;
wire n_12929;
wire n_136;
wire n_6437;
wire n_2874;
wire n_6684;
wire n_6025;
wire n_16740;
wire n_18874;
wire n_18908;
wire n_17578;
wire n_19694;
wire n_14451;
wire n_10122;
wire n_9762;
wire n_3739;
wire n_16218;
wire n_6062;
wire n_3271;
wire n_20641;
wire n_15414;
wire n_5096;
wire n_20231;
wire n_7905;
wire n_11247;
wire n_7204;
wire n_17318;
wire n_20330;
wire n_6877;
wire n_10116;
wire n_14743;
wire n_16985;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_1378;
wire n_18033;
wire n_5268;
wire n_17684;
wire n_5240;
wire n_5718;
wire n_9915;
wire n_13006;
wire n_1876;
wire n_18631;
wire n_12459;
wire n_19242;
wire n_11075;
wire n_5001;
wire n_700;
wire n_4174;
wire n_18491;
wire n_15516;
wire n_4582;
wire n_20320;
wire n_6520;
wire n_7623;
wire n_380;
wire n_15567;
wire n_19695;
wire n_9335;
wire n_20068;
wire n_1108;
wire n_17406;
wire n_16090;
wire n_17949;
wire n_6637;
wire n_11510;
wire n_16843;
wire n_17779;
wire n_10185;
wire n_3909;
wire n_10809;
wire n_13316;
wire n_13140;
wire n_15308;
wire n_5541;
wire n_12501;
wire n_407;
wire n_2810;
wire n_12755;
wire n_20580;
wire n_6703;
wire n_1555;
wire n_10657;
wire n_20713;
wire n_10627;
wire n_762;
wire n_1253;
wire n_19187;
wire n_7265;
wire n_14805;
wire n_11516;
wire n_11520;
wire n_15376;
wire n_6878;
wire n_11137;
wire n_8181;
wire n_16733;
wire n_6527;
wire n_2748;
wire n_11544;
wire n_14234;
wire n_1376;
wire n_20349;
wire n_20967;
wire n_9253;
wire n_6533;
wire n_14126;
wire n_18831;
wire n_7164;
wire n_15164;
wire n_1506;
wire n_18671;
wire n_12011;
wire n_5300;
wire n_11268;
wire n_13707;
wire n_12742;
wire n_20835;
wire n_9953;
wire n_10315;
wire n_18688;
wire n_12317;
wire n_18751;
wire n_3510;
wire n_7046;
wire n_13928;
wire n_17571;
wire n_18446;
wire n_21020;
wire n_8940;
wire n_15541;
wire n_18948;
wire n_18026;
wire n_16727;
wire n_12590;
wire n_14503;
wire n_17211;
wire n_11213;
wire n_19252;
wire n_13519;
wire n_2100;
wire n_5538;
wire n_16314;
wire n_944;
wire n_19468;
wire n_2888;
wire n_1920;
wire n_7811;
wire n_7097;
wire n_2567;
wire n_20158;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_14130;
wire n_17485;
wire n_6713;
wire n_13163;
wire n_12953;
wire n_17044;
wire n_2066;
wire n_2762;
wire n_7851;
wire n_13106;
wire n_13776;
wire n_12222;
wire n_6866;
wire n_11412;
wire n_7332;
wire n_20111;
wire n_471;
wire n_7477;
wire n_19406;
wire n_10268;
wire n_13640;
wire n_6415;
wire n_12397;
wire n_2021;
wire n_1563;
wire n_3052;
wire n_16104;
wire n_1633;
wire n_4621;
wire n_13086;
wire n_183;
wire n_2261;
wire n_12613;
wire n_20260;
wire n_9079;
wire n_9782;
wire n_10049;
wire n_13012;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_13099;
wire n_9950;
wire n_19597;
wire n_11580;
wire n_3867;
wire n_3397;
wire n_12683;
wire n_1646;
wire n_6392;
wire n_13389;
wire n_11642;
wire n_6720;
wire n_11752;
wire n_10785;
wire n_14726;
wire n_13439;
wire n_17940;
wire n_3971;
wire n_14415;
wire n_20953;
wire n_286;
wire n_4979;
wire n_2113;
wire n_15201;
wire n_3711;
wire n_19066;
wire n_14903;
wire n_9536;
wire n_9848;
wire n_6571;
wire n_16159;
wire n_8324;
wire n_20338;
wire n_9841;
wire n_10147;
wire n_9772;
wire n_1496;
wire n_2812;
wire n_14847;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_8014;
wire n_12213;
wire n_12646;
wire n_2132;
wire n_14159;
wire n_5991;
wire n_8623;
wire n_18404;
wire n_8651;
wire n_10699;
wire n_5000;
wire n_1795;
wire n_14358;
wire n_5132;
wire n_3498;
wire n_2350;
wire n_19502;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_9591;
wire n_7171;
wire n_2187;
wire n_1413;
wire n_8413;
wire n_2481;
wire n_158;
wire n_9471;
wire n_20169;
wire n_20737;
wire n_21042;
wire n_1365;
wire n_3675;
wire n_20141;
wire n_12601;
wire n_16361;
wire n_18708;
wire n_8069;
wire n_320;
wire n_10743;
wire n_6432;
wire n_20189;
wire n_2055;
wire n_17829;
wire n_10481;
wire n_13562;
wire n_1609;
wire n_20275;
wire n_7589;
wire n_13568;
wire n_4447;
wire n_218;
wire n_9832;
wire n_5793;
wire n_18456;
wire n_3057;
wire n_12856;
wire n_18907;
wire n_6699;
wire n_13683;
wire n_13630;
wire n_20695;
wire n_3983;
wire n_19626;
wire n_8254;
wire n_10141;
wire n_14661;
wire n_10305;
wire n_16801;
wire n_16728;
wire n_326;
wire n_3773;
wire n_20667;
wire n_1278;
wire n_11429;
wire n_9033;
wire n_14624;
wire n_17576;
wire n_11908;
wire n_3788;
wire n_20781;
wire n_16494;
wire n_18099;
wire n_20707;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_9247;
wire n_3349;
wire n_16739;
wire n_18778;
wire n_7466;
wire n_1205;
wire n_2716;
wire n_11660;
wire n_15675;
wire n_3439;
wire n_18797;
wire n_19036;
wire n_12355;
wire n_3602;
wire n_233;
wire n_8954;
wire n_19640;
wire n_19008;
wire n_12458;
wire n_20766;
wire n_7494;
wire n_1586;
wire n_11280;
wire n_16435;
wire n_16589;
wire n_9680;
wire n_8398;
wire n_5641;
wire n_13046;
wire n_16292;
wire n_4461;
wire n_2660;
wire n_3426;
wire n_17360;
wire n_8528;
wire n_13644;
wire n_20895;
wire n_20241;
wire n_8475;
wire n_17240;
wire n_297;
wire n_20816;
wire n_13545;
wire n_3896;
wire n_14913;
wire n_13197;
wire n_9054;
wire n_4551;
wire n_178;
wire n_10117;
wire n_13252;
wire n_6956;
wire n_10126;
wire n_2284;
wire n_11920;
wire n_19879;
wire n_5420;
wire n_6497;
wire n_16915;
wire n_20628;
wire n_14237;
wire n_6701;
wire n_1239;
wire n_16770;
wire n_10209;
wire n_560;
wire n_8558;
wire n_13769;
wire n_18464;
wire n_9593;
wire n_18670;
wire n_14433;
wire n_3423;
wire n_13626;
wire n_17344;
wire n_10299;
wire n_21055;
wire n_16732;
wire n_14195;
wire n_1800;
wire n_11811;
wire n_12417;
wire n_18505;
wire n_10618;
wire n_2946;
wire n_16691;
wire n_7953;
wire n_16086;
wire n_6876;
wire n_15746;
wire n_17470;
wire n_16446;
wire n_1734;
wire n_7193;
wire n_2840;
wire n_4482;
wire n_5957;
wire n_18772;
wire n_20020;
wire n_20152;
wire n_3024;
wire n_9879;
wire n_8647;
wire n_6362;
wire n_17119;
wire n_8543;
wire n_1854;
wire n_666;
wire n_15637;
wire n_11184;
wire n_6833;
wire n_785;
wire n_14720;
wire n_999;
wire n_12985;
wire n_12232;
wire n_15316;
wire n_5085;
wire n_19926;
wire n_4113;
wire n_13729;
wire n_6430;
wire n_11435;
wire n_873;
wire n_16902;
wire n_6296;
wire n_342;
wire n_5602;
wire n_18828;
wire n_20194;
wire n_11120;
wire n_20481;
wire n_10895;
wire n_4865;
wire n_15611;
wire n_13002;
wire n_5822;
wire n_17095;
wire n_3586;
wire n_4160;
wire n_15111;
wire n_15151;
wire n_6385;
wire n_12571;
wire n_4137;
wire n_1078;
wire n_13022;
wire n_15949;
wire n_4545;
wire n_8200;
wire n_15771;
wire n_15590;
wire n_5713;
wire n_9905;
wire n_16971;
wire n_18628;
wire n_14142;
wire n_8586;
wire n_618;
wire n_12540;
wire n_12001;
wire n_4385;
wire n_7779;
wire n_13275;
wire n_11489;
wire n_20807;
wire n_2337;
wire n_15753;
wire n_16582;
wire n_13760;
wire n_12479;
wire n_8370;
wire n_3732;
wire n_19102;
wire n_17583;
wire n_18925;
wire n_13663;
wire n_10569;
wire n_4558;
wire n_14055;
wire n_16153;
wire n_7349;
wire n_9875;
wire n_10713;
wire n_19874;
wire n_16325;
wire n_12306;
wire n_12637;
wire n_7122;
wire n_180;
wire n_10203;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_11000;
wire n_9803;
wire n_15738;
wire n_8564;
wire n_12114;
wire n_8343;
wire n_7828;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_15106;
wire n_20101;
wire n_13550;
wire n_19520;
wire n_985;
wire n_5506;
wire n_8042;
wire n_16382;
wire n_7727;
wire n_5908;
wire n_17828;
wire n_12325;
wire n_8379;
wire n_643;
wire n_8034;
wire n_17771;
wire n_2383;
wire n_10225;
wire n_682;
wire n_9474;
wire n_7702;
wire n_17533;
wire n_14930;
wire n_3390;
wire n_16374;
wire n_2298;
wire n_19913;
wire n_2320;
wire n_19866;
wire n_11523;
wire n_17370;
wire n_18320;
wire n_8362;
wire n_6971;
wire n_3336;
wire n_8632;
wire n_7739;
wire n_7945;
wire n_8361;
wire n_5903;
wire n_3541;
wire n_14937;
wire n_12344;
wire n_18664;
wire n_725;
wire n_8611;
wire n_6540;
wire n_16360;
wire n_2198;
wire n_15634;
wire n_3067;
wire n_20711;
wire n_473;
wire n_1852;
wire n_5912;
wire n_6086;
wire n_818;
wire n_5803;
wire n_8878;
wire n_5270;
wire n_8492;
wire n_4301;
wire n_10392;
wire n_19197;
wire n_15076;
wire n_6820;
wire n_879;
wire n_11245;
wire n_7107;
wire n_14225;
wire n_7610;
wire n_18913;
wire n_9921;
wire n_1050;
wire n_11005;
wire n_2578;
wire n_1201;
wire n_17432;
wire n_7823;
wire n_8833;
wire n_14605;
wire n_6157;
wire n_2665;
wire n_4879;
wire n_19019;
wire n_1090;
wire n_9894;
wire n_9274;
wire n_20186;
wire n_4927;
wire n_18905;
wire n_14285;
wire n_12171;
wire n_1801;
wire n_20407;
wire n_8690;
wire n_18581;
wire n_16826;
wire n_5390;
wire n_17032;
wire n_5267;
wire n_15377;
wire n_1641;
wire n_16562;
wire n_4151;
wire n_6923;
wire n_8009;
wire n_8195;
wire n_8588;
wire n_843;
wire n_16027;
wire n_17563;
wire n_13520;
wire n_4682;
wire n_11012;
wire n_6673;
wire n_14480;
wire n_14024;
wire n_11798;
wire n_15312;
wire n_6534;
wire n_8805;
wire n_15576;
wire n_1955;
wire n_6246;
wire n_10989;
wire n_14702;
wire n_13315;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_20644;
wire n_5207;
wire n_7934;
wire n_2658;
wire n_12957;
wire n_4601;
wire n_18001;
wire n_4518;
wire n_7009;
wire n_3376;
wire n_683;
wire n_7463;
wire n_19319;
wire n_18485;
wire n_4308;
wire n_11851;
wire n_16068;
wire n_1420;
wire n_21009;
wire n_19139;
wire n_20367;
wire n_13628;
wire n_2833;
wire n_7398;
wire n_12757;
wire n_5223;
wire n_20229;
wire n_414;
wire n_571;
wire n_11738;
wire n_11595;
wire n_5801;
wire n_14163;
wire n_16723;
wire n_12349;
wire n_6054;
wire n_3405;
wire n_2313;
wire n_11603;
wire n_17167;
wire n_19815;
wire n_1022;
wire n_12577;
wire n_3532;
wire n_2609;
wire n_8169;
wire n_11802;
wire n_9984;
wire n_3131;
wire n_820;
wire n_20343;
wire n_12135;
wire n_15761;
wire n_7969;
wire n_8793;
wire n_17894;
wire n_10388;
wire n_6312;
wire n_13108;
wire n_20670;
wire n_15701;
wire n_10510;
wire n_2624;
wire n_2054;
wire n_1552;
wire n_13429;
wire n_6193;
wire n_13897;
wire n_6734;
wire n_6535;
wire n_17174;
wire n_15893;
wire n_17915;
wire n_8059;
wire n_19602;
wire n_9562;
wire n_17780;
wire n_17595;
wire n_18210;
wire n_493;
wire n_17655;
wire n_6014;
wire n_14016;
wire n_10241;
wire n_15451;
wire n_6457;
wire n_15953;
wire n_9955;
wire n_8372;
wire n_6270;
wire n_8737;
wire n_5996;
wire n_7288;
wire n_19329;
wire n_19382;
wire n_6276;
wire n_739;
wire n_1028;
wire n_15661;
wire n_12328;
wire n_530;
wire n_8723;
wire n_12559;
wire n_10767;
wire n_5652;
wire n_17254;
wire n_1645;
wire n_16235;
wire n_15386;
wire n_3301;
wire n_12109;
wire n_2910;
wire n_14457;
wire n_9531;
wire n_10521;
wire n_6934;
wire n_4401;
wire n_12058;
wire n_2586;
wire n_19239;
wire n_268;
wire n_10872;
wire n_12083;
wire n_19618;
wire n_3100;
wire n_10374;
wire n_12045;
wire n_10345;
wire n_8959;
wire n_20259;
wire n_12471;
wire n_4973;
wire n_13781;
wire n_13802;
wire n_14736;
wire n_4402;
wire n_15351;
wire n_16619;
wire n_2487;
wire n_1834;
wire n_10601;
wire n_2534;
wire n_6211;
wire n_8109;
wire n_3576;
wire n_12040;
wire n_9389;
wire n_15562;
wire n_19641;
wire n_8725;
wire n_8007;
wire n_13911;
wire n_14313;
wire n_17560;
wire n_19865;
wire n_18791;
wire n_3570;
wire n_17404;
wire n_18836;
wire n_2793;
wire n_6764;
wire n_7871;
wire n_541;
wire n_16679;
wire n_15982;
wire n_20192;
wire n_7016;
wire n_17019;
wire n_12100;
wire n_4554;
wire n_7571;
wire n_13584;
wire n_13107;
wire n_1663;
wire n_10774;
wire n_6955;
wire n_5952;
wire n_16253;
wire n_10407;
wire n_10577;
wire n_2086;
wire n_14481;
wire n_16171;
wire n_15148;
wire n_8494;
wire n_7919;
wire n_663;
wire n_2966;
wire n_19633;
wire n_18156;
wire n_20611;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_13367;
wire n_20757;
wire n_10843;
wire n_10771;
wire n_18882;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_19827;
wire n_2543;
wire n_11983;
wire n_17065;
wire n_15885;
wire n_15053;
wire n_4875;
wire n_13284;
wire n_8903;
wire n_16946;
wire n_2758;
wire n_12596;
wire n_17155;
wire n_5036;
wire n_17777;
wire n_11215;
wire n_5790;
wire n_2471;
wire n_1067;
wire n_19702;
wire n_11591;
wire n_5118;
wire n_4849;
wire n_2039;
wire n_7133;
wire n_761;
wire n_19316;
wire n_8882;
wire n_14308;
wire n_18279;
wire n_17788;
wire n_15532;
wire n_2734;
wire n_13600;
wire n_8067;
wire n_8385;
wire n_20288;
wire n_18765;
wire n_4917;
wire n_8142;
wire n_19516;
wire n_15381;
wire n_15090;
wire n_11204;
wire n_153;
wire n_648;
wire n_6836;
wire n_12939;
wire n_10415;
wire n_17105;
wire n_18276;
wire n_12374;
wire n_17922;
wire n_17150;
wire n_17519;
wire n_15398;
wire n_16081;
wire n_10227;
wire n_16767;
wire n_2463;
wire n_1792;
wire n_504;
wire n_2062;
wire n_4489;
wire n_822;
wire n_17466;
wire n_17476;
wire n_5472;
wire n_10884;
wire n_13375;
wire n_839;
wire n_7236;
wire n_8345;
wire n_16722;
wire n_1575;
wire n_9343;
wire n_19669;
wire n_9131;
wire n_13286;
wire n_3903;
wire n_5072;
wire n_8529;
wire n_13384;
wire n_11325;
wire n_17342;
wire n_18885;
wire n_10325;
wire n_6361;
wire n_17251;
wire n_1315;
wire n_997;
wire n_18619;
wire n_5940;
wire n_5260;
wire n_6751;
wire n_6232;
wire n_20995;
wire n_15144;
wire n_18186;
wire n_2990;
wire n_2034;
wire n_10505;
wire n_3932;
wire n_12979;
wire n_14140;
wire n_7457;
wire n_6736;
wire n_19337;
wire n_15262;
wire n_11672;
wire n_19089;
wire n_9982;
wire n_11552;
wire n_13682;
wire n_19385;
wire n_20447;
wire n_7639;
wire n_6214;
wire n_9006;
wire n_9221;
wire n_18717;
wire n_19542;
wire n_4365;
wire n_10514;
wire n_14603;
wire n_7049;
wire n_18416;
wire n_6143;
wire n_2736;
wire n_10091;
wire n_7749;
wire n_11195;
wire n_20547;
wire n_6225;
wire n_4373;
wire n_8860;
wire n_2664;
wire n_20616;
wire n_12401;
wire n_4154;
wire n_13304;
wire n_10593;
wire n_15078;
wire n_16608;
wire n_2360;
wire n_18076;
wire n_4453;
wire n_15484;
wire n_8686;
wire n_8563;
wire n_4571;
wire n_20091;
wire n_10197;
wire n_4886;
wire n_6198;
wire n_15792;
wire n_10950;
wire n_9411;
wire n_1019;
wire n_8765;
wire n_15946;
wire n_5164;
wire n_13688;
wire n_19475;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_6827;
wire n_19099;
wire n_1768;
wire n_2369;
wire n_11679;
wire n_17058;
wire n_6281;
wire n_13005;
wire n_2587;
wire n_17322;
wire n_13313;
wire n_18206;
wire n_9675;
wire n_6822;
wire n_4956;
wire n_255;
wire n_18917;
wire n_16503;
wire n_5878;
wire n_18709;
wire n_10075;
wire n_2674;
wire n_17045;
wire n_1613;
wire n_20844;
wire n_17790;
wire n_14351;
wire n_12873;
wire n_12767;
wire n_1779;
wire n_17892;
wire n_18030;
wire n_19155;
wire n_19425;
wire n_9511;
wire n_20235;
wire n_16386;
wire n_10798;
wire n_2673;
wire n_11630;
wire n_14185;
wire n_18881;
wire n_4678;
wire n_13211;
wire n_16937;
wire n_2548;
wire n_9622;
wire n_12198;
wire n_9761;
wire n_7646;
wire n_3779;
wire n_14870;
wire n_12617;
wire n_17707;
wire n_1063;
wire n_19158;
wire n_10669;
wire n_8790;
wire n_21072;
wire n_18029;
wire n_8305;
wire n_4303;
wire n_1912;
wire n_15800;
wire n_1891;
wire n_6634;
wire n_12666;
wire n_17189;
wire n_4868;
wire n_11617;
wire n_19605;
wire n_20184;
wire n_17375;
wire n_14969;
wire n_13565;
wire n_8127;
wire n_5217;
wire n_9115;
wire n_7861;
wire n_472;
wire n_13788;
wire n_4245;
wire n_11422;
wire n_2524;
wire n_208;
wire n_3894;
wire n_12594;
wire n_10542;
wire n_275;
wire n_11376;
wire n_20548;
wire n_5750;
wire n_7648;
wire n_1232;
wire n_996;
wire n_10752;
wire n_5654;
wire n_10868;
wire n_9594;
wire n_2229;
wire n_6400;
wire n_5554;
wire n_9503;
wire n_250;
wire n_18768;
wire n_7551;
wire n_11793;
wire n_4599;
wire n_4222;
wire n_10017;
wire n_1434;
wire n_8093;
wire n_20380;
wire n_9385;
wire n_15104;
wire n_7737;
wire n_20753;
wire n_523;
wire n_3249;
wire n_15971;
wire n_16880;
wire n_2915;
wire n_10572;
wire n_17204;
wire n_9885;
wire n_8115;
wire n_20663;
wire n_4047;
wire n_11670;
wire n_484;
wire n_10642;
wire n_2719;
wire n_10517;
wire n_13852;
wire n_12451;
wire n_16982;
wire n_3033;
wire n_9182;
wire n_10620;
wire n_18091;
wire n_1582;
wire n_8182;
wire n_20728;
wire n_4417;
wire n_796;
wire n_1374;
wire n_16955;
wire n_9581;
wire n_18525;
wire n_17352;
wire n_20956;
wire n_6158;
wire n_15028;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_14734;
wire n_2509;
wire n_5486;
wire n_7260;
wire n_6894;
wire n_6843;
wire n_5851;
wire n_5432;
wire n_20834;
wire n_1463;
wire n_7625;
wire n_6806;
wire n_924;
wire n_9542;
wire n_16486;
wire n_3517;
wire n_20646;
wire n_10829;
wire n_11356;
wire n_524;
wire n_16753;
wire n_1214;
wire n_20324;
wire n_3526;
wire n_17646;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_11678;
wire n_6088;
wire n_10236;
wire n_4683;
wire n_11162;
wire n_18690;
wire n_2873;
wire n_15698;
wire n_3330;
wire n_3514;
wire n_18133;
wire n_1457;
wire n_14402;
wire n_13552;
wire n_8552;
wire n_4600;
wire n_14389;
wire n_9403;
wire n_14558;
wire n_18681;
wire n_9878;
wire n_10139;
wire n_17312;
wire n_270;
wire n_4106;
wire n_20850;
wire n_285;
wire n_12548;
wire n_202;
wire n_9735;
wire n_20140;
wire n_754;
wire n_2323;
wire n_7327;
wire n_12727;
wire n_1277;
wire n_19220;
wire n_5998;
wire n_8318;
wire n_14742;
wire n_20560;
wire n_19094;
wire n_4954;
wire n_15707;
wire n_19410;
wire n_167;
wire n_2906;
wire n_6250;
wire n_12372;
wire n_11392;
wire n_3283;
wire n_15597;
wire n_17259;
wire n_259;
wire n_15066;
wire n_18764;
wire n_18919;
wire n_7864;
wire n_10650;
wire n_4734;
wire n_7955;
wire n_2370;
wire n_2914;
wire n_17953;
wire n_12952;
wire n_6858;
wire n_6050;
wire n_18445;
wire n_4515;
wire n_10417;
wire n_2539;
wire n_8620;
wire n_1145;
wire n_4809;
wire n_4012;
wire n_10253;
wire n_16051;
wire n_15533;
wire n_5212;
wire n_1207;
wire n_13136;
wire n_6823;
wire n_3606;
wire n_12449;
wire n_15261;
wire n_11966;
wire n_14205;
wire n_4320;
wire n_7223;
wire n_14266;
wire n_12770;
wire n_5251;
wire n_3324;
wire n_10977;
wire n_19508;
wire n_17851;
wire n_13220;
wire n_8141;
wire n_3230;
wire n_12826;
wire n_6024;
wire n_4768;
wire n_16953;
wire n_5368;
wire n_3828;
wire n_16773;
wire n_17692;
wire n_16973;
wire n_1850;
wire n_9908;
wire n_8004;
wire n_14763;
wire n_3607;
wire n_2098;
wire n_2616;
wire n_10212;
wire n_20144;
wire n_438;
wire n_14208;
wire n_6714;
wire n_10539;
wire n_12937;
wire n_7446;
wire n_2902;
wire n_4360;
wire n_9317;
wire n_17146;
wire n_8198;
wire n_16168;
wire n_19003;
wire n_12201;
wire n_16755;
wire n_13240;
wire n_19159;
wire n_1021;
wire n_13187;
wire n_13594;
wire n_10516;
wire n_1142;
wire n_11675;
wire n_260;
wire n_7523;
wire n_14035;
wire n_10432;
wire n_14345;
wire n_7559;
wire n_9037;
wire n_20879;
wire n_1599;
wire n_11988;
wire n_18823;
wire n_18921;
wire n_19976;
wire n_2527;
wire n_15172;
wire n_7257;
wire n_3126;
wire n_20889;
wire n_2759;
wire n_10869;
wire n_5007;
wire n_4881;
wire n_10314;
wire n_16945;
wire n_4737;
wire n_9218;
wire n_4357;
wire n_19628;
wire n_7729;
wire n_20441;
wire n_12373;
wire n_19175;
wire n_15544;
wire n_21028;
wire n_3588;
wire n_16897;
wire n_5274;
wire n_6399;
wire n_17474;
wire n_5939;
wire n_9506;
wire n_13629;
wire n_135;
wire n_11569;
wire n_10256;
wire n_4775;
wire n_15976;
wire n_1691;
wire n_8250;
wire n_14315;
wire n_20700;
wire n_21018;
wire n_12181;
wire n_6648;
wire n_12115;
wire n_804;
wire n_12567;
wire n_3093;
wire n_12175;
wire n_17783;
wire n_6910;
wire n_955;
wire n_8466;
wire n_18737;
wire n_9015;
wire n_15482;
wire n_2166;
wire n_4709;
wire n_12754;
wire n_4223;
wire n_20236;
wire n_19895;
wire n_3538;
wire n_11990;
wire n_3839;
wire n_5490;
wire n_13728;
wire n_3875;
wire n_8876;
wire n_19936;
wire n_2415;
wire n_20335;
wire n_3120;
wire n_9070;
wire n_15993;
wire n_16709;
wire n_4794;
wire n_9933;
wire n_15108;
wire n_5215;
wire n_437;
wire n_18441;
wire n_19140;
wire n_10874;
wire n_9486;
wire n_14113;
wire n_12425;
wire n_8267;
wire n_2462;
wire n_6773;
wire n_16814;
wire n_15758;
wire n_615;
wire n_4838;
wire n_19785;
wire n_3604;
wire n_8545;
wire n_17588;
wire n_19621;
wire n_12300;
wire n_159;
wire n_12527;
wire n_21123;
wire n_12110;
wire n_21106;
wire n_9790;
wire n_11404;
wire n_4267;
wire n_20171;
wire n_16026;
wire n_7793;
wire n_9053;
wire n_16337;
wire n_2083;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_11007;
wire n_9880;
wire n_18886;
wire n_15859;
wire n_19670;
wire n_7425;
wire n_5958;
wire n_18353;
wire n_9499;
wire n_7829;
wire n_18626;
wire n_10081;
wire n_799;
wire n_10145;
wire n_8262;
wire n_10167;
wire n_12656;
wire n_5809;
wire n_934;
wire n_7531;
wire n_12219;
wire n_12729;
wire n_356;
wire n_13921;
wire n_6473;
wire n_13345;
wire n_4806;
wire n_4015;
wire n_15129;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_13216;
wire n_4219;
wire n_4723;
wire n_11226;
wire n_9371;
wire n_8701;
wire n_2896;
wire n_1042;
wire n_2311;
wire n_13398;
wire n_14148;
wire n_12644;
wire n_6290;
wire n_20965;
wire n_205;
wire n_20336;
wire n_4234;
wire n_17382;
wire n_19071;
wire n_1363;
wire n_1111;
wire n_5821;
wire n_6622;
wire n_19513;
wire n_5522;
wire n_13169;
wire n_10287;
wire n_20806;
wire n_3699;
wire n_16584;
wire n_7125;
wire n_6532;
wire n_9479;
wire n_6267;
wire n_9480;
wire n_20318;
wire n_19453;
wire n_8085;
wire n_2757;
wire n_2168;
wire n_15026;
wire n_20836;
wire n_14273;
wire n_19002;
wire n_7203;
wire n_9641;
wire n_10039;
wire n_13866;
wire n_1259;
wire n_20857;
wire n_1177;
wire n_18412;
wire n_5771;
wire n_18812;
wire n_8887;
wire n_1618;
wire n_12091;
wire n_15716;
wire n_4911;
wire n_15168;
wire n_5516;
wire n_18978;
wire n_3019;
wire n_11826;
wire n_19745;
wire n_18942;
wire n_11825;
wire n_9111;
wire n_6772;
wire n_15499;
wire n_9618;
wire n_17794;
wire n_10383;
wire n_10856;
wire n_20992;
wire n_14532;
wire n_12935;
wire n_18981;
wire n_9065;
wire n_14463;
wire n_17124;
wire n_6159;
wire n_5857;
wire n_7979;
wire n_9674;
wire n_6617;
wire n_814;
wire n_18462;
wire n_5120;
wire n_19665;
wire n_2399;
wire n_16558;
wire n_8467;
wire n_18308;
wire n_20610;
wire n_19750;
wire n_11093;
wire n_2027;
wire n_16205;
wire n_17202;
wire n_10303;
wire n_15071;
wire n_3922;
wire n_8640;
wire n_1467;
wire n_7447;
wire n_247;
wire n_2159;
wire n_8431;
wire n_1744;
wire n_5916;
wire n_10421;
wire n_14376;
wire n_13855;
wire n_5099;
wire n_681;
wire n_11179;
wire n_19422;
wire n_18393;
wire n_14777;
wire n_9416;
wire n_7365;
wire n_20635;
wire n_2599;
wire n_3988;
wire n_8089;
wire n_2075;
wire n_13771;
wire n_13845;
wire n_11921;
wire n_3761;
wire n_15443;
wire n_14224;
wire n_10285;
wire n_7275;
wire n_19501;
wire n_15039;
wire n_12099;
wire n_6856;
wire n_13572;
wire n_777;
wire n_10084;
wire n_8541;
wire n_12924;
wire n_17148;
wire n_8762;
wire n_18682;
wire n_3035;
wire n_17285;
wire n_13104;
wire n_15176;
wire n_11647;
wire n_6240;
wire n_15222;
wire n_2254;
wire n_6693;
wire n_10101;
wire n_3418;
wire n_10566;
wire n_8188;
wire n_19046;
wire n_16450;
wire n_6586;
wire n_17164;
wire n_19655;
wire n_8923;
wire n_20296;
wire n_281;
wire n_3326;
wire n_11389;
wire n_8624;
wire n_15150;
wire n_12429;
wire n_18290;
wire n_15547;
wire n_1883;
wire n_11315;
wire n_3224;
wire n_1969;
wire n_20160;
wire n_7429;
wire n_13506;
wire n_20605;
wire n_6468;
wire n_7709;
wire n_12923;
wire n_15112;
wire n_16931;
wire n_10362;
wire n_1222;
wire n_19945;
wire n_19288;
wire n_14213;
wire n_11962;
wire n_3803;
wire n_13885;
wire n_14928;
wire n_7782;
wire n_7432;
wire n_4913;
wire n_18732;
wire n_10093;
wire n_13924;
wire n_4428;
wire n_745;
wire n_9684;
wire n_12591;
wire n_4463;
wire n_19182;
wire n_10600;
wire n_11994;
wire n_8175;
wire n_6810;
wire n_11316;
wire n_17386;
wire n_15938;
wire n_18904;
wire n_12948;
wire n_18306;
wire n_16517;
wire n_15636;
wire n_2690;
wire n_3090;
wire n_12467;
wire n_12756;
wire n_11463;
wire n_20455;
wire n_17209;
wire n_18793;
wire n_6305;
wire n_14641;
wire n_17335;
wire n_11069;
wire n_15751;
wire n_10894;
wire n_7412;
wire n_8168;
wire n_5045;
wire n_5237;
wire n_15465;
wire n_7751;
wire n_20900;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_13603;
wire n_8873;
wire n_10311;
wire n_18461;
wire n_7591;
wire n_3564;
wire n_5769;
wire n_7911;
wire n_3795;
wire n_17293;
wire n_11586;
wire n_11786;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2959;
wire n_6239;
wire n_10181;
wire n_15950;
wire n_5768;
wire n_11330;
wire n_6199;
wire n_3282;
wire n_852;
wire n_4192;
wire n_11979;
wire n_12253;
wire n_15380;
wire n_1748;
wire n_6789;
wire n_1466;
wire n_11888;
wire n_2581;
wire n_15902;
wire n_9259;
wire n_16366;
wire n_10755;
wire n_14274;
wire n_11835;
wire n_10525;
wire n_12776;
wire n_7405;
wire n_3650;
wire n_6825;
wire n_15282;
wire n_7614;
wire n_9150;
wire n_6952;
wire n_1480;
wire n_17194;
wire n_20396;
wire n_14907;
wire n_6173;
wire n_16588;
wire n_4190;
wire n_3060;
wire n_11048;
wire n_11933;
wire n_6486;
wire n_11900;
wire n_12620;
wire n_11106;
wire n_19275;
wire n_10983;
wire n_11266;
wire n_15659;
wire n_12673;
wire n_5017;
wire n_18729;
wire n_736;
wire n_14549;
wire n_2265;
wire n_19299;
wire n_1475;
wire n_3174;
wire n_19469;
wire n_3314;
wire n_14798;
wire n_18114;
wire n_15023;
wire n_13030;
wire n_16643;
wire n_3789;
wire n_12324;
wire n_12817;
wire n_11255;
wire n_16511;
wire n_18592;
wire n_11751;
wire n_10834;
wire n_8577;
wire n_9361;
wire n_16828;
wire n_6626;
wire n_4537;
wire n_10890;
wire n_5838;
wire n_771;
wire n_14188;
wire n_3893;
wire n_18094;
wire n_2307;
wire n_20587;
wire n_12316;
wire n_8952;
wire n_3453;
wire n_6980;
wire n_18895;
wire n_17724;
wire n_15506;
wire n_18424;
wire n_1492;
wire n_4065;
wire n_16689;
wire n_15572;
wire n_12949;
wire n_20025;
wire n_1324;
wire n_20339;
wire n_7179;
wire n_13499;
wire n_19009;
wire n_4279;
wire n_16925;
wire n_13560;
wire n_6257;
wire n_17500;
wire n_18912;
wire n_14073;
wire n_16410;
wire n_2698;
wire n_15693;
wire n_17255;
wire n_7658;
wire n_20677;
wire n_2329;
wire n_3455;
wire n_20714;
wire n_18974;
wire n_10921;
wire n_10177;
wire n_6286;
wire n_15677;
wire n_17070;
wire n_11915;
wire n_1987;
wire n_7217;
wire n_2368;
wire n_6377;
wire n_10492;
wire n_16176;
wire n_12061;
wire n_5401;
wire n_4595;
wire n_20261;
wire n_16048;
wire n_19631;
wire n_5816;
wire n_790;
wire n_14175;
wire n_15373;
wire n_20480;
wire n_18002;
wire n_5543;
wire n_12359;
wire n_15328;
wire n_4054;
wire n_17421;
wire n_13615;
wire n_10741;
wire n_2477;
wire n_10037;
wire n_8949;
wire n_2279;
wire n_10760;
wire n_9454;
wire n_11838;
wire n_4732;
wire n_14768;
wire n_5942;
wire n_5764;
wire n_13702;
wire n_8983;
wire n_4969;
wire n_8121;
wire n_11100;
wire n_15283;
wire n_20071;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_18808;
wire n_20415;
wire n_13867;
wire n_566;
wire n_2607;
wire n_11632;
wire n_3343;
wire n_7255;
wire n_3309;
wire n_19279;
wire n_173;
wire n_10658;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_17235;
wire n_3134;
wire n_4909;
wire n_14399;
wire n_15931;
wire n_3769;
wire n_8194;
wire n_17126;
wire n_4070;
wire n_9900;
wire n_12033;
wire n_14534;
wire n_16489;
wire n_13447;
wire n_7647;
wire n_12465;
wire n_14771;
wire n_5868;
wire n_10808;
wire n_7145;
wire n_3667;
wire n_20590;
wire n_8448;
wire n_5257;
wire n_12684;
wire n_13319;
wire n_9489;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_20591;
wire n_13019;
wire n_6961;
wire n_576;
wire n_8732;
wire n_14610;
wire n_9359;
wire n_4368;
wire n_5272;
wire n_16816;
wire n_6919;
wire n_19451;
wire n_8420;
wire n_4430;
wire n_3238;
wire n_18017;
wire n_18887;
wire n_4544;
wire n_3175;
wire n_7809;
wire n_16804;
wire n_5811;
wire n_2886;
wire n_16498;
wire n_10452;
wire n_8746;
wire n_10051;
wire n_3006;
wire n_4531;
wire n_12498;
wire n_9401;
wire n_543;
wire n_11335;
wire n_12625;
wire n_3456;
wire n_4532;
wire n_7564;
wire n_10396;
wire n_10955;
wire n_8185;
wire n_13062;
wire n_6633;
wire n_14931;
wire n_16847;
wire n_10308;
wire n_847;
wire n_17183;
wire n_12532;
wire n_15974;
wire n_14051;
wire n_4257;
wire n_7636;
wire n_4341;
wire n_20623;
wire n_5480;
wire n_12876;
wire n_8066;
wire n_18695;
wire n_12544;
wire n_13793;
wire n_6425;
wire n_14594;
wire n_10581;
wire n_20474;
wire n_519;
wire n_11724;
wire n_11507;
wire n_18703;
wire n_10647;
wire n_19932;
wire n_20664;
wire n_16413;
wire n_7301;
wire n_15824;
wire n_7262;
wire n_15089;
wire n_17490;
wire n_10769;
wire n_1739;
wire n_2642;
wire n_12215;
wire n_17564;
wire n_13218;
wire n_17967;
wire n_1789;
wire n_14965;
wire n_2174;
wire n_4209;
wire n_6282;
wire n_17082;
wire n_11800;
wire n_9870;
wire n_18481;
wire n_13396;
wire n_2046;
wire n_7059;
wire n_14947;
wire n_1606;
wire n_5600;
wire n_395;
wire n_20636;
wire n_6737;
wire n_213;
wire n_20802;
wire n_4888;
wire n_5767;
wire n_7670;
wire n_17904;
wire n_17681;
wire n_3991;
wire n_13813;
wire n_17977;
wire n_16944;
wire n_8505;
wire n_15509;
wire n_1617;
wire n_10157;
wire n_2600;
wire n_10923;
wire n_10038;
wire n_4759;
wire n_14666;
wire n_18635;
wire n_14793;
wire n_16057;
wire n_15913;
wire n_4887;
wire n_3751;
wire n_16901;
wire n_9229;
wire n_14196;
wire n_7487;
wire n_4585;
wire n_18273;
wire n_1785;
wire n_3406;
wire n_20445;
wire n_20414;
wire n_20109;
wire n_1381;
wire n_15406;
wire n_6268;
wire n_5604;
wire n_3470;
wire n_7663;
wire n_12308;
wire n_10846;
wire n_14854;
wire n_13024;
wire n_6529;
wire n_973;
wire n_4762;
wire n_3844;
wire n_11192;
wire n_20070;
wire n_11229;
wire n_4490;
wire n_8295;
wire n_1054;
wire n_7977;
wire n_15166;
wire n_14719;
wire n_5387;
wire n_11848;
wire n_7652;
wire n_4644;
wire n_8956;
wire n_8673;
wire n_14631;
wire n_4131;
wire n_11876;
wire n_16120;
wire n_12667;
wire n_18726;
wire n_15121;
wire n_2488;
wire n_828;
wire n_6134;
wire n_14824;
wire n_18602;
wire n_12878;
wire n_15886;
wire n_19697;
wire n_18048;
wire n_11666;
wire n_5325;
wire n_19429;
wire n_8960;
wire n_12361;
wire n_5004;
wire n_10233;
wire n_4926;
wire n_17988;
wire n_16734;
wire n_5876;
wire n_2550;
wire n_6160;
wire n_5813;
wire n_6235;
wire n_6212;
wire n_6816;
wire n_17950;
wire n_7374;
wire n_12753;
wire n_2291;
wire n_19317;
wire n_9549;
wire n_2165;
wire n_15402;
wire n_15539;
wire n_4210;
wire n_18469;
wire n_788;
wire n_18677;
wire n_18181;
wire n_15485;
wire n_13481;
wire n_17475;
wire n_12482;
wire n_8451;
wire n_6089;
wire n_16363;
wire n_11780;
wire n_5133;
wire n_14607;
wire n_7553;
wire n_5990;
wire n_1625;
wire n_318;
wire n_17853;
wire n_19767;
wire n_11467;
wire n_1412;
wire n_13351;
wire n_1922;
wire n_12997;
wire n_16169;
wire n_10625;
wire n_4877;
wire n_9312;
wire n_12818;
wire n_16572;
wire n_9151;
wire n_14576;
wire n_14981;
wire n_1904;
wire n_16541;
wire n_8830;
wire n_16994;
wire n_2395;
wire n_9324;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_14790;
wire n_8021;
wire n_11092;
wire n_1170;
wire n_9736;
wire n_7041;
wire n_19961;
wire n_6881;
wire n_18256;
wire n_15629;
wire n_16997;
wire n_9402;
wire n_13276;
wire n_7866;
wire n_7334;
wire n_3379;
wire n_4379;
wire n_16998;
wire n_18203;
wire n_8773;
wire n_5947;
wire n_8570;
wire n_16868;
wire n_1452;
wire n_10096;
wire n_668;
wire n_15333;
wire n_19163;
wire n_3743;
wire n_15762;
wire n_8079;
wire n_14106;
wire n_12560;
wire n_19704;
wire n_18190;
wire n_16077;
wire n_1003;
wire n_12477;
wire n_15422;
wire n_20258;
wire n_12523;
wire n_291;
wire n_16054;
wire n_10449;
wire n_14806;
wire n_8778;
wire n_5893;
wire n_20930;
wire n_11345;
wire n_15989;
wire n_16700;
wire n_17502;
wire n_17529;
wire n_2397;
wire n_19507;
wire n_6669;
wire n_17338;
wire n_17538;
wire n_1892;
wire n_6251;
wire n_1212;
wire n_14901;
wire n_4566;
wire n_4371;
wire n_12771;
wire n_10805;
wire n_7358;
wire n_8240;
wire n_7707;
wire n_18328;
wire n_2552;
wire n_9603;
wire n_8853;
wire n_19674;
wire n_5083;
wire n_15159;
wire n_20727;
wire n_14599;
wire n_11559;
wire n_7673;
wire n_15674;
wire n_11686;
wire n_18212;
wire n_7187;
wire n_12480;
wire n_10511;
wire n_20279;
wire n_9012;
wire n_5122;
wire n_11992;
wire n_18535;
wire n_17572;
wire n_2472;
wire n_13754;
wire n_10613;
wire n_6641;
wire n_3845;
wire n_3203;
wire n_13285;
wire n_383;
wire n_18758;
wire n_11814;
wire n_4298;
wire n_10594;
wire n_11622;
wire n_8445;
wire n_1781;
wire n_13413;
wire n_3690;
wire n_8464;
wire n_17668;
wire n_13608;
wire n_11952;
wire n_4211;
wire n_20647;
wire n_16424;
wire n_17666;
wire n_8376;
wire n_5032;
wire n_11506;
wire n_17275;
wire n_7071;
wire n_10797;
wire n_18526;
wire n_20077;
wire n_16695;
wire n_8848;
wire n_6288;
wire n_1862;
wire n_14573;
wire n_20143;
wire n_8894;
wire n_16118;
wire n_17511;
wire n_18452;
wire n_19878;
wire n_19671;
wire n_4128;
wire n_18230;
wire n_19925;
wire n_2955;
wire n_10784;
wire n_11035;
wire n_14009;
wire n_11174;
wire n_13759;
wire n_17201;
wire n_14911;
wire n_10234;
wire n_9230;
wire n_4101;
wire n_3866;
wire n_18816;
wire n_20654;
wire n_11705;
wire n_6409;
wire n_17006;
wire n_11003;
wire n_19128;
wire n_7657;
wire n_18254;
wire n_574;
wire n_17658;
wire n_15279;
wire n_6839;
wire n_9614;
wire n_8967;
wire n_16872;
wire n_1896;
wire n_21045;
wire n_17893;
wire n_8084;
wire n_8856;
wire n_12778;
wire n_12685;
wire n_18335;
wire n_10734;
wire n_20047;
wire n_6051;
wire n_19376;
wire n_8219;
wire n_5507;
wire n_15898;
wire n_10608;
wire n_195;
wire n_19664;
wire n_1328;
wire n_10746;
wire n_18838;
wire n_3519;
wire n_7504;
wire n_7099;
wire n_18889;
wire n_5642;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_14342;
wire n_9926;
wire n_1699;
wire n_8338;
wire n_1631;
wire n_12024;
wire n_18679;
wire n_156;
wire n_6566;
wire n_20505;
wire n_18343;
wire n_9462;
wire n_10900;
wire n_7998;
wire n_8666;
wire n_3053;
wire n_204;
wire n_11438;
wire n_18041;
wire n_14539;
wire n_10052;
wire n_3128;
wire n_18734;
wire n_13667;
wire n_4277;
wire n_16464;
wire n_4614;
wire n_1002;
wire n_11387;
wire n_18357;
wire n_13971;
wire n_15929;
wire n_11099;
wire n_12305;
wire n_7450;
wire n_6081;
wire n_13436;
wire n_20901;
wire n_329;
wire n_3821;
wire n_20786;
wire n_7780;
wire n_8523;
wire n_10476;
wire n_10559;
wire n_13797;
wire n_12439;
wire n_15522;
wire n_258;
wire n_13575;
wire n_7421;
wire n_16239;
wire n_19893;
wire n_2965;
wire n_12366;
wire n_11112;
wire n_14915;
wire n_10114;
wire n_1251;
wire n_18747;
wire n_1989;
wire n_2689;
wire n_10269;
wire n_6238;
wire n_18946;
wire n_8380;
wire n_13371;
wire n_17885;
wire n_16547;
wire n_1672;
wire n_16471;
wire n_4645;
wire n_17127;
wire n_20360;
wire n_18495;
wire n_3308;
wire n_6326;
wire n_19858;
wire n_17600;
wire n_2851;
wire n_17399;
wire n_4474;
wire n_20602;
wire n_10943;
wire n_10453;
wire n_15048;
wire n_7329;
wire n_13909;
wire n_7029;
wire n_18655;
wire n_4770;
wire n_14469;
wire n_5093;
wire n_18975;
wire n_4586;
wire n_19065;
wire n_15304;
wire n_14470;
wire n_3500;
wire n_6603;
wire n_5402;
wire n_11190;
wire n_13957;
wire n_2680;
wire n_16683;
wire n_3264;
wire n_10649;
wire n_2993;
wire n_20416;
wire n_2879;
wire n_15369;
wire n_11453;
wire n_416;
wire n_1430;
wire n_12806;
wire n_18112;
wire n_2729;
wire n_4302;
wire n_18851;
wire n_7127;
wire n_4547;
wire n_13718;
wire n_8321;
wire n_2376;
wire n_7805;
wire n_9807;
wire n_2790;
wire n_7542;
wire n_12354;
wire n_7053;
wire n_11614;
wire n_14807;
wire n_11143;
wire n_19183;
wire n_8037;
wire n_4610;
wire n_13029;
wire n_15093;
wire n_18878;
wire n_5263;
wire n_15293;
wire n_8997;
wire n_17843;
wire n_16698;
wire n_1682;
wire n_20005;
wire n_11349;
wire n_7001;
wire n_13875;
wire n_6129;
wire n_10574;
wire n_13066;
wire n_5590;
wire n_17844;
wire n_2621;
wire n_9286;
wire n_338;
wire n_15404;
wire n_10380;
wire n_13491;
wire n_9358;
wire n_1761;
wire n_16817;
wire n_1018;
wire n_7428;
wire n_12581;
wire n_17012;
wire n_16108;
wire n_8068;
wire n_2390;
wire n_6891;
wire n_20531;
wire n_625;
wire n_18153;
wire n_1107;
wire n_15750;
wire n_10528;
wire n_8097;
wire n_5481;
wire n_13120;
wire n_8114;
wire n_14572;
wire n_8126;
wire n_15441;
wire n_1241;
wire n_14378;
wire n_11736;
wire n_18267;
wire n_17964;
wire n_507;
wire n_9809;
wire n_14636;
wire n_3144;
wire n_9613;
wire n_17139;
wire n_4567;
wire n_17496;
wire n_9897;
wire n_11767;
wire n_6128;
wire n_11807;
wire n_3639;
wire n_11944;
wire n_3121;
wire n_11474;
wire n_3015;
wire n_3870;
wire n_1085;
wire n_19177;
wire n_11692;
wire n_1900;
wire n_620;
wire n_6096;
wire n_19535;
wire n_863;
wire n_6992;
wire n_303;
wire n_12863;
wire n_2433;
wire n_5830;
wire n_1495;
wire n_6681;
wire n_4227;
wire n_11737;
wire n_533;
wire n_15326;
wire n_2456;
wire n_20715;
wire n_13466;
wire n_13689;
wire n_14115;
wire n_17917;
wire n_20821;
wire n_12792;
wire n_19359;
wire n_844;
wire n_8176;
wire n_7215;
wire n_7441;
wire n_20761;
wire n_2382;
wire n_237;
wire n_780;
wire n_1918;
wire n_8327;
wire n_4119;
wire n_9811;
wire n_1140;
wire n_5843;
wire n_15702;
wire n_8539;
wire n_15566;
wire n_11068;
wire n_17144;
wire n_18042;
wire n_3012;
wire n_13768;
wire n_3850;
wire n_11476;
wire n_21011;
wire n_19861;
wire n_13111;
wire n_1216;
wire n_11957;
wire n_8204;
wire n_19661;
wire n_9199;
wire n_12155;
wire n_15221;
wire n_11210;
wire n_7162;
wire n_17315;
wire n_9808;
wire n_18069;
wire n_8958;
wire n_11333;
wire n_1432;
wire n_13692;
wire n_16483;
wire n_18409;
wire n_13126;
wire n_851;
wire n_10579;
wire n_3900;
wire n_10707;
wire n_15682;
wire n_17363;
wire n_9265;
wire n_12332;
wire n_18949;
wire n_11352;
wire n_3862;
wire n_12641;
wire n_930;
wire n_10556;
wire n_8572;
wire n_17548;
wire n_19546;
wire n_8424;
wire n_20929;
wire n_8147;
wire n_4993;
wire n_16950;
wire n_3678;
wire n_10080;
wire n_20902;
wire n_3549;
wire n_3914;
wire n_10766;
wire n_6398;
wire n_11222;
wire n_7461;
wire n_17186;
wire n_1692;
wire n_20487;
wire n_11650;
wire n_14310;
wire n_2611;
wire n_18776;
wire n_15690;
wire n_13531;
wire n_4745;
wire n_14215;
wire n_6319;
wire n_20964;
wire n_10217;
wire n_6966;
wire n_9791;
wire n_9449;
wire n_9149;
wire n_9686;
wire n_19121;
wire n_19462;
wire n_7838;
wire n_9844;
wire n_6724;
wire n_17401;
wire n_6776;
wire n_9458;
wire n_15994;
wire n_20783;
wire n_8455;
wire n_2087;
wire n_9128;
wire n_746;
wire n_292;
wire n_12816;
wire n_14730;
wire n_6710;
wire n_1787;
wire n_18355;
wire n_3172;
wire n_16076;
wire n_2659;
wire n_4033;
wire n_20752;
wire n_10446;
wire n_15010;
wire n_6553;
wire n_10219;
wire n_4508;
wire n_16803;
wire n_3614;
wire n_19983;
wire n_20536;
wire n_4141;
wire n_13877;
wire n_20453;
wire n_6893;
wire n_12377;
wire n_12007;
wire n_5179;
wire n_15240;
wire n_5685;
wire n_14032;
wire n_14822;
wire n_9094;
wire n_19054;
wire n_13524;
wire n_14075;
wire n_4364;
wire n_11049;
wire n_9510;
wire n_20810;
wire n_14817;
wire n_12319;
wire n_14178;
wire n_1841;
wire n_16138;
wire n_12388;
wire n_6206;
wire n_18967;
wire n_7893;
wire n_2954;
wire n_9429;
wire n_489;
wire n_11599;
wire n_15740;
wire n_18997;
wire n_251;
wire n_974;
wire n_4367;
wire n_5134;
wire n_4866;
wire n_18483;
wire n_8123;
wire n_16080;
wire n_14472;
wire n_17015;
wire n_13659;
wire n_307;
wire n_14946;
wire n_13473;
wire n_16815;
wire n_12165;
wire n_16262;
wire n_13497;
wire n_9661;
wire n_9799;
wire n_18665;
wire n_5373;
wire n_7403;
wire n_17553;
wire n_18521;
wire n_3320;
wire n_16975;
wire n_2144;
wire n_6033;
wire n_1247;
wire n_19949;
wire n_10364;
wire n_6060;
wire n_15734;
wire n_9895;
wire n_10288;
wire n_6709;
wire n_11602;
wire n_13843;
wire n_11865;
wire n_15263;
wire n_18577;
wire n_2980;
wire n_1728;
wire n_3311;
wire n_18415;
wire n_11613;
wire n_18540;
wire n_18804;
wire n_7221;
wire n_11870;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_3704;
wire n_8423;
wire n_670;
wire n_379;
wire n_16539;
wire n_20976;
wire n_19817;
wire n_5088;
wire n_441;
wire n_12123;
wire n_18455;
wire n_5392;
wire n_1743;
wire n_8548;
wire n_207;
wire n_15774;
wire n_13738;
wire n_7185;
wire n_17905;
wire n_10889;
wire n_17687;
wire n_6234;
wire n_4153;
wire n_15459;
wire n_5089;
wire n_11394;
wire n_20390;
wire n_16630;
wire n_18792;
wire n_3759;
wire n_9964;
wire n_16870;
wire n_9719;
wire n_16822;
wire n_2617;
wire n_6619;
wire n_13200;
wire n_19619;
wire n_13876;
wire n_19859;
wire n_18601;
wire n_7233;
wire n_17985;
wire n_2122;
wire n_4543;
wire n_11186;
wire n_12996;
wire n_2067;
wire n_8402;
wire n_14097;
wire n_20384;
wire n_15125;
wire n_19775;
wire n_5398;
wire n_20282;
wire n_2194;
wire n_4640;
wire n_16688;
wire n_7202;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_8595;
wire n_11181;
wire n_9040;
wire n_10817;
wire n_12277;
wire n_12062;
wire n_13386;
wire n_16405;
wire n_18600;
wire n_17776;
wire n_15844;
wire n_19103;
wire n_707;
wire n_5051;
wire n_10132;
wire n_2783;
wire n_8520;
wire n_18472;
wire n_9456;
wire n_6366;
wire n_1015;
wire n_6304;
wire n_13605;
wire n_7547;
wire n_5552;
wire n_6074;
wire n_15083;
wire n_15257;
wire n_11286;
wire n_8030;
wire n_16671;
wire n_14511;
wire n_9219;
wire n_17676;
wire n_19500;
wire n_5242;
wire n_1188;
wire n_7527;
wire n_15776;
wire n_7948;
wire n_2618;
wire n_20974;
wire n_7096;
wire n_11863;
wire n_9206;
wire n_19492;
wire n_8485;
wire n_15847;
wire n_3781;
wire n_17031;
wire n_11225;
wire n_20698;
wire n_5127;
wire n_15239;
wire n_4313;
wire n_13113;
wire n_4670;
wire n_3713;
wire n_1863;
wire n_5536;
wire n_15928;
wire n_7293;
wire n_11862;
wire n_4297;
wire n_5810;
wire n_3356;
wire n_20434;
wire n_2190;
wire n_4991;
wire n_13360;
wire n_17735;
wire n_3070;
wire n_15065;
wire n_13044;
wire n_3245;
wire n_12859;
wire n_16025;
wire n_2894;
wire n_9559;
wire n_9709;
wire n_2452;
wire n_8626;
wire n_17294;
wire n_13217;
wire n_10810;
wire n_17656;
wire n_20224;
wire n_8166;
wire n_9356;
wire n_4252;
wire n_5009;
wire n_15689;
wire n_16532;
wire n_20353;
wire n_16833;
wire n_18533;
wire n_12846;
wire n_15467;
wire n_15346;
wire n_7762;
wire n_13840;
wire n_11501;
wire n_17182;
wire n_4446;
wire n_9342;
wire n_19796;
wire n_18053;
wire n_12234;
wire n_1797;
wire n_4425;
wire n_15863;
wire n_744;
wire n_7936;
wire n_215;
wire n_13117;
wire n_1331;
wire n_12042;
wire n_6031;
wire n_16084;
wire n_4237;
wire n_5297;
wire n_20421;
wire n_4828;
wire n_15138;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_10622;
wire n_20566;
wire n_1580;
wire n_2448;
wire n_11639;
wire n_2211;
wire n_8955;
wire n_17888;
wire n_9551;
wire n_5904;
wire n_19039;
wire n_4697;
wire n_16069;
wire n_13230;
wire n_3277;
wire n_10880;
wire n_14612;
wire n_5463;
wire n_18172;
wire n_18049;
wire n_8628;
wire n_13559;
wire n_15400;
wire n_20514;
wire n_15723;
wire n_7481;
wire n_11447;
wire n_6484;
wire n_3340;
wire n_14517;
wire n_5483;
wire n_12534;
wire n_9539;
wire n_8617;
wire n_14297;
wire n_9268;
wire n_9718;
wire n_6639;
wire n_11258;
wire n_358;
wire n_11168;
wire n_18433;
wire n_12148;
wire n_12142;
wire n_9527;
wire n_19568;
wire n_3256;
wire n_15115;
wire n_16269;
wire n_7689;
wire n_19189;
wire n_9952;
wire n_11612;
wire n_20173;
wire n_13782;
wire n_2520;
wire n_13612;
wire n_7010;
wire n_9798;
wire n_20139;
wire n_20079;
wire n_1025;
wire n_17162;
wire n_10537;
wire n_14684;
wire n_19801;
wire n_20827;
wire n_687;
wire n_480;
wire n_13920;
wire n_6555;
wire n_16495;
wire n_4306;
wire n_13130;
wire n_4006;
wire n_12812;
wire n_3102;
wire n_1499;
wire n_4098;
wire n_9635;
wire n_15542;
wire n_19849;
wire n_17284;
wire n_4972;
wire n_1476;
wire n_6036;
wire n_9405;
wire n_16561;
wire n_15255;
wire n_3925;
wire n_17991;
wire n_11481;
wire n_651;
wire n_2850;
wire n_12057;
wire n_12050;
wire n_9726;
wire n_11774;
wire n_14357;
wire n_9540;
wire n_13972;
wire n_13767;
wire n_7824;
wire n_18992;
wire n_3843;
wire n_16909;
wire n_19698;
wire n_4805;
wire n_19781;
wire n_15838;
wire n_10675;
wire n_2386;
wire n_19751;
wire n_9626;
wire n_4822;
wire n_11327;
wire n_6946;
wire n_7947;
wire n_18192;
wire n_4635;
wire n_1450;
wire n_12824;
wire n_12392;
wire n_14545;
wire n_3740;
wire n_1815;
wire n_16858;
wire n_7039;
wire n_8027;
wire n_17974;
wire n_17962;
wire n_14677;
wire n_8406;
wire n_5994;
wire n_14037;
wire n_11265;
wire n_19306;
wire n_9754;
wire n_17802;
wire n_8849;
wire n_13071;
wire n_14127;
wire n_11901;
wire n_3345;
wire n_12848;
wire n_10307;
wire n_4906;
wire n_11754;
wire n_13825;
wire n_6840;
wire n_8535;
wire n_8348;
wire n_6915;
wire n_17825;
wire n_12320;
wire n_20532;
wire n_18548;
wire n_11413;
wire n_13953;
wire n_13040;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_19431;
wire n_10367;
wire n_833;
wire n_14602;
wire n_17035;
wire n_8294;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_20347;
wire n_2413;
wire n_13765;
wire n_18798;
wire n_2605;
wire n_7887;
wire n_9298;
wire n_5884;
wire n_4882;
wire n_10006;
wire n_5728;
wire n_1035;
wire n_13334;
wire n_3475;
wire n_14902;
wire n_18867;
wire n_14450;
wire n_2044;
wire n_15633;
wire n_3886;
wire n_732;
wire n_7521;
wire n_20650;
wire n_16933;
wire n_15110;
wire n_9943;
wire n_7569;
wire n_13745;
wire n_10966;
wire n_14697;
wire n_2968;
wire n_1882;
wire n_13646;
wire n_12130;
wire n_15049;
wire n_13031;
wire n_17819;
wire n_467;
wire n_17902;
wire n_2177;
wire n_18536;
wire n_16884;
wire n_6516;
wire n_14567;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7411;
wire n_13314;
wire n_7326;
wire n_21032;
wire n_14277;
wire n_19689;
wire n_19742;
wire n_16524;
wire n_8005;
wire n_5105;
wire n_3920;
wire n_20239;
wire n_15446;
wire n_5879;
wire n_11303;
wire n_5027;
wire n_775;
wire n_16995;
wire n_5688;
wire n_9030;
wire n_11216;
wire n_15652;
wire n_13638;
wire n_6630;
wire n_5759;
wire n_10409;
wire n_4631;
wire n_18124;
wire n_5999;
wire n_2110;
wire n_11346;
wire n_12530;
wire n_3822;
wire n_18379;
wire n_16199;
wire n_17604;
wire n_16129;
wire n_15575;
wire n_9583;
wire n_10349;
wire n_17303;
wire n_13035;
wire n_10636;
wire n_6403;
wire n_17196;
wire n_9862;
wire n_5451;
wire n_6578;
wire n_5460;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_11165;
wire n_3595;
wire n_6875;
wire n_9617;
wire n_18036;
wire n_18998;
wire n_941;
wire n_9749;
wire n_5517;
wire n_13654;
wire n_19457;
wire n_20057;
wire n_19283;
wire n_19960;
wire n_18716;
wire n_5695;
wire n_18199;
wire n_1940;
wire n_3683;
wire n_11410;
wire n_18672;
wire n_4452;
wire n_284;
wire n_3887;
wire n_5587;
wire n_10845;
wire n_18158;
wire n_15630;
wire n_8907;
wire n_2963;
wire n_5674;
wire n_7499;
wire n_9423;
wire n_526;
wire n_19840;
wire n_674;
wire n_4079;
wire n_1749;
wire n_15227;
wire n_1653;
wire n_10063;
wire n_6559;
wire n_4088;
wire n_8777;
wire n_11149;
wire n_2669;
wire n_6068;
wire n_12236;
wire n_18855;
wire n_4366;
wire n_18565;
wire n_13554;
wire n_6080;
wire n_14372;
wire n_13421;
wire n_7927;
wire n_20462;
wire n_2688;
wire n_6150;
wire n_13795;
wire n_14989;
wire n_1910;
wire n_16792;
wire n_19290;
wire n_20401;
wire n_2018;
wire n_2672;
wire n_5780;
wire n_3433;
wire n_3597;
wire n_13864;
wire n_5743;
wire n_1956;
wire n_12273;
wire n_15809;
wire n_6022;
wire n_2828;
wire n_16320;
wire n_14331;
wire n_19366;
wire n_7691;
wire n_296;
wire n_7745;
wire n_17509;
wire n_3645;
wire n_5705;
wire n_7335;
wire n_12400;
wire n_17099;
wire n_10472;
wire n_19986;
wire n_16718;
wire n_6116;
wire n_18060;
wire n_8780;
wire n_16867;
wire n_1805;
wire n_19199;
wire n_15736;
wire n_16036;
wire n_6757;
wire n_10218;
wire n_5875;
wire n_18388;
wire n_3714;
wire n_9093;
wire n_184;
wire n_15200;
wire n_20156;
wire n_19906;
wire n_12950;
wire n_3676;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_3125;
wire n_12250;
wire n_19962;
wire n_14792;
wire n_5618;
wire n_15760;
wire n_12904;
wire n_6495;
wire n_14669;
wire n_12444;
wire n_11163;
wire n_9425;
wire n_13373;
wire n_20800;
wire n_11730;
wire n_11916;
wire n_3502;
wire n_11311;
wire n_14525;
wire n_14435;
wire n_7993;
wire n_11151;
wire n_1008;
wire n_13153;
wire n_15195;
wire n_581;
wire n_13091;
wire n_12079;
wire n_4628;
wire n_7343;
wire n_21064;
wire n_5982;
wire n_16548;
wire n_13306;
wire n_9344;
wire n_14657;
wire n_7109;
wire n_16082;
wire n_19599;
wire n_12125;
wire n_341;
wire n_1270;
wire n_549;
wire n_6155;
wire n_18107;
wire n_2901;
wire n_17546;
wire n_15165;
wire n_8530;
wire n_15434;
wire n_3621;
wire n_5529;
wire n_6349;
wire n_8500;
wire n_8713;
wire n_14554;
wire n_8297;
wire n_8926;
wire n_14974;
wire n_18489;
wire n_8025;
wire n_5354;
wire n_15498;
wire n_7898;
wire n_11357;
wire n_11027;
wire n_1788;
wire n_20600;
wire n_18330;
wire n_17097;
wire n_7070;
wire n_20659;
wire n_5276;
wire n_11160;
wire n_13043;
wire n_3804;
wire n_3211;
wire n_18020;
wire n_2440;
wire n_2096;
wire n_14892;
wire n_2215;
wire n_13468;
wire n_15830;
wire n_4073;
wire n_8880;
wire n_20395;
wire n_16675;
wire n_13831;
wire n_16105;
wire n_4001;
wire n_8471;
wire n_14529;
wire n_15940;
wire n_18219;
wire n_12906;
wire n_12490;
wire n_6273;
wire n_14424;
wire n_7094;
wire n_20562;
wire n_3111;
wire n_12751;
wire n_10640;
wire n_1813;
wire n_315;
wire n_11897;
wire n_1573;
wire n_19489;
wire n_758;
wire n_10272;
wire n_15070;
wire n_5907;
wire n_784;
wire n_4339;
wire n_19403;
wire n_6182;
wire n_6754;
wire n_14916;
wire n_1076;
wire n_1348;
wire n_12242;
wire n_2445;
wire n_4023;
wire n_3632;
wire n_20905;
wire n_309;
wire n_16241;
wire n_16296;
wire n_5478;
wire n_13382;
wire n_10176;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_17498;
wire n_17316;
wire n_21087;
wire n_9061;
wire n_18143;
wire n_7995;
wire n_17515;
wire n_10254;
wire n_1991;
wire n_14955;
wire n_10332;
wire n_16117;
wire n_17289;
wire n_614;
wire n_12173;
wire n_10257;
wire n_9668;
wire n_17056;
wire n_6592;
wire n_16626;
wire n_2541;
wire n_10195;
wire n_1113;
wire n_1615;
wire n_2372;
wire n_2105;
wire n_20177;
wire n_1806;
wire n_8803;
wire n_10866;
wire n_1673;
wire n_17298;
wire n_4473;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_19515;
wire n_18399;
wire n_3018;
wire n_8818;
wire n_16525;
wire n_20446;
wire n_6962;
wire n_16800;
wire n_18135;
wire n_14716;
wire n_5040;
wire n_18225;
wire n_15384;
wire n_4695;
wire n_15362;
wire n_12542;
wire n_16040;
wire n_15187;
wire n_458;
wire n_11499;
wire n_3628;
wire n_14390;
wire n_20180;
wire n_9433;
wire n_11746;
wire n_658;
wire n_362;
wire n_16526;
wire n_10430;
wire n_12934;
wire n_18310;
wire n_18127;
wire n_19565;
wire n_13941;
wire n_15805;
wire n_3872;
wire n_16449;
wire n_14694;
wire n_1777;
wire n_9552;
wire n_7395;
wire n_20370;
wire n_15888;
wire n_20911;
wire n_3441;
wire n_19902;
wire n_4146;
wire n_15795;
wire n_6609;
wire n_7635;
wire n_2115;
wire n_8567;
wire n_18244;
wire n_10667;
wire n_1347;
wire n_18037;
wire n_18157;
wire n_3534;
wire n_450;
wire n_8578;
wire n_2670;
wire n_13975;
wire n_896;
wire n_15624;
wire n_20435;
wire n_4557;
wire n_20217;
wire n_20118;
wire n_17467;
wire n_1337;
wire n_2148;
wire n_7788;
wire n_16903;
wire n_17688;
wire n_4663;
wire n_15718;
wire n_18738;
wire n_16024;
wire n_5136;
wire n_12303;
wire n_1705;
wire n_3149;
wire n_18493;
wire n_14844;
wire n_12597;
wire n_9757;
wire n_11886;
wire n_19223;
wire n_8761;
wire n_14316;
wire n_7630;
wire n_17049;
wire n_18337;
wire n_1581;
wire n_3058;
wire n_5355;
wire n_13706;
wire n_375;
wire n_998;
wire n_12039;
wire n_10663;
wire n_17880;
wire n_20000;
wire n_20269;
wire n_11792;
wire n_17486;
wire n_16059;
wire n_18901;
wire n_1368;
wire n_3722;
wire n_15412;
wire n_1339;
wire n_14356;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_19644;
wire n_15535;
wire n_7541;
wire n_7913;
wire n_13890;
wire n_11965;
wire n_15158;
wire n_5669;
wire n_3334;
wire n_14852;
wire n_15006;
wire n_18325;
wire n_8875;
wire n_5515;
wire n_11588;
wire n_18364;
wire n_11592;
wire n_3083;
wire n_12290;
wire n_9801;
wire n_12718;
wire n_8649;
wire n_2259;
wire n_11235;
wire n_5059;
wire n_9424;
wire n_9333;
wire n_18185;
wire n_18896;
wire n_11673;
wire n_1233;
wire n_4493;
wire n_17812;
wire n_17816;
wire n_7161;
wire n_9004;
wire n_6364;
wire n_15663;
wire n_16920;
wire n_6848;
wire n_2479;
wire n_886;
wire n_13548;
wire n_16810;
wire n_675;
wire n_9200;
wire n_15035;
wire n_7806;
wire n_3432;
wire n_11059;
wire n_14047;
wire n_16200;
wire n_3480;
wire n_7676;
wire n_11683;
wire n_5467;
wire n_7241;
wire n_15612;
wire n_1169;
wire n_789;
wire n_19896;
wire n_9207;
wire n_13592;
wire n_1916;
wire n_10356;
wire n_12717;
wire n_7644;
wire n_9276;
wire n_14186;
wire n_8829;
wire n_2818;
wire n_18871;
wire n_17038;
wire n_20882;
wire n_18227;
wire n_14540;
wire n_3668;
wire n_1515;
wire n_817;
wire n_14272;
wire n_13260;
wire n_11718;
wire n_2671;
wire n_18266;
wire n_19519;
wire n_17197;
wire n_19161;
wire n_9728;
wire n_4103;
wire n_18021;
wire n_8101;
wire n_13712;
wire n_15549;
wire n_17256;
wire n_1366;
wire n_8749;
wire n_13349;
wire n_8937;
wire n_13233;
wire n_7067;
wire n_12087;
wire n_16323;
wire n_4416;
wire n_15555;
wire n_10998;
wire n_12936;
wire n_13300;
wire n_16461;
wire n_11743;
wire n_12765;
wire n_3930;
wire n_17412;
wire n_9610;
wire n_5471;
wire n_3081;
wire n_10756;
wire n_5497;
wire n_9139;
wire n_5519;
wire n_1961;
wire n_3270;
wire n_15236;
wire n_17153;
wire n_4814;
wire n_8801;
wire n_17203;
wire n_18439;
wire n_15983;
wire n_20484;
wire n_11879;
wire n_13900;
wire n_10782;
wire n_12386;
wire n_13679;
wire n_6862;
wire n_11842;
wire n_20805;
wire n_12746;
wire n_14023;
wire n_20069;
wire n_11320;
wire n_15728;
wire n_645;
wire n_17252;
wire n_10251;
wire n_16658;
wire n_15253;
wire n_721;
wire n_18000;
wire n_1276;
wire n_21088;
wire n_10737;
wire n_10475;
wire n_3252;
wire n_6647;
wire n_18743;
wire n_8040;
wire n_6941;
wire n_7239;
wire n_16523;
wire n_7826;
wire n_9981;
wire n_8102;
wire n_10541;
wire n_11419;
wire n_11171;
wire n_3859;
wire n_5592;
wire n_3150;
wire n_5491;
wire n_9825;
wire n_19349;
wire n_15315;
wire n_17029;
wire n_16623;
wire n_1034;
wire n_1652;
wire n_7078;
wire n_12352;
wire n_18531;
wire n_11459;
wire n_9043;
wire n_11998;
wire n_8269;
wire n_7006;
wire n_4031;
wire n_3571;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_17121;
wire n_14706;
wire n_11662;
wire n_16013;
wire n_4340;
wire n_7812;
wire n_9766;
wire n_6778;
wire n_11877;
wire n_5526;
wire n_5202;
wire n_12074;
wire n_15819;
wire n_3817;
wire n_17709;
wire n_612;
wire n_333;
wire n_7165;
wire n_9777;
wire n_20596;
wire n_20729;
wire n_6830;
wire n_2061;
wire n_2685;
wire n_16737;
wire n_12252;
wire n_17694;
wire n_9666;
wire n_10028;
wire n_15842;
wire n_11532;
wire n_12868;
wire n_1391;
wire n_9605;
wire n_17310;
wire n_1006;
wire n_16033;
wire n_14755;
wire n_4995;
wire n_5873;
wire n_6514;
wire n_17200;
wire n_10083;
wire n_1245;
wire n_16592;
wire n_3429;
wire n_3758;
wire n_2326;
wire n_4109;
wire n_11494;
wire n_1872;
wire n_14090;
wire n_5926;
wire n_16226;
wire n_14347;
wire n_9724;
wire n_652;
wire n_8403;
wire n_20386;
wire n_18154;
wire n_3716;
wire n_11570;
wire n_15945;
wire n_2926;
wire n_798;
wire n_13631;
wire n_16820;
wire n_7781;
wire n_14746;
wire n_10295;
wire n_8296;
wire n_6429;
wire n_4235;
wire n_21067;
wire n_18125;
wire n_11122;
wire n_6775;
wire n_2185;
wire n_20561;
wire n_4345;
wire n_17216;
wire n_9205;
wire n_9418;
wire n_17304;
wire n_12205;
wire n_8676;
wire n_15119;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_10341;
wire n_12606;
wire n_5812;
wire n_15008;
wire n_9973;
wire n_20975;
wire n_5804;
wire n_3240;
wire n_14253;
wire n_16520;
wire n_3362;
wire n_4130;
wire n_14212;
wire n_9020;
wire n_9619;
wire n_10161;
wire n_13003;
wire n_8652;
wire n_16708;
wire n_20132;
wire n_12843;
wire n_4456;
wire n_9691;
wire n_2365;
wire n_9133;
wire n_1399;
wire n_5981;
wire n_20311;
wire n_7784;
wire n_16965;
wire n_19017;
wire n_10902;
wire n_15477;
wire n_17351;
wire n_4020;
wire n_17997;
wire n_19148;
wire n_6933;
wire n_1970;
wire n_17623;
wire n_3724;
wire n_9353;
wire n_20961;
wire n_4055;
wire n_5444;
wire n_11590;
wire n_5737;
wire n_8439;
wire n_6908;
wire n_5615;
wire n_17157;
wire n_10323;
wire n_6083;
wire n_8499;
wire n_767;
wire n_13322;
wire n_8772;
wire n_19117;
wire n_6278;
wire n_11430;
wire n_7195;
wire n_15072;
wire n_18159;
wire n_3342;
wire n_6101;
wire n_20829;
wire n_3796;
wire n_16488;
wire n_3884;
wire n_13850;
wire n_16411;
wire n_13835;
wire n_5550;
wire n_3375;
wire n_15224;
wire n_20094;
wire n_155;
wire n_15029;
wire n_2363;
wire n_12687;
wire n_14460;
wire n_19594;
wire n_15640;
wire n_17863;
wire n_7115;
wire n_17123;
wire n_1020;
wire n_16216;
wire n_15382;
wire n_12022;
wire n_172;
wire n_11535;
wire n_12624;
wire n_11808;
wire n_8789;
wire n_7520;
wire n_1279;
wire n_9377;
wire n_2511;
wire n_9224;
wire n_11577;
wire n_15045;
wire n_17253;
wire n_16577;
wire n_16802;
wire n_19687;
wire n_20750;
wire n_7222;
wire n_8678;
wire n_12981;
wire n_1255;
wire n_20202;
wire n_2335;
wire n_10289;
wire n_9145;
wire n_12716;
wire n_13079;
wire n_15130;
wire n_1401;
wire n_8901;
wire n_4494;
wire n_9887;
wire n_7206;
wire n_8869;
wire n_552;
wire n_11729;
wire n_14012;
wire n_8272;
wire n_3577;
wire n_6625;
wire n_4636;
wire n_16764;
wire n_6826;
wire n_11727;
wire n_327;
wire n_6341;
wire n_4386;
wire n_10183;
wire n_13693;
wire n_8870;
wire n_5041;
wire n_11433;
wire n_8178;
wire n_5524;
wire n_926;
wire n_13434;
wire n_8234;
wire n_17605;
wire n_2178;
wire n_2765;
wire n_12759;
wire n_14418;
wire n_186;
wire n_17741;
wire n_11840;
wire n_2241;
wire n_9774;
wire n_2531;
wire n_11987;
wire n_11052;
wire n_3377;
wire n_18420;
wire n_1518;
wire n_13476;
wire n_14803;
wire n_11169;
wire n_855;
wire n_20630;
wire n_8862;
wire n_13229;
wire n_2059;
wire n_14092;
wire n_8184;
wire n_13950;
wire n_6911;
wire n_14219;
wire n_13344;
wire n_19015;
wire n_18106;
wire n_10353;
wire n_10151;
wire n_12138;
wire n_3374;
wire n_7776;
wire n_8001;
wire n_12521;
wire n_11931;
wire n_11036;
wire n_8064;
wire n_14117;
wire n_13721;
wire n_15295;
wire n_6095;
wire n_4323;
wire n_13535;
wire n_5376;
wire n_13704;
wire n_18719;
wire n_5488;
wire n_9099;
wire n_1105;
wire n_10034;
wire n_11336;
wire n_18167;
wire n_8787;
wire n_9543;
wire n_8131;
wire n_19126;
wire n_19788;
wire n_14633;
wire n_16264;
wire n_14538;
wire n_7448;
wire n_4480;
wire n_6787;
wire n_20102;
wire n_17608;
wire n_16230;
wire n_6423;
wire n_8150;
wire n_5891;
wire n_9168;
wire n_2418;
wire n_1377;
wire n_18365;
wire n_12159;
wire n_20479;
wire n_3222;
wire n_325;
wire n_1740;
wire n_12259;
wire n_11665;
wire n_9367;
wire n_13402;
wire n_11685;
wire n_20940;
wire n_15662;
wire n_16923;
wire n_11801;
wire n_10230;
wire n_12117;
wire n_17938;
wire n_11573;
wire n_4374;
wire n_6176;
wire n_14395;
wire n_1408;
wire n_15042;
wire n_1693;
wire n_20520;
wire n_6969;
wire n_13060;
wire n_15651;
wire n_9496;
wire n_15214;
wire n_8914;
wire n_14082;
wire n_8821;
wire n_17380;
wire n_11446;
wire n_17064;
wire n_13586;
wire n_15163;
wire n_12772;
wire n_15979;
wire n_5362;
wire n_8209;
wire n_388;
wire n_18810;
wire n_4580;
wire n_15867;
wire n_17263;
wire n_21117;
wire n_18687;
wire n_20609;
wire n_21034;
wire n_12145;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_8963;
wire n_9191;
wire n_16177;
wire n_16617;
wire n_8550;
wire n_7449;
wire n_17009;
wire n_1502;
wire n_3501;
wire n_12889;
wire n_15793;
wire n_19769;
wire n_13096;
wire n_16857;
wire n_3216;
wire n_9913;
wire n_11626;
wire n_11178;
wire n_13684;
wire n_4844;
wire n_9329;
wire n_12608;
wire n_17740;
wire n_2661;
wire n_13008;
wire n_1649;
wire n_13742;
wire n_1297;
wire n_9627;
wire n_10271;
wire n_18586;
wire n_11295;
wire n_5729;
wire n_4677;
wire n_4525;
wire n_17944;
wire n_10402;
wire n_3364;
wire n_2643;
wire n_755;
wire n_9585;
wire n_15232;
wire n_17151;
wire n_1898;
wire n_8797;
wire n_21057;
wire n_11126;
wire n_3671;
wire n_9606;
wire n_15768;
wire n_19013;
wire n_476;
wire n_12026;
wire n_20576;
wire n_4104;
wire n_10047;
wire n_982;
wire n_20994;
wire n_3064;
wire n_13977;
wire n_16980;
wire n_3199;
wire n_11396;
wire n_7050;
wire n_7590;
wire n_17361;
wire n_403;
wire n_3016;
wire n_6739;
wire n_17297;
wire n_1319;
wire n_3669;
wire n_2480;
wire n_14869;
wire n_1700;
wire n_1332;
wire n_5385;
wire n_10523;
wire n_10377;
wire n_17562;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3459;
wire n_15013;
wire n_17343;
wire n_14739;
wire n_13724;
wire n_17030;
wire n_1966;
wire n_9708;
wire n_9130;
wire n_9988;
wire n_1513;
wire n_20397;
wire n_4524;
wire n_15374;
wire n_10173;
wire n_4657;
wire n_12075;
wire n_15478;
wire n_8837;
wire n_10999;
wire n_17451;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_8784;
wire n_20820;
wire n_3964;
wire n_20839;
wire n_15415;
wire n_8768;
wire n_8086;
wire n_20014;
wire n_16485;
wire n_16447;
wire n_9010;
wire n_11637;
wire n_2492;
wire n_12183;
wire n_13432;
wire n_20240;
wire n_4876;
wire n_15217;
wire n_241;
wire n_19791;
wire n_12519;
wire n_2900;
wire n_12955;
wire n_8307;
wire n_15290;
wire n_2622;
wire n_3447;
wire n_19709;
wire n_13214;
wire n_10412;
wire n_1950;
wire n_5928;
wire n_7830;
wire n_16642;
wire n_2249;
wire n_19048;
wire n_3463;
wire n_15399;
wire n_2785;
wire n_730;
wire n_1524;
wire n_19727;
wire n_469;
wire n_5504;
wire n_9345;
wire n_19069;
wire n_11820;
wire n_19591;
wire n_4239;
wire n_10509;
wire n_8010;
wire n_17539;
wire n_18718;
wire n_18367;
wire n_20583;
wire n_8950;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_9487;
wire n_18303;
wire n_13588;
wire n_5494;
wire n_12413;
wire n_17547;
wire n_18725;
wire n_7935;
wire n_2416;
wire n_17086;
wire n_12726;
wire n_12784;
wire n_20437;
wire n_9851;
wire n_15281;
wire n_4706;
wire n_3879;
wire n_6850;
wire n_12761;
wire n_4764;
wire n_2408;
wire n_13899;
wire n_17704;
wire n_4990;
wire n_11370;
wire n_19997;
wire n_949;
wire n_16266;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_2760;
wire n_4919;
wire n_15145;
wire n_15448;
wire n_8049;
wire n_13666;
wire n_7266;
wire n_1151;
wire n_20813;
wire n_19176;
wire n_4251;
wire n_2393;
wire n_18079;
wire n_3566;
wire n_5800;
wire n_17622;
wire n_19018;
wire n_15155;
wire n_4173;
wire n_5309;
wire n_15501;
wire n_19543;
wire n_16856;
wire n_19723;
wire n_12160;
wire n_2230;
wire n_9824;
wire n_14582;
wire n_7442;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_14508;
wire n_3783;
wire n_19701;
wire n_11654;
wire n_15208;
wire n_14562;
wire n_3643;
wire n_8681;
wire n_20308;
wire n_19753;
wire n_9884;
wire n_15972;
wire n_6026;
wire n_1143;
wire n_15453;
wire n_16484;
wire n_17384;
wire n_7136;
wire n_19799;
wire n_4960;
wire n_9693;
wire n_11546;
wire n_1153;
wire n_9273;
wire n_894;
wire n_1380;
wire n_20135;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_18104;
wire n_19717;
wire n_1023;
wire n_10932;
wire n_4327;
wire n_14799;
wire n_3190;
wire n_11697;
wire n_3695;
wire n_13555;
wire n_17018;
wire n_10487;
wire n_14853;
wire n_2820;
wire n_21082;
wire n_12512;
wire n_15043;
wire n_11937;
wire n_16596;
wire n_638;
wire n_4370;
wire n_17390;
wire n_19141;
wire n_5638;
wire n_16881;
wire n_5058;
wire n_13558;
wire n_9075;
wire n_13954;
wire n_2777;
wire n_11763;
wire n_7167;
wire n_5849;
wire n_3233;
wire n_8906;
wire n_1603;
wire n_7146;
wire n_4478;
wire n_18849;
wire n_2935;
wire n_4246;
wire n_14625;
wire n_7618;
wire n_2863;
wire n_19426;
wire n_4632;
wire n_16372;
wire n_11941;
wire n_12031;
wire n_20772;
wire n_11704;
wire n_2920;
wire n_9582;
wire n_8268;
wire n_17067;
wire n_15291;
wire n_20410;
wire n_1290;
wire n_4375;
wire n_15244;
wire n_617;
wire n_14340;
wire n_13743;
wire n_20190;
wire n_3368;
wire n_13951;
wire n_8008;
wire n_19409;
wire n_3117;
wire n_19804;
wire n_13376;
wire n_14377;
wire n_7159;
wire n_3490;
wire n_1622;
wire n_2751;
wire n_1968;
wire n_11282;
wire n_673;
wire n_2842;
wire n_7615;
wire n_3603;
wire n_1978;
wire n_10182;
wire n_14795;
wire n_20773;
wire n_17830;
wire n_8309;
wire n_15685;
wire n_17632;
wire n_19169;
wire n_1164;
wire n_8874;
wire n_12174;
wire n_17288;
wire n_5035;
wire n_1336;
wire n_5453;
wire n_5339;
wire n_17003;
wire n_12289;
wire n_12041;
wire n_13736;
wire n_13254;
wire n_12819;
wire n_17098;
wire n_14810;
wire n_3241;
wire n_16322;
wire n_280;
wire n_12433;
wire n_10413;
wire n_20411;
wire n_17889;
wire n_19466;
wire n_13328;
wire n_16259;
wire n_12550;
wire n_6185;
wire n_15452;
wire n_8344;
wire n_692;
wire n_18674;
wire n_7711;
wire n_4457;
wire n_17173;
wire n_2150;
wire n_17051;
wire n_6643;
wire n_4062;
wire n_6695;
wire n_11593;
wire n_1481;
wire n_4584;
wire n_15074;
wire n_12563;
wire n_2530;
wire n_2299;
wire n_17350;
wire n_16639;
wire n_13624;
wire n_5277;
wire n_792;
wire n_1262;
wire n_13407;
wire n_9447;
wire n_13404;
wire n_18425;
wire n_6213;
wire n_15857;
wire n_14818;
wire n_229;
wire n_18427;
wire n_7958;
wire n_4605;
wire n_5747;
wire n_15714;
wire n_13994;
wire n_11470;
wire n_11294;
wire n_994;
wire n_2428;
wire n_13219;
wire n_17620;
wire n_13737;
wire n_12630;
wire n_20314;
wire n_19683;
wire n_12789;
wire n_12679;
wire n_14084;
wire n_4999;
wire n_13932;
wire n_2872;
wire n_353;
wire n_1678;
wire n_2589;
wire n_15600;
wire n_4086;
wire n_10988;
wire n_13249;
wire n_12338;
wire n_11014;
wire n_5687;
wire n_17169;
wire n_6153;
wire n_15545;
wire n_11310;
wire n_16670;
wire n_3782;
wire n_12675;
wire n_15797;
wire n_6202;
wire n_15353;
wire n_13968;
wire n_7688;
wire n_20389;
wire n_17719;
wire n_9567;
wire n_11773;
wire n_19334;
wire n_5740;
wire n_2501;
wire n_13731;
wire n_12013;
wire n_18349;
wire n_15818;
wire n_16192;
wire n_18667;
wire n_13160;
wire n_7772;
wire n_2028;
wire n_3114;
wire n_11144;
wire n_13385;
wire n_10926;
wire n_20597;
wire n_2773;
wire n_11841;
wire n_2402;
wire n_16342;
wire n_9022;
wire n_387;
wire n_10400;
wire n_13567;
wire n_2808;
wire n_13687;
wire n_8908;
wire n_18068;
wire n_2392;
wire n_9161;
wire n_3272;
wire n_12241;
wire n_10792;
wire n_5898;
wire n_7113;
wire n_13779;
wire n_16124;
wire n_607;
wire n_13722;
wire n_13225;
wire n_18756;
wire n_19022;
wire n_6657;
wire n_10994;
wire n_5617;
wire n_5946;
wire n_1268;
wire n_20392;
wire n_14595;
wire n_14638;
wire n_13039;
wire n_20403;
wire n_702;
wire n_4933;
wire n_4144;
wire n_18564;
wire n_2375;
wire n_6380;
wire n_4895;
wire n_15288;
wire n_9867;
wire n_6163;
wire n_4726;
wire n_10005;
wire n_5573;
wire n_6331;
wire n_311;
wire n_5068;
wire n_15906;
wire n_7363;
wire n_17411;
wire n_2569;
wire n_19218;
wire n_14260;
wire n_10061;
wire n_16790;
wire n_12086;
wire n_269;
wire n_11887;
wire n_14189;
wire n_12281;
wire n_20086;
wire n_4510;
wire n_14552;
wire n_18121;
wire n_446;
wire n_5273;
wire n_10136;
wire n_7588;
wire n_1710;
wire n_18542;
wire n_10369;
wire n_2355;
wire n_18805;
wire n_11703;
wire n_7697;
wire n_17710;
wire n_9027;
wire n_3002;
wire n_18486;
wire n_10194;
wire n_7192;
wire n_1099;
wire n_12807;
wire n_4899;
wire n_3146;
wire n_759;
wire n_4156;
wire n_1727;
wire n_14704;
wire n_14293;
wire n_10223;
wire n_15417;
wire n_3132;
wire n_8881;
wire n_16459;
wire n_9404;
wire n_19629;
wire n_3681;
wire n_13301;
wire n_778;
wire n_2351;
wire n_550;
wire n_17416;
wire n_19165;
wire n_13049;
wire n_1152;
wire n_4579;
wire n_13338;
wire n_6496;
wire n_9352;
wire n_14083;
wire n_17365;
wire n_16167;
wire n_12019;
wire n_2704;
wire n_3729;
wire n_6968;
wire n_13416;
wire n_12255;
wire n_7377;
wire n_9681;
wire n_8353;
wire n_12503;
wire n_2048;
wire n_7723;
wire n_3775;
wire n_9098;
wire n_13053;
wire n_13752;
wire n_14125;
wire n_4753;
wire n_1289;
wire n_1831;
wire n_6292;
wire n_7759;
wire n_16020;
wire n_5754;
wire n_2515;
wire n_1600;
wire n_838;
wire n_1941;
wire n_3637;
wire n_9853;
wire n_16165;
wire n_17403;
wire n_13324;
wire n_16967;
wire n_17961;
wire n_7777;
wire n_12339;
wire n_16482;
wire n_8302;
wire n_14616;
wire n_5756;
wire n_14784;
wire n_20904;
wire n_15301;
wire n_7693;
wire n_11150;
wire n_19082;
wire n_3194;
wire n_2085;
wire n_6408;
wire n_6015;
wire n_18346;
wire n_2097;
wire n_10215;
wire n_19205;
wire n_16844;
wire n_15811;
wire n_20063;
wire n_4203;
wire n_12105;
wire n_16132;
wire n_5789;
wire n_21063;
wire n_5400;
wire n_7558;
wire n_5347;
wire n_14744;
wire n_2957;
wire n_8103;
wire n_8719;
wire n_9778;
wire n_15218;
wire n_14441;
wire n_13159;
wire n_3820;
wire n_14769;
wire n_14732;
wire n_13337;
wire n_5509;
wire n_15433;
wire n_14230;
wire n_11699;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_11817;
wire n_1479;
wire n_14199;
wire n_20754;
wire n_16842;
wire n_1638;
wire n_14722;
wire n_5349;
wire n_14101;
wire n_6472;
wire n_9532;
wire n_3499;
wire n_15586;
wire n_10680;
wire n_16711;
wire n_12564;
wire n_17713;
wire n_18558;
wire n_17306;
wire n_2585;
wire n_16892;
wire n_3361;
wire n_6073;
wire n_20119;
wire n_8834;
wire n_9989;
wire n_8417;
wire n_1732;
wire n_2678;
wire n_17628;
wire n_11621;
wire n_16590;
wire n_18258;
wire n_4556;
wire n_2183;
wire n_11558;
wire n_389;
wire n_18457;
wire n_1707;
wire n_5079;
wire n_20122;
wire n_9406;
wire n_10089;
wire n_19577;
wire n_11113;
wire n_17389;
wire n_2421;
wire n_9160;
wire n_11051;
wire n_13308;
wire n_7712;
wire n_1818;
wire n_6580;
wire n_14791;
wire n_13923;
wire n_14927;
wire n_265;
wire n_20950;
wire n_8599;
wire n_8781;
wire n_5375;
wire n_18145;
wire n_1264;
wire n_7915;
wire n_12655;
wire n_13882;
wire n_3075;
wire n_17650;
wire n_12779;
wire n_1102;
wire n_14085;
wire n_19646;
wire n_15427;
wire n_8244;
wire n_17963;
wire n_12688;
wire n_17368;
wire n_11334;
wire n_20084;
wire n_6795;
wire n_6121;
wire n_457;
wire n_3430;
wire n_2063;
wire n_18825;
wire n_20400;
wire n_11080;
wire n_8367;
wire n_10761;
wire n_14074;
wire n_3484;
wire n_14043;
wire n_13445;
wire n_411;
wire n_4971;
wire n_9521;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_4661;
wire n_3041;
wire n_357;
wire n_412;
wire n_8898;
wire n_1421;
wire n_2423;
wire n_5422;
wire n_8905;
wire n_8145;
wire n_21036;
wire n_7424;
wire n_10216;
wire n_17896;
wire n_9863;
wire n_3832;
wire n_15348;
wire n_10616;
wire n_3525;
wire n_11182;
wire n_20859;
wire n_15754;
wire n_3684;
wire n_10175;
wire n_1681;
wire n_13576;
wire n_5332;
wire n_7149;
wire n_589;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_8211;
wire n_16515;
wire n_1383;
wire n_603;
wire n_19210;
wire n_12788;
wire n_10450;
wire n_15254;
wire n_245;
wire n_13238;
wire n_319;
wire n_690;
wire n_5367;
wire n_20253;
wire n_12866;
wire n_6629;
wire n_16122;
wire n_11158;
wire n_20163;
wire n_19436;
wire n_1837;
wire n_13970;
wire n_10536;
wire n_189;
wire n_9284;
wire n_4953;
wire n_18898;
wire n_7596;
wire n_18572;
wire n_17220;
wire n_11578;
wire n_1246;
wire n_11015;
wire n_5265;
wire n_7549;
wire n_4802;
wire n_17231;
wire n_5733;
wire n_1187;
wire n_14046;
wire n_6918;
wire n_1298;
wire n_9773;
wire n_17971;
wire n_13170;
wire n_8682;
wire n_19887;
wire n_8290;
wire n_13664;
wire n_20130;
wire n_19807;
wire n_17554;
wire n_8890;
wire n_12962;
wire n_12094;
wire n_279;
wire n_9784;
wire n_12964;
wire n_3063;
wire n_14120;
wire n_2288;
wire n_14412;
wire n_14499;
wire n_8275;
wire n_7474;
wire n_7124;
wire n_16911;
wire n_14609;
wire n_9192;
wire n_4581;
wire n_6008;
wire n_665;
wire n_11607;
wire n_2107;
wire n_12838;
wire n_16785;
wire n_18019;
wire n_3679;
wire n_738;
wire n_672;
wire n_11896;
wire n_20692;
wire n_2735;
wire n_14332;
wire n_4214;
wire n_5290;
wire n_15067;
wire n_15223;
wire n_13861;
wire n_19649;
wire n_989;
wire n_2233;
wire n_19872;
wire n_14583;
wire n_11401;
wire n_20933;
wire n_18850;
wire n_4892;
wire n_12514;
wire n_18095;
wire n_16034;
wire n_16389;
wire n_9564;
wire n_11199;
wire n_9127;
wire n_19931;
wire n_8048;
wire n_21116;
wire n_14840;
wire n_4950;
wire n_19900;
wire n_14970;
wire n_7755;
wire n_13135;
wire n_20310;
wire n_15005;
wire n_17156;
wire n_1404;
wire n_16326;
wire n_18698;
wire n_15123;
wire n_3627;
wire n_5214;
wire n_18092;
wire n_5845;
wire n_8868;
wire n_9889;
wire n_293;
wire n_20254;
wire n_13464;
wire n_4454;
wire n_11669;
wire n_2332;
wire n_6005;
wire n_1295;
wire n_2571;
wire n_3049;
wire n_5436;
wire n_12271;
wire n_19839;
wire n_3066;
wire n_12803;
wire n_2045;
wire n_6085;
wire n_11849;
wire n_16874;
wire n_5140;
wire n_19575;
wire n_1597;
wire n_8656;
wire n_9183;
wire n_5847;
wire n_9461;
wire n_6383;
wire n_12773;
wire n_7308;
wire n_12736;
wire n_18814;
wire n_17702;
wire n_5050;
wire n_9062;
wire n_1461;
wire n_10265;
wire n_1830;
wire n_6567;
wire n_16063;
wire n_5658;
wire n_13599;
wire n_15211;
wire n_7290;
wire n_13077;
wire n_19982;
wire n_5546;
wire n_19762;
wire n_7822;
wire n_15643;
wire n_680;
wire n_5289;
wire n_14251;
wire n_15911;
wire n_18236;
wire n_12239;
wire n_16628;
wire n_11085;
wire n_16047;
wire n_19760;
wire n_1274;
wire n_7632;
wire n_17075;
wire n_475;
wire n_17387;
wire n_2703;
wire n_6314;
wire n_13162;
wire n_19442;
wire n_5610;
wire n_8576;
wire n_916;
wire n_1884;
wire n_20665;
wire n_18943;
wire n_2683;
wire n_18361;
wire n_4180;
wire n_15309;
wire n_18932;
wire n_17299;
wire n_7289;
wire n_15790;
wire n_16521;
wire n_14488;
wire n_4642;
wire n_13952;
wire n_7473;
wire n_15890;
wire n_1750;
wire n_16468;
wire n_3544;
wire n_6845;
wire n_10451;
wire n_10768;
wire n_3852;
wire n_16429;
wire n_19213;
wire n_5233;
wire n_16611;
wire n_19311;
wire n_20934;
wire n_7483;
wire n_13868;
wire n_5710;
wire n_1491;
wire n_3219;
wire n_274;
wire n_5333;
wire n_5799;
wire n_8976;
wire n_13694;
wire n_10312;
wire n_4587;
wire n_16682;
wire n_14325;
wire n_19130;
wire n_16453;
wire n_14998;
wire n_8844;
wire n_19576;
wire n_6357;
wire n_3479;
wire n_5499;
wire n_9123;
wire n_19454;
wire n_4150;
wire n_20295;
wire n_12545;
wire n_8669;
wire n_4285;
wire n_12531;
wire n_11290;
wire n_19978;
wire n_9922;
wire n_20543;
wire n_1908;
wire n_712;
wire n_8769;
wire n_9463;
wire n_18607;
wire n_18165;
wire n_12916;
wire n_1392;
wire n_15198;
wire n_16860;
wire n_6087;
wire n_17852;
wire n_13246;
wire n_19143;
wire n_19647;
wire n_20755;
wire n_10135;
wire n_20533;
wire n_7664;
wire n_14329;
wire n_16782;
wire n_16432;
wire n_14428;
wire n_18272;
wire n_8990;
wire n_1914;
wire n_8208;
wire n_12692;
wire n_7714;
wire n_12976;
wire n_14660;
wire n_20221;
wire n_2130;
wire n_13984;
wire n_19899;
wire n_18359;
wire n_9843;
wire n_20100;
wire n_3187;
wire n_19391;
wire n_11619;
wire n_479;
wire n_5564;
wire n_16779;
wire n_18807;
wire n_3082;
wire n_15641;
wire n_2473;
wire n_12946;
wire n_16298;
wire n_19293;
wire n_16830;
wire n_13449;
wire n_14620;
wire n_18342;
wire n_6103;
wire n_18362;
wire n_2565;
wire n_1237;
wire n_12286;
wire n_5883;
wire n_14134;
wire n_13995;
wire n_3078;
wire n_12146;
wire n_7680;
wire n_6666;
wire n_5117;
wire n_9362;
wire n_13483;
wire n_1531;
wire n_17822;
wire n_6207;
wire n_9712;
wire n_18649;
wire n_13614;
wire n_11202;
wire n_9460;
wire n_18246;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_17444;
wire n_11227;
wire n_5975;
wire n_18837;
wire n_14502;
wire n_15367;
wire n_1951;
wire n_12557;
wire n_2558;
wire n_7061;
wire n_9068;
wire n_3104;
wire n_6661;
wire n_17857;
wire n_19848;
wire n_14750;
wire n_10228;
wire n_14518;
wire n_15704;
wire n_20406;
wire n_4952;
wire n_5699;
wire n_9348;
wire n_11125;
wire n_15209;
wire n_5920;
wire n_20197;
wire n_2112;
wire n_9632;
wire n_21126;
wire n_19214;
wire n_2237;
wire n_11951;
wire n_5211;
wire n_9257;
wire n_19164;
wire n_5535;
wire n_14467;
wire n_7783;
wire n_6057;
wire n_14898;
wire n_9049;
wire n_18615;
wire n_17980;
wire n_7990;
wire n_10433;
wire n_18562;
wire n_10231;
wire n_10929;
wire n_15300;
wire n_18830;
wire n_14656;
wire n_3968;
wire n_17262;
wire n_2841;
wire n_3332;
wire n_8300;
wire n_7501;
wire n_11383;
wire n_19736;
wire n_2998;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_13540;
wire n_2822;
wire n_13642;
wire n_14764;
wire n_17329;
wire n_2937;
wire n_4293;
wire n_18497;
wire n_16290;
wire n_4039;
wire n_14632;
wire n_6926;
wire n_17413;
wire n_9067;
wire n_703;
wire n_20529;
wire n_18334;
wire n_3385;
wire n_15372;
wire n_227;
wire n_17358;
wire n_12735;
wire n_14510;
wire n_7917;
wire n_4942;
wire n_15388;
wire n_536;
wire n_10425;
wire n_12254;
wire n_4348;
wire n_1602;
wire n_9299;
wire n_3139;
wire n_11298;
wire n_16232;
wire n_9244;
wire n_14667;
wire n_5261;
wire n_16871;
wire n_17292;
wire n_12124;
wire n_12494;
wire n_3636;
wire n_16529;
wire n_3823;
wire n_3403;
wire n_12051;
wire n_9911;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_14802;
wire n_18031;
wire n_13637;
wire n_7572;
wire n_16603;
wire n_2944;
wire n_2780;
wire n_1202;
wire n_627;
wire n_2033;
wire n_4121;
wire n_16838;
wire n_18593;
wire n_11363;
wire n_3984;
wire n_8728;
wire n_20693;
wire n_19438;
wire n_6200;
wire n_12612;
wire n_8407;
wire n_13423;
wire n_11636;
wire n_14926;
wire n_17048;
wire n_18463;
wire n_6902;
wire n_12798;
wire n_16993;
wire n_7197;
wire n_3737;
wire n_16685;
wire n_11313;
wire n_17602;
wire n_15182;
wire n_9072;
wire n_12635;
wire n_2300;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_551;
wire n_4521;
wire n_13139;
wire n_19133;
wire n_19257;
wire n_12874;
wire n_8511;
wire n_2283;
wire n_5206;
wire n_582;
wire n_13356;
wire n_20309;
wire n_2508;
wire n_10344;
wire n_9459;
wire n_5298;
wire n_17366;
wire n_3417;
wire n_8246;
wire n_9655;
wire n_3626;
wire n_12048;
wire n_17566;
wire n_20354;
wire n_8925;
wire n_7881;
wire n_4789;
wire n_19953;
wire n_12829;
wire n_17854;
wire n_1081;
wire n_9678;
wire n_18833;
wire n_2493;
wire n_9560;
wire n_15036;
wire n_12528;
wire n_4565;
wire n_7032;
wire n_16061;
wire n_9303;
wire n_19226;
wire n_12371;
wire n_20852;
wire n_18257;
wire n_14866;
wire n_6884;
wire n_7752;
wire n_8201;
wire n_3512;
wire n_1860;
wire n_8046;
wire n_6287;
wire n_14575;
wire n_14005;
wire n_4172;
wire n_8414;
wire n_5567;
wire n_8292;
wire n_9138;
wire n_11936;
wire n_12071;
wire n_11543;
wire n_6067;
wire n_2280;
wire n_12578;
wire n_18339;
wire n_12311;
wire n_13253;
wire n_456;
wire n_13647;
wire n_9179;
wire n_2468;
wire n_2171;
wire n_11056;
wire n_14241;
wire n_16275;
wire n_2035;
wire n_7196;
wire n_10916;
wire n_14693;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_8187;
wire n_10108;
wire n_10661;
wire n_19245;
wire n_5817;
wire n_16587;
wire n_18731;
wire n_16400;
wire n_9504;
wire n_5417;
wire n_18876;
wire n_14118;
wire n_19235;
wire n_9285;
wire n_15068;
wire n_13088;
wire n_10963;
wire n_11146;
wire n_3097;
wire n_4395;
wire n_10788;
wire n_16161;
wire n_1215;
wire n_11830;
wire n_14577;
wire n_3748;
wire n_13026;
wire n_10471;
wire n_20916;
wire n_211;
wire n_1804;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5989;
wire n_13116;
wire n_1769;
wire n_4319;
wire n_9360;
wire n_14323;
wire n_10099;
wire n_20041;
wire n_10193;
wire n_14096;
wire n_4874;
wire n_516;
wire n_1997;
wire n_10140;
wire n_7867;
wire n_19930;
wire n_10149;
wire n_3167;
wire n_4748;
wire n_13828;
wire n_16441;
wire n_19434;
wire n_10576;
wire n_4025;
wire n_1321;
wire n_16984;
wire n_14301;
wire n_19342;
wire n_10682;
wire n_752;
wire n_7543;
wire n_9659;
wire n_17491;
wire n_12204;
wire n_13643;
wire n_20369;
wire n_17302;
wire n_2412;
wire n_14774;
wire n_19476;
wire n_3107;
wire n_9013;
wire n_9427;
wire n_226;
wire n_20381;
wire n_7019;
wire n_5315;
wire n_3708;
wire n_15540;
wire n_1778;
wire n_584;
wire n_10237;
wire n_9538;
wire n_19294;
wire n_19668;
wire n_16491;
wire n_19398;
wire n_4082;
wire n_979;
wire n_14471;
wire n_3381;
wire n_11170;
wire n_20935;
wire n_19733;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_4466;
wire n_3955;
wire n_1887;
wire n_19277;
wire n_15040;
wire n_18307;
wire n_11457;
wire n_7199;
wire n_15731;
wire n_2170;
wire n_4721;
wire n_19798;
wire n_9924;
wire n_9159;
wire n_16662;
wire n_16225;
wire n_3840;
wire n_7166;
wire n_5369;
wire n_9476;
wire n_16496;
wire n_3809;
wire n_801;
wire n_19080;
wire n_14800;
wire n_7923;
wire n_11058;
wire n_6327;
wire n_5853;
wire n_3468;
wire n_12203;
wire n_15606;
wire n_20456;
wire n_11403;
wire n_19280;
wire n_272;
wire n_14099;
wire n_20465;
wire n_18685;
wire n_11741;
wire n_4561;
wire n_3291;
wire n_8095;
wire n_18860;
wire n_11365;
wire n_13291;
wire n_14756;
wire n_1472;
wire n_17237;
wire n_8735;
wire n_15073;
wire n_2475;
wire n_8902;
wire n_12869;
wire n_8796;
wire n_2715;
wire n_14413;
wire n_18204;
wire n_5044;
wire n_210;
wire n_3755;
wire n_4536;
wire n_11141;
wire n_14753;
wire n_8549;
wire n_14161;
wire n_5459;
wire n_19072;
wire n_10716;
wire n_224;
wire n_11238;
wire n_11406;
wire n_2854;
wire n_16000;
wire n_10443;
wire n_19485;
wire n_3341;
wire n_19686;
wire n_16557;
wire n_19232;
wire n_12954;
wire n_1116;
wire n_5024;
wire n_2747;
wire n_19452;
wire n_1511;
wire n_15393;
wire n_8593;
wire n_10912;
wire n_20699;
wire n_19752;
wire n_10469;
wire n_17626;
wire n_9649;
wire n_19095;
wire n_15864;
wire n_3731;
wire n_4412;
wire n_7649;
wire n_18645;
wire n_15628;
wire n_16788;
wire n_12004;
wire n_6704;
wire n_9090;
wire n_2003;
wire n_2533;
wire n_9696;
wire n_14181;
wire n_9996;
wire n_4810;
wire n_21102;
wire n_10405;
wire n_9498;
wire n_10390;
wire n_1370;
wire n_9836;
wire n_5005;
wire n_14570;
wire n_20196;
wire n_16191;
wire n_12912;
wire n_8596;
wire n_9938;
wire n_16467;
wire n_20503;
wire n_10867;
wire n_11847;
wire n_16697;
wire n_20846;
wire n_10092;
wire n_3620;
wire n_18067;
wire n_2767;
wire n_5474;
wire n_16371;
wire n_181;
wire n_9743;
wire n_9121;
wire n_16661;
wire n_11237;
wire n_12005;
wire n_16493;
wire n_1300;
wire n_1960;
wire n_10738;
wire n_5700;
wire n_16961;
wire n_2862;
wire n_4325;
wire n_14501;
wire n_4711;
wire n_16780;
wire n_12302;
wire n_11432;
wire n_20080;
wire n_3307;
wire n_3288;
wire n_9216;
wire n_9563;
wire n_17493;
wire n_15229;
wire n_7941;
wire n_13010;
wire n_5662;
wire n_14738;
wire n_8858;
wire n_3880;
wire n_3904;
wire n_15504;
wire n_13703;
wire n_3008;
wire n_4821;
wire n_10813;
wire n_19705;
wire n_15403;
wire n_14291;
wire n_14761;
wire n_7074;
wire n_11707;
wire n_10899;
wire n_11728;
wire n_16137;
wire n_171;
wire n_14388;
wire n_19831;
wire n_14932;
wire n_6184;
wire n_1040;
wire n_4138;
wire n_1444;
wire n_12723;
wire n_10334;
wire n_2882;
wire n_14674;
wire n_11688;
wire n_9794;
wire n_16062;
wire n_10726;
wire n_16210;
wire n_13486;
wire n_20798;
wire n_9550;
wire n_20688;
wire n_6711;
wire n_11696;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_10635;
wire n_11681;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_6007;
wire n_10852;
wire n_14893;
wire n_13789;
wire n_1772;
wire n_14354;
wire n_19652;
wire n_6879;
wire n_15442;
wire n_9896;
wire n_9612;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_6303;
wire n_19985;
wire n_3092;
wire n_7692;
wire n_5397;
wire n_9272;
wire n_13055;
wire n_9645;
wire n_14283;
wire n_880;
wire n_5566;
wire n_16392;
wire n_9697;
wire n_15307;
wire n_20459;
wire n_4388;
wire n_10901;
wire n_15855;
wire n_19224;
wire n_7131;
wire n_17943;
wire n_13839;
wire n_9929;
wire n_13898;
wire n_7042;
wire n_9859;
wire n_2809;
wire n_19504;
wire n_16375;
wire n_932;
wire n_2276;
wire n_5492;
wire n_8077;
wire n_11242;
wire n_2465;
wire n_15445;
wire n_12917;
wire n_14711;
wire n_16586;
wire n_17158;
wire n_2972;
wire n_7391;
wire n_13819;
wire n_13990;
wire n_15745;
wire n_3721;
wire n_11253;
wire n_13193;
wire n_2425;
wire n_15648;
wire n_5692;
wire n_15887;
wire n_7981;
wire n_13037;
wire n_1601;
wire n_12188;
wire n_17603;
wire n_5473;
wire n_12575;
wire n_14698;
wire n_10372;
wire n_1011;
wire n_4286;
wire n_18754;
wire n_3638;
wire n_18537;
wire n_13127;
wire n_12598;
wire n_4858;
wire n_5370;
wire n_13561;
wire n_7378;
wire n_15922;
wire n_16938;
wire n_15987;
wire n_7836;
wire n_12626;
wire n_10960;
wire n_10712;
wire n_2387;
wire n_4318;
wire n_16849;
wire n_8910;
wire n_20337;
wire n_16412;
wire n_16070;
wire n_5227;
wire n_14091;
wire n_14842;
wire n_15981;
wire n_20162;
wire n_10100;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_5359;
wire n_19407;
wire n_5282;
wire n_13539;
wire n_499;
wire n_10162;
wire n_9840;
wire n_15471;
wire n_4738;
wire n_19534;
wire n_11399;
wire n_20599;
wire n_6215;
wire n_12676;
wire n_8252;
wire n_20300;
wire n_3663;
wire n_9491;
wire n_10337;
wire n_12999;
wire n_10264;
wire n_6569;
wire n_16710;
wire n_15355;
wire n_9992;
wire n_14089;
wire n_8278;
wire n_18090;
wire n_443;
wire n_12362;
wire n_5716;
wire n_12360;
wire n_139;
wire n_13570;
wire n_6605;
wire n_16356;
wire n_16182;
wire n_16103;
wire n_8683;
wire n_956;
wire n_6544;
wire n_21014;
wire n_15241;
wire n_6332;
wire n_399;
wire n_7130;
wire n_15729;
wire n_6680;
wire n_3575;
wire n_6310;
wire n_9695;
wire n_13411;
wire n_19947;
wire n_16240;
wire n_11526;
wire n_20422;
wire n_1937;
wire n_6259;
wire n_3004;
wire n_15371;
wire n_9800;
wire n_1285;
wire n_10745;
wire n_193;
wire n_12733;
wire n_18634;
wire n_5445;
wire n_7227;
wire n_16650;
wire n_14299;
wire n_18247;
wire n_7813;
wire n_13332;
wire n_16280;
wire n_9085;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_11302;
wire n_9899;
wire n_18678;
wire n_16898;
wire n_12261;
wire n_11561;
wire n_19264;
wire n_14198;
wire n_5628;
wire n_5245;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_9042;
wire n_1754;
wire n_9570;
wire n_11054;
wire n_9644;
wire n_1172;
wire n_2775;
wire n_18423;
wire n_6769;
wire n_16301;
wire n_20405;
wire n_6844;
wire n_18366;
wire n_13582;
wire n_8700;
wire n_19810;
wire n_13255;
wire n_18691;
wire n_2657;
wire n_18961;
wire n_7802;
wire n_16869;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_15851;
wire n_5860;
wire n_6416;
wire n_7515;
wire n_3387;
wire n_10408;
wire n_17718;
wire n_13424;
wire n_4349;
wire n_20751;
wire n_6945;
wire n_8378;
wire n_18176;
wire n_6491;
wire n_10562;
wire n_10893;
wire n_449;
wire n_7914;
wire n_17017;
wire n_6447;
wire n_4390;
wire n_459;
wire n_17088;
wire n_1782;
wire n_11517;
wire n_13716;
wire n_9523;
wire n_4380;
wire n_4609;
wire n_7325;
wire n_14561;
wire n_18248;
wire n_723;
wire n_1393;
wire n_7674;
wire n_20769;
wire n_9829;
wire n_20906;
wire n_13914;
wire n_11579;
wire n_19347;
wire n_17803;
wire n_14119;
wire n_18689;
wire n_7983;
wire n_641;
wire n_18110;
wire n_16397;
wire n_19856;
wire n_11640;
wire n_9153;
wire n_4700;
wire n_4002;
wire n_14825;
wire n_21092;
wire n_11656;
wire n_3815;
wire n_14007;
wire n_2982;
wire n_8653;
wire n_19031;
wire n_17837;
wire n_18164;
wire n_17407;
wire n_8601;
wire n_1043;
wire n_2869;
wire n_12835;
wire n_7079;
wire n_11572;
wire n_9789;
wire n_16694;
wire n_16893;
wire n_5820;
wire n_20266;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_14426;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_16653;
wire n_10012;
wire n_196;
wire n_14957;
wire n_17706;
wire n_12348;
wire n_10939;
wire n_17506;
wire n_3112;
wire n_954;
wire n_10008;
wire n_2051;
wire n_9795;
wire n_16538;
wire n_3196;
wire n_16834;
wire n_19955;
wire n_664;
wire n_13203;
wire n_5126;
wire n_8659;
wire n_6732;
wire n_2381;
wire n_1967;
wire n_1280;
wire n_15408;
wire n_544;
wire n_15184;
wire n_13052;
wire n_7668;
wire n_7435;
wire n_20215;
wire n_17265;
wire n_18507;
wire n_3923;
wire n_5603;
wire n_6560;
wire n_17614;
wire n_9847;
wire n_13846;
wire n_15961;
wire n_20832;
wire n_7848;
wire n_13312;
wire n_2596;
wire n_8337;
wire n_3986;
wire n_18779;
wire n_5909;
wire n_11289;
wire n_147;
wire n_18471;
wire n_1211;
wire n_11157;
wire n_16178;
wire n_14718;
wire n_11013;
wire n_7653;
wire n_12885;
wire n_1644;
wire n_8347;
wire n_1252;
wire n_18963;
wire n_773;
wire n_17955;
wire n_16845;
wire n_15605;
wire n_17612;
wire n_6655;
wire n_718;
wire n_12073;
wire n_20148;
wire n_8899;
wire n_2573;
wire n_6480;
wire n_5837;
wire n_11836;
wire n_2336;
wire n_5412;
wire n_20804;
wire n_8481;
wire n_3483;
wire n_11747;
wire n_1925;
wire n_20662;
wire n_7420;
wire n_15914;
wire n_20451;
wire n_16954;
wire n_19908;
wire n_10115;
wire n_16749;
wire n_19505;
wire n_17102;
wire n_12585;
wire n_12963;
wire n_12029;
wire n_16769;
wire n_9827;
wire n_1574;
wire n_18057;
wire n_14748;
wire n_20391;
wire n_1981;
wire n_17683;
wire n_15318;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_531;
wire n_20081;
wire n_16636;
wire n_6283;
wire n_4939;
wire n_11758;
wire n_17864;
wire n_9400;
wire n_18863;
wire n_10744;
wire n_691;
wire n_6819;
wire n_4903;
wire n_17004;
wire n_20209;
wire n_4382;
wire n_423;
wire n_6898;
wire n_14838;
wire n_17691;
wire n_15620;
wire n_20142;
wire n_16905;
wire n_11958;
wire n_16717;
wire n_10009;
wire n_7244;
wire n_16293;
wire n_4626;
wire n_10072;
wire n_12699;
wire n_20629;
wire n_8750;
wire n_13657;
wire n_20501;
wire n_9104;
wire n_8637;
wire n_4638;
wire n_8792;
wire n_7286;
wire n_7857;
wire n_13871;
wire n_18149;
wire n_3719;
wire n_16840;
wire n_17534;
wire n_3888;
wire n_9960;
wire n_14843;
wire n_5295;
wire n_13881;
wire n_8390;
wire n_1181;
wire n_16072;
wire n_17994;
wire n_10002;
wire n_9601;
wire n_20794;
wire n_13137;
wire n_13226;
wire n_18652;
wire n_15951;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_20833;
wire n_17465;
wire n_18735;
wire n_12006;
wire n_3943;
wire n_7964;
wire n_11322;
wire n_11484;
wire n_9972;
wire n_2908;
wire n_8594;
wire n_14183;
wire n_9541;
wire n_18653;
wire n_1184;
wire n_17084;
wire n_14528;
wire n_1073;
wire n_4549;
wire n_19570;
wire n_1062;
wire n_5102;
wire n_9974;
wire n_18597;
wire n_16889;
wire n_1974;
wire n_8425;
wire n_13001;
wire n_6959;
wire n_11803;
wire n_4331;
wire n_4159;
wire n_16458;
wire n_13784;
wire n_21115;
wire n_11139;
wire n_3451;
wire n_8051;
wire n_11021;
wire n_17613;
wire n_2832;
wire n_1944;
wire n_267;
wire n_5656;
wire n_1988;
wire n_15996;
wire n_6561;
wire n_5865;
wire n_13271;
wire n_12096;
wire n_2277;
wire n_16507;
wire n_10125;
wire n_14770;
wire n_787;
wire n_16829;
wire n_13761;
wire n_1522;
wire n_4760;
wire n_13190;
wire n_10693;
wire n_14461;
wire n_1314;
wire n_8755;
wire n_13174;
wire n_16028;
wire n_20039;
wire n_18061;
wire n_5407;
wire n_2988;
wire n_12814;
wire n_11553;
wire n_4560;
wire n_14322;
wire n_17561;
wire n_12009;
wire n_13916;
wire n_7761;
wire n_5042;
wire n_859;
wire n_1889;
wire n_6090;
wire n_18829;
wire n_3641;
wire n_16707;
wire n_16674;
wire n_19399;
wire n_15171;
wire n_3183;
wire n_11926;
wire n_8383;
wire n_2885;
wire n_14585;
wire n_7437;
wire n_11460;
wire n_8895;
wire n_20500;
wire n_4987;
wire n_1396;
wire n_4988;
wire n_10728;
wire n_15109;
wire n_6620;
wire n_9220;
wire n_16676;
wire n_20645;
wire n_4540;
wire n_19315;
wire n_13965;
wire n_17130;
wire n_8665;
wire n_21053;
wire n_3652;
wire n_14640;
wire n_9444;
wire n_17809;
wire n_10497;
wire n_12082;
wire n_13966;
wire n_14936;
wire n_12322;
wire n_1416;
wire n_19812;
wire n_21062;
wire n_18063;
wire n_8303;
wire n_13981;
wire n_5871;
wire n_17221;
wire n_6052;
wire n_7769;
wire n_11416;
wire n_14360;
wire n_9193;
wire n_19326;
wire n_20183;
wire n_8852;
wire n_20366;
wire n_20578;
wire n_20277;
wire n_6488;
wire n_9755;
wire n_19243;
wire n_4502;
wire n_7005;
wire n_5334;
wire n_1590;
wire n_4115;
wire n_16942;
wire n_5019;
wire n_17907;
wire n_14828;
wire n_1819;
wire n_9162;
wire n_15264;
wire n_947;
wire n_7341;
wire n_5792;
wire n_20890;
wire n_19114;
wire n_468;
wire n_19321;
wire n_182;
wire n_696;
wire n_482;
wire n_1833;
wire n_16142;
wire n_12833;
wire n_2499;
wire n_16091;
wire n_6649;
wire n_15424;
wire n_8357;
wire n_1382;
wire n_2970;
wire n_4264;
wire n_5954;
wire n_10326;
wire n_14827;
wire n_3192;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_20306;
wire n_13363;
wire n_8587;
wire n_7285;
wire n_1972;
wire n_4718;
wire n_10725;
wire n_6324;
wire n_5489;
wire n_15653;
wire n_10274;
wire n_17969;
wire n_4029;
wire n_14780;
wire n_12340;
wire n_10799;
wire n_8922;
wire n_3193;
wire n_18240;
wire n_8498;
wire n_669;
wire n_4170;
wire n_12184;
wire n_19138;
wire n_12472;
wire n_13048;
wire n_20814;
wire n_12266;
wire n_19388;
wire n_12432;
wire n_517;
wire n_6041;
wire n_8526;
wire n_13593;
wire n_8319;
wire n_6859;
wire n_10732;
wire n_20528;
wire n_16851;
wire n_15310;
wire n_144;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_12122;
wire n_18065;
wire n_14889;
wire n_20538;
wire n_17773;
wire n_8214;
wire n_18265;
wire n_8516;
wire n_815;
wire n_12310;
wire n_11343;
wire n_8989;
wire n_7746;
wire n_11362;
wire n_20278;
wire n_1433;
wire n_3912;
wire n_16119;
wire n_10720;
wire n_19221;
wire n_19586;
wire n_20550;
wire n_15050;
wire n_17469;
wire n_12827;
wire n_18422;
wire n_21065;
wire n_9217;
wire n_20060;
wire n_6747;
wire n_2903;
wire n_12804;
wire n_3812;
wire n_11347;
wire n_7957;
wire n_2378;
wire n_5530;
wire n_16440;
wire n_6718;
wire n_965;
wire n_13804;
wire n_17357;
wire n_12418;
wire n_19074;
wire n_8087;
wire n_4056;
wire n_10238;
wire n_17887;
wire n_5993;
wire n_19956;
wire n_9948;
wire n_7687;
wire n_18583;
wire n_2142;
wire n_15396;
wire n_4043;
wire n_15038;
wire n_3170;
wire n_1455;
wire n_836;
wire n_6975;
wire n_3464;
wire n_7703;
wire n_11760;
wire n_15781;
wire n_10395;
wire n_1483;
wire n_8722;
wire n_17376;
wire n_970;
wire n_15306;
wire n_713;
wire n_3179;
wire n_12187;
wire n_7665;
wire n_4836;
wire n_7677;
wire n_15978;
wire n_10366;
wire n_14017;
wire n_6663;
wire n_14145;
wire n_1419;
wire n_13406;
wire n_10431;
wire n_8622;
wire n_11485;
wire n_3528;
wire n_12453;
wire n_15984;
wire n_4207;
wire n_20551;
wire n_2404;
wire n_9597;
wire n_10614;
wire n_10786;
wire n_16067;
wire n_18123;
wire n_8947;
wire n_15079;
wire n_9983;
wire n_5943;
wire n_6556;
wire n_20049;
wire n_4880;
wire n_15784;
wire n_4051;
wire n_13070;
wire n_17799;
wire n_2996;
wire n_15231;
wire n_6365;
wire n_11417;
wire n_7111;
wire n_5284;
wire n_8786;
wire n_9414;
wire n_11677;
wire n_3246;
wire n_980;
wire n_1869;
wire n_3623;
wire n_11898;
wire n_14749;
wire n_7284;
wire n_3615;
wire n_17675;
wire n_20058;
wire n_13457;
wire n_18479;
wire n_2811;
wire n_9152;
wire n_145;
wire n_2146;
wire n_3276;
wire n_7064;
wire n_19658;
wire n_19907;
wire n_9533;
wire n_18588;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_7799;
wire n_5698;
wire n_21110;
wire n_8871;
wire n_1456;
wire n_14627;
wire n_15552;
wire n_14735;
wire n_15808;
wire n_15103;
wire n_20948;
wire n_2129;
wire n_17647;
wire n_18916;
wire n_553;
wire n_13547;
wire n_578;
wire n_18976;
wire n_8371;
wire n_2975;
wire n_8547;
wire n_11538;
wire n_10815;
wire n_11008;
wire n_4075;
wire n_600;
wire n_20412;
wire n_10424;
wire n_15500;
wire n_502;
wire n_19883;
wire n_16522;
wire n_15543;
wire n_14823;
wire n_5209;
wire n_15807;
wire n_10684;
wire n_13154;
wire n_5704;
wire n_16074;
wire n_4889;
wire n_20780;
wire n_17456;
wire n_19923;
wire n_18666;
wire n_18694;
wire n_3618;
wire n_10184;
wire n_3705;
wire n_1709;
wire n_19472;
wire n_18984;
wire n_11885;
wire n_3974;
wire n_16644;
wire n_9208;
wire n_7792;
wire n_11657;
wire n_13124;
wire n_16327;
wire n_10924;
wire n_14991;
wire n_2853;
wire n_3350;
wire n_8633;
wire n_12897;
wire n_9392;
wire n_7390;
wire n_6111;
wire n_5219;
wire n_920;
wire n_15338;
wire n_18302;
wire n_15866;
wire n_14162;
wire n_15880;
wire n_4261;
wire n_15508;
wire n_18993;
wire n_15292;
wire n_1132;
wire n_501;
wire n_18300;
wire n_18621;
wire n_14566;
wire n_15694;
wire n_7530;
wire n_10129;
wire n_16475;
wire n_1402;
wire n_18347;
wire n_3957;
wire n_13844;
wire n_19198;
wire n_7471;
wire n_19881;
wire n_9328;
wire n_18262;
wire n_10192;
wire n_17137;
wire n_19078;
wire n_20771;
wire n_18139;
wire n_16606;
wire n_11846;
wire n_16560;
wire n_14857;
wire n_7058;
wire n_4648;
wire n_8011;
wire n_19714;
wire n_2214;
wire n_6730;
wire n_11530;
wire n_18498;
wire n_6367;
wire n_8222;
wire n_20232;
wire n_12825;
wire n_2732;
wire n_15907;
wire n_8206;
wire n_8065;
wire n_9914;
wire n_19272;
wire n_18897;
wire n_2949;
wire n_16861;
wire n_7008;
wire n_12918;
wire n_1927;
wire n_16533;
wire n_14600;
wire n_12077;
wire n_16313;
wire n_7139;
wire n_10384;
wire n_17317;
wire n_19265;
wire n_16158;
wire n_19012;
wire n_10885;
wire n_11002;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_16620;
wire n_20348;
wire n_20463;
wire n_19719;
wire n_11648;
wire n_14289;
wire n_18197;
wire n_1572;
wire n_8568;
wire n_17118;
wire n_11734;
wire n_12645;
wire n_18293;
wire n_10003;
wire n_11050;
wire n_17689;
wire n_1388;
wire n_18131;
wire n_14485;
wire n_15277;
wire n_12987;
wire n_4396;
wire n_20871;
wire n_1990;
wire n_12251;
wire n_19408;
wire n_17165;
wire n_16379;
wire n_6667;
wire n_17326;
wire n_9838;
wire n_3491;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_20316;
wire n_8836;
wire n_4228;
wire n_12700;
wire n_12602;
wire n_20549;
wire n_19747;
wire n_3065;
wire n_18796;
wire n_16799;
wire n_11318;
wire n_7060;
wire n_12367;
wire n_17282;
wire n_6750;
wire n_4931;
wire n_20941;
wire n_7790;
wire n_20298;
wire n_20803;
wire n_13492;
wire n_10840;
wire n_5181;
wire n_3208;
wire n_20777;
wire n_14589;
wire n_1342;
wire n_8120;
wire n_21124;
wire n_19532;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_5963;
wire n_19538;
wire n_7532;
wire n_14899;
wire n_12703;
wire n_17311;
wire n_9215;
wire n_5972;
wire n_7065;
wire n_6177;
wire n_5937;
wire n_18278;
wire n_14714;
wire n_15897;
wire n_7267;
wire n_15069;
wire n_12445;
wire n_20120;
wire n_6460;
wire n_9595;
wire n_19680;
wire n_11420;
wire n_1605;
wire n_11527;
wire n_15133;
wire n_18113;
wire n_17899;
wire n_13826;
wire n_2984;
wire n_157;
wire n_18858;
wire n_7619;
wire n_18196;
wire n_2489;
wire n_15832;
wire n_17396;
wire n_13078;
wire n_4145;
wire n_6852;
wire n_15709;
wire n_624;
wire n_13516;
wire n_13557;
wire n_7883;
wire n_5872;
wire n_10397;
wire n_6692;
wire n_9707;
wire n_19105;
wire n_8854;
wire n_12834;
wire n_10202;
wire n_19607;
wire n_12821;
wire n_17653;
wire n_7220;
wire n_2106;
wire n_9262;
wire n_11964;
wire n_12247;
wire n_17033;
wire n_854;
wire n_2091;
wire n_393;
wire n_13065;
wire n_7270;
wire n_8621;
wire n_13753;
wire n_2348;
wire n_19677;
wire n_9806;
wire n_9019;
wire n_14796;
wire n_17793;
wire n_13175;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_17087;
wire n_20615;
wire n_5846;
wire n_9814;
wire n_15361;
wire n_5930;
wire n_17815;
wire n_13823;
wire n_20294;
wire n_11985;
wire n_7458;
wire n_1824;
wire n_3543;
wire n_9856;
wire n_8421;
wire n_19969;
wire n_1776;
wire n_7433;
wire n_3609;
wire n_6334;
wire n_8911;
wire n_9518;
wire n_18509;
wire n_5572;
wire n_10335;
wire n_2570;
wire n_2789;
wire n_17589;
wire n_13658;
wire n_18883;
wire n_807;
wire n_6355;
wire n_7015;
wire n_10567;
wire n_18699;
wire n_7987;
wire n_9009;
wire n_14137;
wire n_802;
wire n_17345;
wire n_20127;
wire n_960;
wire n_7272;
wire n_15505;
wire n_2352;
wire n_12628;
wire n_9722;
wire n_20225;
wire n_5416;
wire n_20892;
wire n_16302;
wire n_11260;
wire n_16305;
wire n_9760;
wire n_6018;
wire n_14320;
wire n_11605;
wire n_13156;
wire n_4611;
wire n_5797;
wire n_7815;
wire n_1052;
wire n_19593;
wire n_11629;
wire n_13119;
wire n_16883;
wire n_20582;
wire n_4399;
wire n_20598;
wire n_8280;
wire n_16094;
wire n_169;
wire n_12156;
wire n_13409;
wire n_2796;
wire n_13832;
wire n_17577;
wire n_5393;
wire n_7352;
wire n_8427;
wire n_4755;
wire n_2771;
wire n_6322;
wire n_2947;
wire n_11466;
wire n_15270;
wire n_928;
wire n_12632;
wire n_6419;
wire n_18715;
wire n_13581;
wire n_748;
wire n_7903;
wire n_16282;
wire n_7089;
wire n_8217;
wire n_20626;
wire n_9331;
wire n_7604;
wire n_2999;
wire n_988;
wire n_15649;
wire n_330;
wire n_328;
wire n_8285;
wire n_8521;
wire n_12446;
wire n_7803;
wire n_20575;
wire n_14526;
wire n_16497;
wire n_11690;
wire n_5986;
wire n_9355;
wire n_16206;
wire n_18642;
wire n_16730;
wire n_7622;
wire n_11968;
wire n_429;
wire n_7839;
wire n_6792;
wire n_19312;
wire n_5794;
wire n_8136;
wire n_20858;
wire n_3476;
wire n_16455;
wire n_11797;
wire n_13672;
wire n_8386;
wire n_6123;
wire n_10802;
wire n_15317;
wire n_1356;
wire n_21100;
wire n_2666;
wire n_20365;
wire n_4409;
wire n_4191;
wire n_11991;
wire n_7072;
wire n_3827;
wire n_11618;
wire n_911;
wire n_19212;
wire n_623;
wire n_11502;
wire n_1403;
wire n_5395;
wire n_18590;
wire n_8857;
wire n_9495;
wire n_10987;
wire n_236;
wire n_12063;
wire n_10551;
wire n_10646;
wire n_13471;
wire n_13021;
wire n_15589;
wire n_15322;
wire n_3790;
wire n_7960;
wire n_14967;
wire n_6152;
wire n_18465;
wire n_17635;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_10538;
wire n_15557;
wire n_10199;
wire n_1694;
wire n_6925;
wire n_17339;
wire n_12334;
wire n_17527;
wire n_11252;
wire n_18358;
wire n_15816;
wire n_14369;
wire n_3062;
wire n_4994;
wire n_7967;
wire n_15998;
wire n_8314;
wire n_384;
wire n_3533;
wire n_7246;
wire n_11086;
wire n_13184;
wire n_3409;
wire n_4381;
wire n_9092;
wire n_4316;
wire n_15900;
wire n_14160;
wire n_4860;
wire n_12994;
wire n_5352;
wire n_10637;
wire n_1157;
wire n_3563;
wire n_20634;
wire n_14637;
wire n_9066;
wire n_763;
wire n_19496;
wire n_12535;
wire n_3442;
wire n_3972;
wire n_14248;
wire n_12582;
wire n_15175;
wire n_1687;
wire n_4934;
wire n_19590;
wire n_2638;
wire n_13988;
wire n_13132;
wire n_1756;
wire n_4350;
wire n_16364;
wire n_18962;
wire n_2340;
wire n_9857;
wire n_8404;
wire n_10056;
wire n_19526;
wire n_6459;
wire n_17300;
wire n_1427;
wire n_14307;
wire n_15678;
wire n_5228;
wire n_1100;
wire n_8606;
wire n_10701;
wire n_7484;
wire n_17397;
wire n_3806;
wire n_9440;
wire n_6753;
wire n_2114;
wire n_5914;
wire n_13879;
wire n_3329;
wire n_11687;
wire n_1175;
wire n_3402;
wire n_1621;
wire n_13522;
wire n_18208;
wire n_6448;
wire n_12524;
wire n_5186;
wire n_19948;
wire n_10454;
wire n_4218;
wire n_9464;
wire n_17532;
wire n_11386;
wire n_4687;
wire n_19033;
wire n_10656;
wire n_394;
wire n_17858;
wire n_3686;
wire n_8741;
wire n_10444;
wire n_11866;
wire n_17020;
wire n_2865;
wire n_17417;
wire n_20387;
wire n_20799;
wire n_13223;
wire n_3259;
wire n_7214;
wire n_11244;
wire n_8806;
wire n_2572;
wire n_1248;
wire n_3677;
wire n_6311;
wire n_8167;
wire n_20722;
wire n_9783;
wire n_4746;
wire n_16957;
wire n_7566;
wire n_18543;
wire n_4215;
wire n_17185;
wire n_12707;
wire n_322;
wire n_17269;
wire n_10546;
wire n_10527;
wire n_9008;
wire n_10143;
wire n_14856;
wire n_8207;
wire n_5344;
wire n_1536;
wire n_3177;
wire n_10186;
wire n_3440;
wire n_20452;
wire n_3658;
wire n_12264;
wire n_16839;
wire n_12464;
wire n_3404;
wire n_3346;
wire n_19497;
wire n_2542;
wire n_10120;
wire n_5892;
wire n_20676;
wire n_20631;
wire n_20056;
wire n_5714;
wire n_9957;
wire n_7975;
wire n_12609;
wire n_17807;
wire n_591;
wire n_10591;
wire n_5634;
wire n_7086;
wire n_7732;
wire n_16332;
wire n_9089;
wire n_8840;
wire n_18327;
wire n_5644;
wire n_20968;
wire n_17767;
wire n_9439;
wire n_19111;
wire n_15405;
wire n_3059;
wire n_15621;
wire n_14773;
wire n_15706;
wire n_16752;
wire n_16180;
wire n_14173;
wire n_19803;
wire n_8179;
wire n_4470;
wire n_10697;
wire n_8111;
wire n_19090;
wire n_17195;
wire n_2868;
wire n_10935;
wire n_13317;
wire n_9631;
wire n_10547;
wire n_18235;
wire n_15432;
wire n_10933;
wire n_19260;
wire n_21098;
wire n_10085;
wire n_19793;
wire n_3328;
wire n_18448;
wire n_9816;
wire n_5343;
wire n_1093;
wire n_8251;
wire n_6518;
wire n_6396;
wire n_14383;
wire n_12195;
wire n_19134;
wire n_14400;
wire n_3469;
wire n_15392;
wire n_14858;
wire n_2835;
wire n_20036;
wire n_5542;
wire n_3099;
wire n_2897;
wire n_8506;
wire n_14725;
wire n_4300;
wire n_18403;
wire n_2024;
wire n_18788;
wire n_10336;
wire n_19297;
wire n_701;
wire n_8635;
wire n_8320;
wire n_9703;
wire n_19052;
wire n_9118;
wire n_16922;
wire n_18237;
wire n_11562;
wire n_3901;
wire n_5180;
wire n_10703;
wire n_11575;
wire n_2973;
wire n_16114;
wire n_16637;
wire n_10198;
wire n_11065;
wire n_2710;
wire n_16393;
wire n_6092;
wire n_12486;
wire n_6462;
wire n_4519;
wire n_18596;
wire n_17849;
wire n_21089;
wire n_5025;
wire n_8872;
wire n_12743;
wire n_240;
wire n_10371;
wire n_3878;
wire n_13578;
wire n_19397;
wire n_4310;
wire n_12610;
wire n_7439;
wire n_17516;
wire n_1902;
wire n_7744;
wire n_2784;
wire n_10346;
wire n_3898;
wire n_20938;
wire n_6702;
wire n_18656;
wire n_10059;
wire n_9961;
wire n_12763;
wire n_16038;
wire n_5924;
wire n_1845;
wire n_20121;
wire n_1533;
wire n_14950;
wire n_7684;
wire n_14834;
wire n_11984;
wire n_1275;
wire n_9692;
wire n_18390;
wire n_13222;
wire n_20008;
wire n_11942;
wire n_11207;
wire n_12280;
wire n_12883;
wire n_19965;
wire n_3824;
wire n_12064;
wire n_10974;
wire n_7313;
wire n_16212;
wire n_5899;
wire n_11482;
wire n_1497;
wire n_15843;
wire n_4479;
wire n_12283;
wire n_6463;
wire n_10351;
wire n_18516;
wire n_4986;
wire n_19400;
wire n_950;
wire n_15789;
wire n_711;
wire n_18421;
wire n_18953;
wire n_11479;
wire n_7036;
wire n_4743;
wire n_9720;
wire n_17206;
wire n_4250;
wire n_8363;
wire n_12208;
wire n_19268;
wire n_19897;
wire n_2188;
wire n_11083;
wire n_14282;
wire n_11907;
wire n_2430;
wire n_12396;
wire n_6084;
wire n_3094;
wire n_741;
wire n_13997;
wire n_13513;
wire n_371;
wire n_5185;
wire n_2964;
wire n_14713;
wire n_308;
wire n_20979;
wire n_865;
wire n_3312;
wire n_1041;
wire n_993;
wire n_3752;
wire n_7380;
wire n_18806;
wire n_12690;
wire n_12813;
wire n_11524;
wire n_9842;
wire n_18375;
wire n_3655;
wire n_5709;
wire n_6277;
wire n_8411;
wire n_8817;
wire n_8461;
wire n_10438;
wire n_3918;
wire n_20706;
wire n_19371;
wire n_11582;
wire n_10946;
wire n_11796;
wire n_9893;
wire n_1310;
wire n_12021;
wire n_5927;
wire n_8691;
wire n_20588;
wire n_9032;
wire n_10275;
wire n_3593;
wire n_14284;
wire n_19029;
wire n_12990;
wire n_1229;
wire n_2582;
wire n_20088;
wire n_6864;
wire n_10204;
wire n_2485;
wire n_18567;
wire n_18894;
wire n_2563;
wire n_19184;
wire n_2875;
wire n_14086;
wire n_1928;
wire n_12672;
wire n_9172;
wire n_14665;
wire n_18614;
wire n_20838;
wire n_12665;
wire n_13719;
wire n_5226;
wire n_7602;
wire n_20037;
wire n_16540;
wire n_9026;
wire n_18136;
wire n_13453;
wire n_7106;
wire n_11700;
wire n_12940;
wire n_7557;
wire n_7408;
wire n_12555;
wire n_16551;
wire n_18727;
wire n_496;
wire n_4335;
wire n_17952;
wire n_6146;
wire n_5677;
wire n_19178;
wire n_4629;
wire n_9515;
wire n_13183;
wire n_5235;
wire n_15650;
wire n_1129;
wire n_1464;
wire n_19206;
wire n_7719;
wire n_3217;
wire n_11996;
wire n_8938;
wire n_20841;
wire n_10455;
wire n_7852;
wire n_12526;
wire n_12456;
wire n_3503;
wire n_20962;
wire n_5979;
wire n_1870;
wire n_10121;
wire n_13809;
wire n_364;
wire n_7582;
wire n_16304;
wire n_5521;
wire n_431;
wire n_2654;
wire n_19529;
wire n_11104;
wire n_2319;
wire n_15234;
wire n_10828;
wire n_13390;
wire n_17160;
wire n_5410;
wire n_1762;
wire n_16591;
wire n_3080;
wire n_17435;
wire n_20887;
wire n_10418;
wire n_18983;
wire n_6917;
wire n_14601;
wire n_11850;
wire n_3428;
wire n_19814;
wire n_2345;
wire n_6612;
wire n_10922;

INVx1_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_113),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_95),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_33),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_70),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_18),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_26),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_52),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_68),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_67),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_47),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_20),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_50),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_92),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_28),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_5),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_8),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_4),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_39),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_16),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_87),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_22),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_43),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_23),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_89),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_127),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_69),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_38),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_48),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_17),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_106),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_94),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_35),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_42),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_90),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_79),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_56),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_15),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_49),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_34),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_71),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_76),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_46),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_77),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_84),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_30),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_72),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_54),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_44),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_31),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_61),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_98),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_119),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_59),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_53),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_123),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_99),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_40),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_100),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_12),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_57),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_45),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_65),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_21),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_93),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_82),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_1),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_19),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_149),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_153),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_145),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_235),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_237),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_158),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_146),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_147),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_263),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_157),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_134),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_169),
.B(n_27),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_140),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_159),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_163),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_138),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_139),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_185),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_264),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_265),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_275),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_205),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_278),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_294),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_281),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_282),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_284),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_175),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_293),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_289),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_292),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_271),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_299),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_266),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_272),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_273),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_265),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_264),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_309),
.A2(n_219),
.B1(n_203),
.B2(n_206),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

AND2x2_ASAP7_75t_SL g359 ( 
.A(n_319),
.B(n_150),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_136),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_192),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_164),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_191),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_344),
.A2(n_202),
.B1(n_253),
.B2(n_252),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_218),
.B(n_248),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_141),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_142),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_322),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

NOR2x1_ASAP7_75t_L g395 ( 
.A(n_324),
.B(n_183),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_304),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_312),
.B(n_184),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_308),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_344),
.A2(n_211),
.B1(n_245),
.B2(n_244),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_321),
.B(n_143),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_341),
.A2(n_186),
.B(n_198),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_312),
.B(n_199),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_308),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_321),
.B(n_144),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_214),
.B1(n_227),
.B2(n_221),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_312),
.B(n_216),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_312),
.B(n_220),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_210),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_304),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_311),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_308),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_308),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_344),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_312),
.B(n_208),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_305),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_308),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_311),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_311),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_308),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_332),
.B(n_213),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_308),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_304),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_312),
.B(n_242),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_328),
.A2(n_207),
.B1(n_259),
.B2(n_258),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_305),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_308),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_308),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_308),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_308),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_311),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_332),
.B(n_201),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_328),
.A2(n_204),
.B1(n_257),
.B2(n_256),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_304),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_311),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_328),
.A2(n_193),
.B1(n_254),
.B2(n_251),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_308),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_308),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_308),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_321),
.B(n_262),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_311),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_308),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_308),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_312),
.B(n_195),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_344),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_308),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_321),
.B(n_250),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_312),
.B(n_239),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_312),
.B(n_233),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_308),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_328),
.A2(n_236),
.B1(n_247),
.B2(n_246),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_308),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_332),
.B(n_188),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_312),
.B(n_187),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_308),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_312),
.B(n_249),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_309),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_331),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_321),
.B(n_182),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_349),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_466),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_356),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_363),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_402),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_370),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_397),
.B(n_398),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_378),
.B(n_388),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_421),
.B(n_243),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_427),
.B(n_181),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_189),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_362),
.B(n_180),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_366),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_379),
.B(n_190),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_386),
.B(n_179),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_360),
.B(n_177),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_350),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_387),
.B(n_353),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_395),
.A2(n_162),
.B(n_229),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_380),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

INVx6_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_197),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_350),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_389),
.B(n_176),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_352),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

NAND2x1_ASAP7_75t_L g514 ( 
.A(n_361),
.B(n_352),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_355),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_391),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_437),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_368),
.B(n_215),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_422),
.B(n_174),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_351),
.A2(n_217),
.B1(n_234),
.B2(n_232),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_417),
.B(n_178),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_439),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_443),
.B(n_171),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_376),
.B(n_168),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_383),
.B(n_424),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_393),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_354),
.B(n_222),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_358),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_390),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_371),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_373),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_374),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_418),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_377),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_382),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_361),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_426),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_384),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_364),
.B(n_406),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_435),
.B(n_166),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_444),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_392),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_385),
.B(n_223),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_403),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_372),
.A2(n_196),
.B(n_229),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_457),
.B(n_161),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_468),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_407),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_359),
.B(n_224),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_412),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_365),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_381),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_453),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_463),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_410),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_441),
.B(n_238),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_456),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_367),
.A2(n_154),
.B(n_231),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_465),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_430),
.Y(n_589)
);

BUFx8_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_405),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_434),
.B(n_228),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_442),
.B(n_226),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_445),
.A2(n_229),
.B(n_196),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_411),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_466),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_385),
.B(n_173),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_349),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_388),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_349),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_466),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_356),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_399),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_356),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_349),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_356),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_399),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_356),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_356),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_399),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_349),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_399),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_399),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_356),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_397),
.B(n_225),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_421),
.B(n_151),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_356),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_349),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_378),
.B(n_238),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_362),
.A2(n_196),
.B1(n_229),
.B2(n_238),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_399),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_421),
.B(n_196),
.Y(n_624)
);

INVxp33_ASAP7_75t_SL g625 ( 
.A(n_353),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_399),
.Y(n_626)
);

BUFx8_ASAP7_75t_L g627 ( 
.A(n_357),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_399),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_399),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_356),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_349),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_399),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_466),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_356),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_356),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_349),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_399),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_356),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_397),
.B(n_229),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_466),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_399),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_349),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_388),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_399),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_466),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_362),
.B(n_196),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_362),
.B(n_62),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_356),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_349),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_399),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_349),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_356),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_466),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_466),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_356),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_388),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_362),
.A2(n_63),
.B1(n_105),
.B2(n_332),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_466),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_399),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_421),
.B(n_332),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_399),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_349),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_362),
.B(n_379),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_356),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_399),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_349),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_362),
.B(n_379),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_356),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_349),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_399),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_349),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_421),
.B(n_454),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_397),
.B(n_305),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_378),
.B(n_388),
.Y(n_675)
);

CKINVDCx8_ASAP7_75t_R g676 ( 
.A(n_357),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_356),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_356),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_399),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_349),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_356),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_362),
.B(n_379),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_399),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_356),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_362),
.B(n_379),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_362),
.B(n_379),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_362),
.B(n_379),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_349),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_349),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_356),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_388),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_385),
.B(n_332),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_395),
.A2(n_345),
.B(n_311),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_466),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_421),
.B(n_454),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_349),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_356),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_421),
.B(n_454),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_356),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_356),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_356),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_SL g702 ( 
.A(n_397),
.B(n_398),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_356),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_349),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_349),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_399),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_349),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_362),
.B(n_379),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_421),
.B(n_454),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_356),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_362),
.B(n_379),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_466),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_366),
.A2(n_380),
.B1(n_401),
.B2(n_400),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_356),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_378),
.B(n_388),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_399),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_356),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_356),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_349),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_399),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_421),
.B(n_332),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_356),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_356),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_356),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_349),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_356),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_421),
.B(n_332),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_356),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_356),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_356),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_356),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_356),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_399),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_349),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_399),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_399),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_356),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_356),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_SL g739 ( 
.A(n_397),
.B(n_398),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_399),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_356),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_349),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_399),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_399),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_356),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_356),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_364),
.A2(n_342),
.B(n_341),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_421),
.B(n_454),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_399),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_399),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_421),
.B(n_332),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_356),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_356),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_385),
.B(n_332),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_349),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_421),
.B(n_454),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_349),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_356),
.Y(n_758)
);

INVxp33_ASAP7_75t_SL g759 ( 
.A(n_353),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_466),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_362),
.B(n_379),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_466),
.A2(n_265),
.B1(n_288),
.B2(n_275),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_356),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_356),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_399),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_356),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_356),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_473),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_470),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_633),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_664),
.B(n_668),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_475),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_476),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_682),
.B(n_685),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_484),
.B(n_675),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_477),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_581),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_472),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_674),
.B(n_616),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_595),
.A2(n_591),
.B1(n_580),
.B2(n_596),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_750),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_472),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_474),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_651),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_686),
.B(n_687),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_611),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_611),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_483),
.B(n_583),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_623),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_604),
.B(n_608),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_708),
.B(n_711),
.Y(n_791)
);

NOR2x1p5_ASAP7_75t_L g792 ( 
.A(n_613),
.B(n_626),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_603),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_623),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_761),
.B(n_584),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_592),
.A2(n_588),
.B1(n_543),
.B2(n_545),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_585),
.B(n_673),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_574),
.A2(n_600),
.B1(n_657),
.B2(n_644),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_605),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_607),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_625),
.B(n_759),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_496),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_628),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_577),
.B(n_559),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_578),
.B(n_702),
.Y(n_805)
);

INVx6_ASAP7_75t_L g806 ( 
.A(n_628),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_695),
.B(n_698),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_632),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_632),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_691),
.B(n_516),
.C(n_692),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_645),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_754),
.B(n_482),
.C(n_598),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_586),
.B(n_579),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_493),
.A2(n_502),
.B1(n_518),
.B2(n_515),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_609),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_610),
.B(n_615),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_660),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_709),
.B(n_756),
.C(n_748),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_661),
.B(n_721),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_503),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_660),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_727),
.B(n_751),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_508),
.Y(n_824)
);

NOR2x1p5_ASAP7_75t_L g825 ( 
.A(n_629),
.B(n_637),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_662),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_519),
.Y(n_827)
);

CKINVDCx6p67_ASAP7_75t_R g828 ( 
.A(n_662),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_713),
.B(n_527),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_666),
.B(n_671),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_618),
.B(n_630),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_533),
.B(n_498),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_R g833 ( 
.A(n_471),
.B(n_597),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_666),
.B(n_671),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_498),
.B(n_509),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_634),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_679),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_635),
.B(n_639),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_679),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_526),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_517),
.B(n_536),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_649),
.B(n_653),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_656),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_762),
.B(n_575),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_665),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_491),
.A2(n_499),
.B1(n_617),
.B2(n_624),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_669),
.B(n_677),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_678),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_683),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_540),
.A2(n_550),
.B1(n_542),
.B2(n_548),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_683),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_490),
.A2(n_492),
.B1(n_589),
.B2(n_497),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_706),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_589),
.A2(n_560),
.B1(n_532),
.B2(n_522),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_602),
.B(n_622),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_599),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_684),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_638),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_690),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_697),
.B(n_699),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_700),
.B(n_701),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_641),
.B(n_654),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_524),
.A2(n_551),
.B1(n_620),
.B2(n_703),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_601),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_720),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_606),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_710),
.B(n_714),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_717),
.B(n_718),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_720),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_612),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_736),
.B(n_743),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_655),
.B(n_712),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_722),
.B(n_723),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_619),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_724),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_726),
.B(n_728),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_743),
.B(n_749),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_631),
.Y(n_881)
);

INVx6_ASAP7_75t_L g882 ( 
.A(n_749),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_729),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_566),
.B(n_541),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_730),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_509),
.B(n_512),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_658),
.B(n_676),
.C(n_538),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_636),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_731),
.B(n_767),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_732),
.B(n_737),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_646),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_738),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_643),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_650),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_741),
.B(n_745),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_752),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_753),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_652),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_642),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_512),
.B(n_531),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_565),
.B(n_573),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_663),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_758),
.B(n_763),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_716),
.B(n_733),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_659),
.B(n_694),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_667),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_764),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_670),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_760),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_766),
.B(n_479),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_672),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_680),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_688),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_531),
.B(n_544),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_735),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_614),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_627),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_740),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_689),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_544),
.B(n_546),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_480),
.B(n_485),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_487),
.B(n_488),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_553),
.B(n_554),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_744),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_489),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_546),
.A2(n_571),
.B1(n_549),
.B2(n_547),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_501),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_504),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_505),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_555),
.B(n_556),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_765),
.B(n_478),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_510),
.B(n_582),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_511),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_481),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_696),
.A2(n_757),
.B1(n_755),
.B2(n_742),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_558),
.B(n_567),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_704),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_481),
.B(n_590),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_513),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_506),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_507),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_570),
.B(n_576),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_705),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_520),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_521),
.B(n_528),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_563),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_707),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_576),
.B(n_582),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_547),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_569),
.B(n_564),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_529),
.B(n_537),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_719),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_725),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_534),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_535),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_539),
.B(n_571),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_734),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_549),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_552),
.Y(n_960)
);

AND3x1_ASAP7_75t_L g961 ( 
.A(n_525),
.B(n_530),
.C(n_561),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_557),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_562),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_587),
.A2(n_523),
.B1(n_572),
.B2(n_593),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_693),
.Y(n_965)
);

OAI22x1_ASAP7_75t_L g966 ( 
.A1(n_486),
.A2(n_495),
.B1(n_621),
.B2(n_647),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_494),
.B(n_514),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_739),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_747),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_640),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_500),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_648),
.B(n_594),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_568),
.B(n_264),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_473),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_470),
.Y(n_976)
);

OAI22xp33_ASAP7_75t_L g977 ( 
.A1(n_595),
.A2(n_421),
.B1(n_454),
.B2(n_674),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_473),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_750),
.B(n_388),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_674),
.B(n_616),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_470),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_674),
.B(n_616),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_496),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_473),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_750),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_472),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_674),
.B(n_616),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_633),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_470),
.Y(n_990)
);

INVx4_ASAP7_75t_SL g991 ( 
.A(n_474),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_484),
.B(n_421),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_473),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_484),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_750),
.Y(n_996)
);

BUFx10_ASAP7_75t_L g997 ( 
.A(n_484),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_472),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_496),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_470),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_473),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_473),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_470),
.Y(n_1003)
);

AO22x2_ASAP7_75t_L g1004 ( 
.A1(n_591),
.A2(n_596),
.B1(n_393),
.B2(n_313),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_750),
.B(n_474),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_473),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_674),
.B(n_616),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_625),
.B(n_264),
.Y(n_1008)
);

AND2x6_ASAP7_75t_L g1009 ( 
.A(n_484),
.B(n_675),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_470),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_473),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_470),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_664),
.B(n_668),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_470),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_470),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_470),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_470),
.Y(n_1017)
);

AND2x6_ASAP7_75t_L g1018 ( 
.A(n_484),
.B(n_675),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_473),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_750),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_473),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_750),
.B(n_474),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_472),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_473),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1025)
);

AO22x2_ASAP7_75t_L g1026 ( 
.A1(n_591),
.A2(n_596),
.B1(n_393),
.B2(n_313),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_473),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_664),
.B(n_668),
.Y(n_1028)
);

AND2x6_ASAP7_75t_L g1029 ( 
.A(n_484),
.B(n_675),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_470),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_472),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_496),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_674),
.B(n_616),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_474),
.B(n_651),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_473),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_473),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_473),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_470),
.Y(n_1039)
);

INVxp33_ASAP7_75t_L g1040 ( 
.A(n_762),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_625),
.B(n_264),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_473),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_473),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_664),
.B(n_668),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_664),
.B(n_668),
.Y(n_1045)
);

BUFx10_ASAP7_75t_L g1046 ( 
.A(n_484),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_472),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_664),
.B(n_668),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_473),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_750),
.B(n_474),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_470),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_470),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_595),
.A2(n_592),
.B1(n_583),
.B2(n_580),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_473),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_473),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_470),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_472),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_473),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_625),
.B(n_264),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_496),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_472),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_470),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_474),
.B(n_651),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_484),
.B(n_421),
.Y(n_1066)
);

BUFx10_ASAP7_75t_L g1067 ( 
.A(n_484),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_473),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_472),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_473),
.Y(n_1070)
);

AO22x2_ASAP7_75t_L g1071 ( 
.A1(n_591),
.A2(n_596),
.B1(n_393),
.B2(n_313),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_471),
.B(n_357),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_470),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_473),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_750),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_473),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_664),
.B(n_668),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_750),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_473),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_673),
.B(n_397),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_750),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_L g1082 ( 
.A(n_664),
.B(n_761),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_674),
.B(n_616),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_474),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_R g1085 ( 
.A(n_633),
.B(n_305),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_473),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_470),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_474),
.Y(n_1088)
);

INVx6_ASAP7_75t_L g1089 ( 
.A(n_472),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_472),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_474),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_664),
.B(n_668),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_473),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_496),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_473),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_470),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_474),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_473),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_750),
.B(n_474),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_664),
.B(n_668),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_750),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_473),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_470),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_592),
.B(n_333),
.C(n_332),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_473),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_473),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_470),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_473),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_592),
.B(n_333),
.C(n_332),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_595),
.A2(n_592),
.B1(n_583),
.B2(n_580),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_472),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_625),
.B(n_264),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_484),
.B(n_421),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_750),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_R g1118 ( 
.A(n_633),
.B(n_305),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_484),
.B(n_421),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_473),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_473),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_470),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_625),
.B(n_264),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_664),
.B(n_668),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_473),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_471),
.B(n_357),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_750),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_625),
.B(n_264),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_470),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_470),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_470),
.Y(n_1131)
);

AND2x6_ASAP7_75t_L g1132 ( 
.A(n_484),
.B(n_675),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_474),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_473),
.Y(n_1134)
);

BUFx4f_ASAP7_75t_L g1135 ( 
.A(n_472),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_592),
.B(n_333),
.C(n_332),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_572),
.A2(n_568),
.B(n_648),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_L g1139 ( 
.A(n_664),
.B(n_761),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_484),
.B(n_421),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_633),
.B(n_466),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_470),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_625),
.B(n_264),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_472),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_664),
.B(n_668),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_470),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_664),
.A2(n_682),
.B1(n_685),
.B2(n_668),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_750),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_473),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_664),
.B(n_668),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_484),
.B(n_421),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_470),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_474),
.B(n_651),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_482),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_470),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_674),
.B(n_616),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_664),
.B(n_668),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_625),
.B(n_264),
.Y(n_1158)
);

INVx4_ASAP7_75t_SL g1159 ( 
.A(n_474),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_472),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_625),
.B(n_264),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_473),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_470),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_484),
.B(n_675),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_750),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_484),
.B(n_421),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_470),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_750),
.Y(n_1168)
);

INVxp33_ASAP7_75t_L g1169 ( 
.A(n_762),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_471),
.B(n_357),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_473),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_595),
.A2(n_592),
.B1(n_583),
.B2(n_580),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_473),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_473),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_664),
.A2(n_682),
.B1(n_685),
.B2(n_668),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_664),
.B(n_668),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_470),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_750),
.Y(n_1178)
);

INVxp33_ASAP7_75t_SL g1179 ( 
.A(n_674),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_484),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_674),
.B(n_616),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_470),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_472),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_474),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_484),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_474),
.Y(n_1186)
);

NOR2x1p5_ASAP7_75t_L g1187 ( 
.A(n_474),
.B(n_378),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_470),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_592),
.B(n_333),
.C(n_332),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_470),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_750),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_591),
.A2(n_596),
.B1(n_583),
.B2(n_592),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_664),
.B(n_668),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_750),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_470),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_472),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_474),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_595),
.A2(n_592),
.B1(n_583),
.B2(n_580),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_470),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_674),
.B(n_616),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_595),
.A2(n_592),
.B1(n_583),
.B2(n_580),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_472),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_625),
.B(n_264),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_473),
.Y(n_1204)
);

NOR2x1p5_ASAP7_75t_L g1205 ( 
.A(n_474),
.B(n_378),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_473),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_473),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_473),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_750),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_769),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_977),
.B(n_1179),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_771),
.B(n_774),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1008),
.B(n_1041),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_785),
.B(n_791),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_841),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_812),
.B(n_1115),
.C(n_1060),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1013),
.B(n_1028),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1123),
.B(n_1128),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1044),
.B(n_1045),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_782),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_768),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_772),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1084),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_853),
.B(n_987),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1143),
.B(n_1161),
.C(n_1158),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1203),
.B(n_1048),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1100),
.B(n_1124),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_SL g1229 ( 
.A(n_947),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_810),
.B(n_798),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1082),
.B(n_1139),
.C(n_1147),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1145),
.B(n_1150),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_979),
.B(n_984),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_775),
.B(n_801),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_999),
.B(n_1033),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_L g1236 ( 
.A(n_853),
.B(n_987),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_773),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1157),
.B(n_1176),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1061),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1193),
.B(n_1175),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_776),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_795),
.B(n_804),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_889),
.B(n_968),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_975),
.B(n_982),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_837),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_994),
.B(n_1025),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1135),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1186),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1054),
.B(n_1112),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1030),
.B(n_1051),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_793),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1064),
.B(n_1101),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1104),
.B(n_1113),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1137),
.B(n_1192),
.Y(n_1254)
);

INVx3_ASAP7_75t_R g1255 ( 
.A(n_918),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1094),
.B(n_1172),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1072),
.B(n_1126),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_799),
.Y(n_1258)
);

OAI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1198),
.A2(n_1201),
.B1(n_1106),
.B2(n_1189),
.C(n_1136),
.Y(n_1259)
);

NAND2xp33_ASAP7_75t_L g1260 ( 
.A(n_889),
.B(n_968),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1111),
.B(n_1154),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_780),
.B(n_813),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_797),
.B(n_777),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_797),
.B(n_777),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_950),
.B(n_992),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_797),
.B(n_777),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_800),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1141),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_816),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_817),
.B(n_831),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_802),
.Y(n_1271)
);

AND2x6_ASAP7_75t_L g1272 ( 
.A(n_970),
.B(n_1066),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_819),
.B(n_1116),
.Y(n_1273)
);

INVxp33_ASAP7_75t_L g1274 ( 
.A(n_1119),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_836),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_991),
.B(n_1159),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_838),
.B(n_842),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_847),
.B(n_861),
.Y(n_1278)
);

INVx8_ASAP7_75t_L g1279 ( 
.A(n_1009),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_950),
.B(n_1140),
.Y(n_1280)
);

INVx5_ASAP7_75t_L g1281 ( 
.A(n_1009),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1151),
.B(n_1166),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_834),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_854),
.B(n_846),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_862),
.B(n_869),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_870),
.B(n_876),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_879),
.B(n_890),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1035),
.Y(n_1288)
);

INVx8_ASAP7_75t_L g1289 ( 
.A(n_1009),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_895),
.B(n_904),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1065),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_865),
.B(n_852),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_884),
.B(n_844),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_807),
.B(n_1170),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_843),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1058),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_828),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_875),
.B(n_859),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_891),
.B(n_1005),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_SL g1300 ( 
.A(n_1153),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_911),
.B(n_922),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_784),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_845),
.Y(n_1303)
);

INVx8_ASAP7_75t_L g1304 ( 
.A(n_1018),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_848),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_923),
.B(n_946),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1058),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1062),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1040),
.B(n_1169),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_779),
.B(n_980),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_L g1311 ( 
.A(n_983),
.B(n_1007),
.C(n_988),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_L g1312 ( 
.A(n_889),
.B(n_967),
.Y(n_1312)
);

AO221x1_ASAP7_75t_L g1313 ( 
.A1(n_966),
.A2(n_1004),
.B1(n_1071),
.B2(n_1026),
.C(n_815),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_857),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_858),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_952),
.B(n_860),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_878),
.B(n_883),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_885),
.B(n_892),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1005),
.B(n_1022),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1018),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_821),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1018),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1029),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_824),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1062),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_896),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1080),
.B(n_1029),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_897),
.B(n_898),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_906),
.B(n_855),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_908),
.B(n_926),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_928),
.B(n_929),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_864),
.B(n_910),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_930),
.B(n_934),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1029),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1034),
.B(n_1083),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1156),
.B(n_1181),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_940),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1022),
.B(n_1050),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1200),
.B(n_1183),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_945),
.B(n_955),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_974),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_827),
.Y(n_1342)
);

OR2x2_ASAP7_75t_SL g1343 ( 
.A(n_770),
.B(n_989),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_820),
.B(n_823),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_978),
.B(n_985),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_993),
.B(n_1001),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1002),
.B(n_1006),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_840),
.Y(n_1349)
);

NOR2xp67_ASAP7_75t_L g1350 ( 
.A(n_1202),
.B(n_781),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1011),
.B(n_1019),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_809),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_778),
.B(n_818),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1021),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1024),
.Y(n_1355)
);

NOR3xp33_ASAP7_75t_L g1356 ( 
.A(n_887),
.B(n_805),
.C(n_829),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_788),
.B(n_942),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1027),
.B(n_1036),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1037),
.B(n_1038),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1042),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_794),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1043),
.B(n_1049),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1132),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_939),
.B(n_787),
.Y(n_1364)
);

NOR3xp33_ASAP7_75t_L g1365 ( 
.A(n_832),
.B(n_919),
.C(n_900),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_806),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1055),
.B(n_1056),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1059),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_933),
.B(n_951),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_856),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_957),
.B(n_1091),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_783),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1374)
);

INVx8_ASAP7_75t_L g1375 ( 
.A(n_1132),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_866),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1079),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1088),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1097),
.B(n_1184),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_778),
.B(n_818),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1086),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_863),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_863),
.B(n_867),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1093),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_963),
.B(n_986),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_882),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1095),
.B(n_1098),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_868),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_996),
.B(n_1020),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1132),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1103),
.Y(n_1391)
);

INVxp33_ASAP7_75t_L g1392 ( 
.A(n_867),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1107),
.B(n_1108),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1110),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1120),
.B(n_1121),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1125),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1162),
.B(n_1171),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_872),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1075),
.B(n_1078),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1204),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1206),
.B(n_1207),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1208),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_877),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1133),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_796),
.B(n_1164),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1081),
.B(n_1117),
.C(n_1102),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_881),
.Y(n_1409)
);

AOI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_943),
.A2(n_932),
.B1(n_902),
.B2(n_937),
.C(n_931),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1127),
.B(n_1148),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1165),
.B(n_1168),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1178),
.B(n_1191),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_888),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_L g1415 ( 
.A(n_1164),
.B(n_1187),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1023),
.B(n_1032),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1164),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1085),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_893),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1089),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1023),
.B(n_1032),
.Y(n_1421)
);

NOR2xp67_ASAP7_75t_L g1422 ( 
.A(n_1194),
.B(n_1209),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1118),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1069),
.B(n_1114),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_958),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1069),
.B(n_1114),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_924),
.B(n_927),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_894),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_899),
.B(n_903),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_L g1430 ( 
.A(n_1197),
.B(n_789),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_835),
.B(n_886),
.C(n_921),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1160),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_907),
.Y(n_1433)
);

NAND2x1_ASAP7_75t_L g1434 ( 
.A(n_965),
.B(n_971),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_973),
.B(n_961),
.C(n_964),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1050),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_909),
.B(n_912),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_913),
.B(n_914),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_920),
.B(n_938),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1099),
.B(n_949),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_960),
.B(n_941),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1144),
.B(n_956),
.Y(n_1442)
);

NOR3xp33_ASAP7_75t_L g1443 ( 
.A(n_901),
.B(n_915),
.C(n_935),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1144),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_944),
.B(n_948),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_962),
.B(n_995),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_953),
.B(n_954),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_997),
.B(n_1046),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1067),
.B(n_1180),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1185),
.B(n_959),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_949),
.B(n_1099),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_833),
.B(n_850),
.C(n_936),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_834),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_786),
.B(n_839),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_976),
.B(n_981),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_990),
.B(n_1000),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1003),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_830),
.B(n_873),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_SL g1459 ( 
.A(n_803),
.B(n_1047),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1010),
.B(n_1052),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_880),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_808),
.B(n_874),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1012),
.B(n_1063),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1014),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1015),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1016),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1017),
.B(n_1146),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_826),
.B(n_1090),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_L g1469 ( 
.A(n_851),
.B(n_998),
.Y(n_1469)
);

BUFx5_ASAP7_75t_L g1470 ( 
.A(n_972),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1031),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_811),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_790),
.B(n_792),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1039),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1205),
.B(n_825),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_814),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1053),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_822),
.B(n_849),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1057),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1073),
.B(n_1131),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1087),
.B(n_1199),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1096),
.B(n_1109),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1105),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_905),
.B(n_871),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1196),
.B(n_916),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_925),
.B(n_1195),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_SL g1487 ( 
.A(n_917),
.B(n_1152),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1122),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1129),
.B(n_1163),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1130),
.B(n_1167),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1142),
.A2(n_1177),
.B1(n_1188),
.B2(n_1182),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1155),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1190),
.B(n_969),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1138),
.B(n_972),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_972),
.B(n_977),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1005),
.B(n_1022),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_771),
.B(n_774),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_768),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_768),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_771),
.B(n_774),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_769),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_977),
.B(n_1179),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_771),
.B(n_774),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_771),
.B(n_774),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1008),
.B(n_264),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_L g1507 ( 
.A(n_771),
.B(n_774),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1084),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_977),
.B(n_1179),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_771),
.B(n_774),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_768),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_769),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1008),
.B(n_264),
.Y(n_1513)
);

INVxp33_ASAP7_75t_L g1514 ( 
.A(n_1141),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_853),
.B(n_397),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_771),
.B(n_774),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1517)
);

INVxp33_ASAP7_75t_L g1518 ( 
.A(n_1141),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_768),
.Y(n_1519)
);

XOR2xp5_ASAP7_75t_L g1520 ( 
.A(n_918),
.B(n_466),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_844),
.A2(n_1040),
.B1(n_1169),
.B2(n_359),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_768),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_977),
.B(n_1179),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_977),
.B(n_1179),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_771),
.B(n_774),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1005),
.B(n_1022),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_SL g1527 ( 
.A(n_1106),
.B(n_378),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_771),
.B(n_774),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_769),
.Y(n_1529)
);

BUFx8_ASAP7_75t_L g1530 ( 
.A(n_918),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_977),
.B(n_1179),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_771),
.B(n_774),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_769),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_768),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1008),
.A2(n_1060),
.B(n_1041),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_769),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_775),
.B(n_801),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_769),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_977),
.B(n_1179),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_771),
.B(n_774),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1008),
.B(n_264),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_977),
.B(n_1179),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_782),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_768),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1008),
.B(n_264),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_769),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_768),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1008),
.B(n_264),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_771),
.B(n_774),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_768),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_SL g1551 ( 
.A(n_947),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_771),
.B(n_774),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_768),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_771),
.A2(n_774),
.B1(n_791),
.B2(n_785),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_768),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_769),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_977),
.B(n_1179),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1008),
.B(n_264),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_775),
.B(n_801),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_977),
.B(n_1179),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_782),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_782),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_768),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_977),
.B(n_1179),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_771),
.B(n_774),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_782),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1084),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_768),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1085),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_771),
.B(n_774),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1008),
.B(n_750),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_771),
.B(n_774),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_775),
.B(n_801),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_977),
.B(n_1179),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1008),
.B(n_264),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_768),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_853),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_771),
.B(n_774),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1008),
.B(n_264),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1008),
.B(n_264),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_769),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_771),
.B(n_774),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_768),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_768),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_771),
.B(n_774),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_977),
.B(n_1179),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1008),
.A2(n_1060),
.B1(n_1115),
.B2(n_1041),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_977),
.B(n_1179),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_769),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_L g1590 ( 
.A(n_853),
.B(n_397),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_769),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1008),
.B(n_264),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_768),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_771),
.B(n_774),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1084),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_782),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_768),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1008),
.B(n_264),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_768),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1008),
.B(n_264),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_771),
.B(n_397),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1008),
.B(n_264),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1008),
.B(n_264),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1008),
.B(n_264),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_841),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_768),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_853),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_768),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_771),
.B(n_774),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_768),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_771),
.B(n_774),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_782),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_775),
.B(n_801),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_841),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_771),
.B(n_774),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_769),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1084),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1008),
.B(n_264),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_977),
.B(n_1179),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_769),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1008),
.B(n_264),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_769),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_768),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_775),
.B(n_801),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_771),
.A2(n_785),
.B(n_791),
.C(n_774),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_1141),
.Y(n_1629)
);

NOR2x1p5_ASAP7_75t_L g1630 ( 
.A(n_828),
.B(n_378),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_771),
.B(n_774),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_771),
.B(n_774),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_769),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_771),
.B(n_774),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_984),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_977),
.B(n_1179),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_769),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_771),
.B(n_774),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_769),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_L g1640 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_L g1641 ( 
.A(n_771),
.B(n_774),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1008),
.B(n_264),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_769),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1008),
.B(n_264),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1085),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_782),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1008),
.B(n_264),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1035),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_771),
.B(n_774),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_771),
.B(n_774),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_771),
.B(n_774),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_775),
.B(n_801),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_SL g1653 ( 
.A(n_947),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_768),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_SL g1655 ( 
.A(n_947),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1008),
.B(n_264),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_769),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_775),
.B(n_801),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_768),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_768),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_769),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1084),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1141),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1008),
.B(n_264),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_771),
.B(n_774),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_768),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_768),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_769),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_SL g1670 ( 
.A(n_771),
.B(n_397),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_771),
.B(n_774),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1085),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_775),
.B(n_801),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_782),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_771),
.B(n_774),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_769),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_769),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_771),
.B(n_774),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1008),
.B(n_264),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1141),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1008),
.B(n_264),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_769),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_768),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_768),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_841),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_977),
.B(n_1179),
.Y(n_1686)
);

NAND2xp33_ASAP7_75t_L g1687 ( 
.A(n_771),
.B(n_774),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_841),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_768),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_768),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_782),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_L g1692 ( 
.A(n_771),
.B(n_774),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_768),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1008),
.B(n_264),
.Y(n_1694)
);

BUFx8_ASAP7_75t_L g1695 ( 
.A(n_918),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_768),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_769),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_768),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1082),
.A2(n_1139),
.B(n_774),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_768),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1008),
.B(n_264),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1008),
.B(n_264),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_769),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1008),
.B(n_264),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_782),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_853),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_977),
.B(n_1179),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1084),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_977),
.B(n_1179),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_841),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1008),
.B(n_264),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_768),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_769),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_977),
.B(n_1179),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1008),
.B(n_264),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1141),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_768),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_768),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_768),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_841),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_769),
.Y(n_1725)
);

NOR2xp67_ASAP7_75t_L g1726 ( 
.A(n_853),
.B(n_397),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_771),
.B(n_774),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_771),
.B(n_774),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_775),
.B(n_801),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_782),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1084),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_977),
.B(n_1179),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1008),
.B(n_264),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_771),
.B(n_774),
.Y(n_1734)
);

NOR2xp67_ASAP7_75t_L g1735 ( 
.A(n_853),
.B(n_397),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_771),
.B(n_774),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_771),
.B(n_774),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_768),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_L g1739 ( 
.A(n_771),
.B(n_774),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_984),
.B(n_357),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_768),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_L g1742 ( 
.A(n_771),
.B(n_774),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_977),
.B(n_1179),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_841),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_SL g1745 ( 
.A(n_947),
.Y(n_1745)
);

BUFx5_ASAP7_75t_L g1746 ( 
.A(n_889),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1008),
.A2(n_1115),
.B1(n_1123),
.B2(n_1060),
.C(n_1041),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1035),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1008),
.B(n_264),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_768),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_771),
.A2(n_785),
.B(n_791),
.C(n_774),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_771),
.B(n_774),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_768),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1008),
.B(n_264),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1008),
.B(n_264),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1084),
.Y(n_1756)
);

BUFx5_ASAP7_75t_L g1757 ( 
.A(n_889),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_768),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_977),
.B(n_1179),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_769),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1008),
.B(n_264),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1005),
.B(n_1022),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1084),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_775),
.B(n_801),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_771),
.B(n_774),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_841),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_L g1768 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1008),
.B(n_264),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_977),
.B(n_1179),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_769),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_768),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_769),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_771),
.B(n_774),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_977),
.B(n_1179),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_768),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_L g1777 ( 
.A(n_771),
.B(n_774),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1008),
.B(n_264),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_769),
.Y(n_1779)
);

INVxp33_ASAP7_75t_L g1780 ( 
.A(n_1141),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_841),
.Y(n_1781)
);

NOR3xp33_ASAP7_75t_L g1782 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_769),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_L g1784 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_977),
.B(n_1179),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_977),
.B(n_1179),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1008),
.B(n_264),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_L g1788 ( 
.A(n_771),
.B(n_774),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_977),
.B(n_1179),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_771),
.B(n_774),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_769),
.Y(n_1791)
);

NAND2xp33_ASAP7_75t_L g1792 ( 
.A(n_771),
.B(n_774),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_771),
.B(n_774),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_977),
.B(n_1179),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1008),
.B(n_264),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_768),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_768),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_771),
.B(n_774),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_768),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_775),
.B(n_801),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_771),
.B(n_774),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_768),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_771),
.B(n_774),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_771),
.B(n_774),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1008),
.B(n_264),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_768),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_768),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_769),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_771),
.B(n_774),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_768),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1008),
.B(n_264),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_977),
.B(n_1179),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_977),
.B(n_1179),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_984),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_977),
.B(n_1179),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_771),
.B(n_774),
.Y(n_1818)
);

NAND2xp33_ASAP7_75t_L g1819 ( 
.A(n_771),
.B(n_774),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_771),
.B(n_774),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_769),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_768),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1008),
.B(n_264),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_771),
.B(n_774),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1008),
.B(n_264),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_768),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_768),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1084),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_768),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_771),
.B(n_774),
.Y(n_1830)
);

NAND2xp33_ASAP7_75t_L g1831 ( 
.A(n_771),
.B(n_774),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_771),
.B(n_774),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1005),
.B(n_1022),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_768),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_L g1836 ( 
.A(n_812),
.B(n_307),
.C(n_305),
.Y(n_1836)
);

NAND2xp33_ASAP7_75t_L g1837 ( 
.A(n_771),
.B(n_774),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1008),
.B(n_264),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_977),
.B(n_1179),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_977),
.B(n_1179),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_771),
.B(n_774),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1008),
.B(n_264),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_769),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1008),
.A2(n_1060),
.B1(n_1115),
.B2(n_1041),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1084),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_769),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_977),
.B(n_1179),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_SL g1849 ( 
.A(n_947),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1084),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1008),
.B(n_264),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1085),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_L g1853 ( 
.A(n_771),
.B(n_774),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_841),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_771),
.B(n_774),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_768),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_771),
.B(n_774),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_771),
.B(n_774),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_977),
.B(n_1179),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_771),
.B(n_774),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_782),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_771),
.A2(n_785),
.B(n_791),
.C(n_774),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_768),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_768),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_984),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_768),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_771),
.B(n_774),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_771),
.B(n_774),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_771),
.B(n_774),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_984),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_771),
.B(n_774),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1035),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1141),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1084),
.Y(n_1874)
);

NAND2xp33_ASAP7_75t_L g1875 ( 
.A(n_771),
.B(n_774),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1008),
.B(n_264),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_984),
.B(n_357),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_768),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1085),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_768),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1008),
.B(n_264),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_771),
.B(n_774),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_977),
.B(n_1179),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_771),
.B(n_774),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_771),
.B(n_774),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_782),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_841),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_775),
.B(n_801),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_771),
.B(n_774),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1008),
.B(n_264),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_782),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1008),
.A2(n_1060),
.B1(n_1115),
.B2(n_1041),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1008),
.B(n_264),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_977),
.B(n_1179),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_775),
.B(n_801),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_SL g1896 ( 
.A(n_947),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_841),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_775),
.B(n_801),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_782),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_768),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_977),
.B(n_1179),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_771),
.B(n_774),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1008),
.B(n_1060),
.C(n_1041),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1084),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1084),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_771),
.B(n_774),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_771),
.B(n_774),
.Y(n_1908)
);

AO221x1_ASAP7_75t_L g1909 ( 
.A1(n_977),
.A2(n_524),
.B1(n_351),
.B2(n_966),
.C(n_1147),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_771),
.B(n_774),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1008),
.B(n_264),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_844),
.A2(n_1040),
.B1(n_1169),
.B2(n_359),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1008),
.B(n_264),
.Y(n_1913)
);

AND2x2_ASAP7_75t_SL g1914 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1226),
.B(n_1212),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1210),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1214),
.B(n_1219),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1554),
.B(n_1344),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1329),
.B(n_1240),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1281),
.B(n_1319),
.Y(n_1920)
);

INVx2_ASAP7_75t_SL g1921 ( 
.A(n_1220),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1293),
.B(n_1617),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1213),
.B(n_1218),
.Y(n_1923)
);

INVxp33_ASAP7_75t_L g1924 ( 
.A(n_1740),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1245),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1281),
.B(n_1338),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1227),
.B(n_1228),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1232),
.B(n_1238),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1221),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1216),
.B(n_1587),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_SL g1931 ( 
.A1(n_1517),
.A2(n_1603),
.B(n_1720),
.C(n_1640),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1691),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1535),
.B(n_1845),
.Y(n_1933)
);

OAI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1231),
.A2(n_1751),
.B(n_1628),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1892),
.B(n_1215),
.Y(n_1935)
);

OAI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1497),
.A2(n_1500),
.B1(n_1504),
.B2(n_1503),
.Y(n_1936)
);

OAI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1510),
.A2(n_1516),
.B1(n_1528),
.B2(n_1525),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1608),
.B(n_1685),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1222),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1356),
.B(n_1862),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1747),
.B(n_1688),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1237),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1897),
.B(n_1234),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1257),
.B(n_1298),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1241),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1506),
.A2(n_1513),
.B1(n_1545),
.B2(n_1541),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1711),
.B(n_1724),
.Y(n_1948)
);

NOR2xp67_ASAP7_75t_SL g1949 ( 
.A(n_1891),
.B(n_1899),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1549),
.B(n_1552),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1744),
.B(n_1767),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1244),
.A2(n_1250),
.B1(n_1252),
.B2(n_1246),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1781),
.B(n_1854),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1565),
.B(n_1570),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1225),
.A2(n_1578),
.B1(n_1582),
.B2(n_1572),
.Y(n_1955)
);

NOR2xp67_ASAP7_75t_L g1956 ( 
.A(n_1418),
.B(n_1423),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1585),
.B(n_1594),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1887),
.B(n_1230),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1612),
.B(n_1614),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1618),
.B(n_1631),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1279),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1537),
.B(n_1559),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1573),
.B(n_1616),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1632),
.B(n_1634),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1253),
.A2(n_1254),
.B1(n_1909),
.B2(n_1284),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1308),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1638),
.B(n_1649),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1650),
.B(n_1651),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1666),
.B(n_1671),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1675),
.B(n_1678),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1727),
.B(n_1728),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1251),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1734),
.B(n_1736),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1627),
.B(n_1652),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1332),
.B(n_1737),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1521),
.A2(n_1912),
.B1(n_1262),
.B2(n_1313),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1258),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1752),
.B(n_1765),
.Y(n_1978)
);

NOR2x2_ASAP7_75t_L g1979 ( 
.A(n_1496),
.B(n_1526),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1292),
.A2(n_1309),
.B1(n_1502),
.B2(n_1211),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1658),
.B(n_1673),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1774),
.B(n_1790),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1793),
.B(n_1798),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1267),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1802),
.B(n_1805),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1806),
.B(n_1811),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1239),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1818),
.B(n_1820),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1824),
.B(n_1830),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1269),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1832),
.B(n_1842),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1855),
.B(n_1857),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1858),
.B(n_1860),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1729),
.B(n_1764),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1275),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1867),
.B(n_1868),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1869),
.B(n_1871),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1877),
.B(n_1635),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1295),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1321),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1882),
.B(n_1884),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1308),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1279),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1816),
.B(n_1865),
.Y(n_2004)
);

OA22x2_ASAP7_75t_L g2005 ( 
.A1(n_1407),
.A2(n_1256),
.B1(n_1523),
.B2(n_1509),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1524),
.A2(n_1539),
.B1(n_1542),
.B2(n_1531),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1217),
.A2(n_1641),
.B(n_1507),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1885),
.B(n_1889),
.Y(n_2008)
);

NOR3xp33_ASAP7_75t_L g2009 ( 
.A(n_1722),
.B(n_1782),
.C(n_1768),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1903),
.B(n_1907),
.Y(n_2010)
);

NOR2xp67_ASAP7_75t_L g2011 ( 
.A(n_1281),
.B(n_1577),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1908),
.B(n_1910),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1242),
.B(n_1687),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1303),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1410),
.B(n_1766),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1307),
.Y(n_2016)
);

OAI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1548),
.A2(n_1575),
.B(n_1558),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1784),
.A2(n_1901),
.B1(n_1904),
.B2(n_1840),
.Y(n_2018)
);

A2O1A1Ixp33_ASAP7_75t_L g2019 ( 
.A1(n_1692),
.A2(n_1739),
.B(n_1777),
.C(n_1742),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1324),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1320),
.B(n_1323),
.Y(n_2021)
);

NAND2x1p5_ASAP7_75t_L g2022 ( 
.A(n_1339),
.B(n_1557),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1342),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1579),
.A2(n_1580),
.B1(n_1598),
.B2(n_1592),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1305),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1261),
.B(n_1270),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1289),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1788),
.B(n_1792),
.Y(n_2028)
);

NOR2x2_ASAP7_75t_L g2029 ( 
.A(n_1496),
.B(n_1526),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1801),
.B(n_1888),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1560),
.A2(n_1564),
.B1(n_1586),
.B2(n_1574),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1277),
.B(n_1278),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1349),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1819),
.B(n_1831),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1837),
.B(n_1853),
.Y(n_2035)
);

NAND2xp33_ASAP7_75t_L g2036 ( 
.A(n_1746),
.B(n_1757),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1875),
.B(n_1601),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1630),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1588),
.A2(n_1636),
.B1(n_1686),
.B2(n_1622),
.Y(n_2039)
);

A2O1A1Ixp33_ASAP7_75t_L g2040 ( 
.A1(n_1259),
.A2(n_1605),
.B(n_1607),
.C(n_1606),
.Y(n_2040)
);

AND2x2_ASAP7_75t_SL g2041 ( 
.A(n_1260),
.B(n_1327),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1708),
.A2(n_1715),
.B1(n_1732),
.B2(n_1710),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1699),
.B(n_1746),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1913),
.B(n_1621),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1569),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_1386),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1911),
.B(n_1624),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1314),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1315),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1361),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1289),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1642),
.A2(n_1644),
.B1(n_1656),
.B2(n_1647),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1665),
.B(n_1679),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1681),
.A2(n_1694),
.B1(n_1703),
.B2(n_1702),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_SL g2055 ( 
.A1(n_1705),
.A2(n_1717),
.B1(n_1733),
.B2(n_1712),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_SL g2056 ( 
.A1(n_1749),
.A2(n_1755),
.B1(n_1761),
.B2(n_1754),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1743),
.B(n_1759),
.Y(n_2057)
);

NOR2x2_ASAP7_75t_L g2058 ( 
.A(n_1762),
.B(n_1834),
.Y(n_2058)
);

NOR2xp67_ASAP7_75t_L g2059 ( 
.A(n_1610),
.B(n_1707),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1370),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1770),
.B(n_1775),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1785),
.B(n_1786),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1769),
.B(n_1778),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1285),
.A2(n_1287),
.B1(n_1290),
.B2(n_1286),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_L g2065 ( 
.A(n_1787),
.B(n_1807),
.C(n_1795),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1789),
.B(n_1794),
.Y(n_2066)
);

INVx8_ASAP7_75t_L g2067 ( 
.A(n_1304),
.Y(n_2067)
);

AND2x6_ASAP7_75t_L g2068 ( 
.A(n_1263),
.B(n_1264),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1301),
.A2(n_1306),
.B(n_1494),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1326),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1813),
.B(n_1823),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1571),
.B(n_1379),
.Y(n_2072)
);

AND2x4_ASAP7_75t_SL g2073 ( 
.A(n_1297),
.B(n_1276),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1825),
.A2(n_1838),
.B1(n_1851),
.B2(n_1843),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1876),
.B(n_1881),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1814),
.A2(n_1815),
.B1(n_1839),
.B2(n_1817),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1890),
.B(n_1893),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_1223),
.Y(n_2078)
);

A2O1A1Ixp33_ASAP7_75t_L g2079 ( 
.A1(n_1335),
.A2(n_1311),
.B(n_1435),
.C(n_1495),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_1223),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1841),
.B(n_1848),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1376),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1304),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_L g2084 ( 
.A(n_1859),
.B(n_1894),
.C(n_1883),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1895),
.B(n_1898),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1282),
.B(n_1316),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1902),
.B(n_1372),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1337),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1294),
.B(n_1272),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1505),
.A2(n_1600),
.B1(n_1662),
.B2(n_1604),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1272),
.B(n_1369),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1341),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1272),
.B(n_1870),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1354),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1274),
.B(n_1427),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_SL g2096 ( 
.A1(n_1527),
.A2(n_1365),
.B(n_1400),
.C(n_1389),
.Y(n_2096)
);

INVx4_ASAP7_75t_L g2097 ( 
.A(n_1375),
.Y(n_2097)
);

BUFx4f_ASAP7_75t_L g2098 ( 
.A(n_1375),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1746),
.B(n_1757),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1355),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1271),
.B(n_1273),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1388),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1746),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1399),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1494),
.A2(n_1312),
.B(n_1434),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_1310),
.B(n_1336),
.Y(n_2106)
);

AND2x6_ASAP7_75t_SL g2107 ( 
.A(n_1473),
.B(n_1762),
.Y(n_2107)
);

INVx4_ASAP7_75t_L g2108 ( 
.A(n_1248),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1317),
.B(n_1318),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1757),
.B(n_1602),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1328),
.B(n_1330),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1360),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1233),
.B(n_1235),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1368),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1377),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1331),
.B(n_1333),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_1248),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1340),
.B(n_1345),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_1415),
.A2(n_1664),
.B1(n_1873),
.B2(n_1475),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1757),
.B(n_1645),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_1508),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1346),
.B(n_1348),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1351),
.B(n_1358),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1359),
.B(n_1362),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1405),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1367),
.B(n_1371),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_SL g2127 ( 
.A(n_1672),
.B(n_1852),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1879),
.B(n_1357),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1374),
.B(n_1387),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1701),
.B(n_1716),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1393),
.B(n_1395),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1409),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1414),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1381),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_1384),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1419),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1800),
.B(n_1804),
.Y(n_2137)
);

BUFx5_ASAP7_75t_L g2138 ( 
.A(n_1391),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1833),
.B(n_1836),
.Y(n_2139)
);

A2O1A1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_1670),
.A2(n_1398),
.B(n_1401),
.C(n_1397),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1403),
.B(n_1648),
.Y(n_2141)
);

AND2x6_ASAP7_75t_SL g2142 ( 
.A(n_1834),
.B(n_1484),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1748),
.B(n_1872),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1428),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1394),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1396),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1461),
.B(n_1402),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1364),
.A2(n_1451),
.B1(n_1459),
.B2(n_1487),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1404),
.A2(n_1499),
.B(n_1498),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1511),
.B(n_1519),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1453),
.B(n_1283),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_1508),
.Y(n_2152)
);

BUFx8_ASAP7_75t_L g2153 ( 
.A(n_1229),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1551),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1522),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1534),
.B(n_1544),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_SL g2157 ( 
.A1(n_1255),
.A2(n_1343),
.B1(n_1520),
.B2(n_1518),
.Y(n_2157)
);

NOR2xp67_ASAP7_75t_L g2158 ( 
.A(n_1366),
.B(n_1420),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1433),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_SL g2160 ( 
.A(n_1247),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1547),
.B(n_1550),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1567),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1514),
.B(n_1629),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1299),
.B(n_1266),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1553),
.B(n_1555),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1288),
.B(n_1291),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1268),
.B(n_1680),
.Y(n_2167)
);

AOI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_1452),
.A2(n_1425),
.B1(n_1568),
.B2(n_1563),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1653),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1576),
.B(n_1583),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1436),
.B(n_1224),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1464),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1584),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1236),
.B(n_1440),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_1567),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1593),
.B(n_1597),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1599),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1472),
.B(n_1382),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1609),
.B(n_1611),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1613),
.B(n_1626),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1595),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1654),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_1441),
.A2(n_1334),
.B1(n_1417),
.B2(n_1363),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1466),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1659),
.B(n_1660),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1479),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_1667),
.A2(n_1683),
.B(n_1668),
.Y(n_2187)
);

OAI22xp33_ASAP7_75t_SL g2188 ( 
.A1(n_1684),
.A2(n_1797),
.B1(n_1721),
.B2(n_1900),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1483),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1302),
.A2(n_1413),
.B1(n_1412),
.B2(n_1411),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1382),
.B(n_1444),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1718),
.B(n_1780),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1689),
.B(n_1690),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_1693),
.B(n_1696),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_1458),
.B(n_1392),
.Y(n_2195)
);

INVx4_ASAP7_75t_L g2196 ( 
.A(n_1595),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1698),
.B(n_1700),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1488),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1501),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1713),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1719),
.B(n_1723),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_1738),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_1741),
.B(n_1750),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1444),
.B(n_1753),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_1758),
.A2(n_1812),
.B1(n_1772),
.B2(n_1880),
.Y(n_2205)
);

NOR2xp67_ASAP7_75t_L g2206 ( 
.A(n_1543),
.B(n_1561),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1776),
.B(n_1796),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1799),
.B(n_1803),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1808),
.A2(n_1863),
.B1(n_1856),
.B2(n_1826),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1431),
.A2(n_1300),
.B1(n_1886),
.B2(n_1861),
.Y(n_2210)
);

INVx2_ASAP7_75t_SL g2211 ( 
.A(n_1620),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1512),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_SL g2213 ( 
.A(n_1322),
.B(n_1390),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_1809),
.A2(n_1829),
.B1(n_1878),
.B2(n_1866),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1432),
.B(n_1265),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_1486),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1822),
.B(n_1827),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1835),
.B(n_1864),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1385),
.B(n_1515),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1655),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1489),
.B(n_1462),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_1280),
.B(n_1373),
.Y(n_2222)
);

NOR3xp33_ASAP7_75t_L g2223 ( 
.A(n_1442),
.B(n_1408),
.C(n_1443),
.Y(n_2223)
);

NAND2x1_ASAP7_75t_L g2224 ( 
.A(n_1491),
.B(n_1493),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1529),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1478),
.B(n_1476),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1378),
.B(n_1406),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1533),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1350),
.B(n_1450),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_1590),
.B(n_1726),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_1457),
.B(n_1465),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1422),
.A2(n_1735),
.B1(n_1446),
.B2(n_1352),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1353),
.B(n_1380),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1471),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1474),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1485),
.B(n_1430),
.Y(n_2236)
);

A2O1A1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_1477),
.A2(n_1492),
.B(n_1426),
.C(n_1424),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_1429),
.A2(n_1490),
.B(n_1482),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1536),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_SL g2240 ( 
.A(n_1562),
.B(n_1566),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1468),
.B(n_1469),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1596),
.B(n_1615),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1538),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1646),
.B(n_1674),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1706),
.B(n_1730),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_1546),
.A2(n_1657),
.B1(n_1847),
.B2(n_1844),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1556),
.B(n_1581),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1589),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_1437),
.A2(n_1481),
.B(n_1480),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1745),
.Y(n_2250)
);

NAND2xp33_ASAP7_75t_L g2251 ( 
.A(n_1470),
.B(n_1296),
.Y(n_2251)
);

INVxp67_ASAP7_75t_SL g2252 ( 
.A(n_1470),
.Y(n_2252)
);

BUFx8_ASAP7_75t_L g2253 ( 
.A(n_1849),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1620),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1591),
.B(n_1669),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1383),
.B(n_1416),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_1530),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1619),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1623),
.Y(n_2259)
);

OAI221xp5_ASAP7_75t_L g2260 ( 
.A1(n_1325),
.A2(n_1347),
.B1(n_1454),
.B2(n_1421),
.C(n_1449),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1663),
.B(n_1906),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1625),
.Y(n_2262)
);

NAND2x1_ASAP7_75t_L g2263 ( 
.A(n_1633),
.B(n_1704),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1896),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1637),
.B(n_1661),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1639),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_1448),
.A2(n_1906),
.B1(n_1905),
.B2(n_1874),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1643),
.B(n_1714),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1663),
.B(n_1905),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1676),
.B(n_1725),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1677),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_1709),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1682),
.B(n_1821),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_1874),
.B(n_1731),
.Y(n_2274)
);

OAI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_1438),
.A2(n_1439),
.B1(n_1445),
.B2(n_1447),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_1455),
.A2(n_1456),
.B(n_1460),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1709),
.B(n_1850),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1697),
.B(n_1771),
.Y(n_2278)
);

INVx4_ASAP7_75t_L g2279 ( 
.A(n_1731),
.Y(n_2279)
);

AOI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_1760),
.A2(n_1779),
.B1(n_1810),
.B2(n_1791),
.Y(n_2280)
);

INVx5_ASAP7_75t_L g2281 ( 
.A(n_1850),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1773),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1695),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1756),
.B(n_1846),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_1756),
.A2(n_1763),
.B1(n_1828),
.B2(n_1846),
.Y(n_2285)
);

O2A1O1Ixp5_ASAP7_75t_L g2286 ( 
.A1(n_1783),
.A2(n_1463),
.B(n_1467),
.C(n_1470),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1763),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1828),
.B(n_1470),
.Y(n_2288)
);

AOI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1221),
.Y(n_2290)
);

AO22x1_ASAP7_75t_L g2291 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_844),
.B2(n_1506),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1569),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2294)
);

OAI22x1_ASAP7_75t_R g2295 ( 
.A1(n_1664),
.A2(n_466),
.B1(n_633),
.B2(n_1873),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1221),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1210),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1221),
.Y(n_2303)
);

OAI221xp5_ASAP7_75t_L g2304 ( 
.A1(n_1747),
.A2(n_1845),
.B1(n_1892),
.B2(n_1587),
.C(n_1535),
.Y(n_2304)
);

BUFx12f_ASAP7_75t_L g2305 ( 
.A(n_1530),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1210),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2311)
);

NOR2xp67_ASAP7_75t_L g2312 ( 
.A(n_1418),
.B(n_750),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_1281),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1281),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_L g2326 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2327)
);

A2O1A1Ixp33_ASAP7_75t_SL g2328 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1603),
.C(n_1517),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1279),
.Y(n_2330)
);

AO22x1_ASAP7_75t_L g2331 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_844),
.B2(n_1506),
.Y(n_2331)
);

NAND3xp33_ASAP7_75t_L g2332 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_1279),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_1747),
.B(n_1845),
.C(n_1587),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2339)
);

AOI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_L g2342 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_1239),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1210),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_1239),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1221),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2348)
);

BUFx8_ASAP7_75t_SL g2349 ( 
.A(n_1664),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1221),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2354)
);

NOR2xp67_ASAP7_75t_L g2355 ( 
.A(n_1418),
.B(n_750),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_1271),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2358)
);

AOI22xp33_ASAP7_75t_L g2359 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_1281),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1221),
.Y(n_2361)
);

O2A1O1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1535),
.C(n_1226),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_1271),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1210),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_1271),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_1569),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1210),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2378)
);

AOI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1210),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1210),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1221),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1221),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2391)
);

INVx3_ASAP7_75t_L g2392 ( 
.A(n_1279),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1221),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1221),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1210),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2398)
);

INVx2_ASAP7_75t_SL g2399 ( 
.A(n_1220),
.Y(n_2399)
);

NAND2xp33_ASAP7_75t_L g2400 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1210),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1221),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1221),
.Y(n_2408)
);

NOR2x1_ASAP7_75t_R g2409 ( 
.A(n_1220),
.B(n_633),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1221),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1221),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1210),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1221),
.Y(n_2415)
);

NAND2xp33_ASAP7_75t_L g2416 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2416)
);

AND2x6_ASAP7_75t_SL g2417 ( 
.A(n_1213),
.B(n_1218),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1210),
.Y(n_2418)
);

OR2x6_ASAP7_75t_L g2419 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2419)
);

NOR3xp33_ASAP7_75t_L g2420 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1221),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_1220),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_SL g2425 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_1569),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1221),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2429)
);

A2O1A1Ixp33_ASAP7_75t_SL g2430 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1603),
.C(n_1517),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2434)
);

AOI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2438)
);

INVx8_ASAP7_75t_L g2439 ( 
.A(n_1279),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1210),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2447)
);

HB1xp67_ASAP7_75t_L g2448 ( 
.A(n_1271),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1221),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_1361),
.Y(n_2452)
);

AOI221xp5_ASAP7_75t_L g2453 ( 
.A1(n_1226),
.A2(n_1747),
.B1(n_1213),
.B2(n_1218),
.C(n_1513),
.Y(n_2453)
);

OAI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_1226),
.A2(n_1231),
.B(n_1344),
.Y(n_2454)
);

A2O1A1Ixp33_ASAP7_75t_L g2455 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1249),
.C(n_1628),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_1569),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_1210),
.Y(n_2463)
);

NOR2x1p5_ASAP7_75t_L g2464 ( 
.A(n_1220),
.B(n_474),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_1220),
.Y(n_2465)
);

INVx4_ASAP7_75t_L g2466 ( 
.A(n_1308),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2467)
);

AOI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2468)
);

AOI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_1308),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_1220),
.Y(n_2471)
);

NOR2xp67_ASAP7_75t_L g2472 ( 
.A(n_1418),
.B(n_750),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_1281),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_1210),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_1221),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1221),
.Y(n_2481)
);

AND2x6_ASAP7_75t_SL g2482 ( 
.A(n_1213),
.B(n_1218),
.Y(n_2482)
);

BUFx8_ASAP7_75t_L g2483 ( 
.A(n_1229),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2484)
);

BUFx2_ASAP7_75t_L g2485 ( 
.A(n_1361),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1221),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1221),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_1220),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_1220),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_1210),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2499)
);

XOR2xp5_ASAP7_75t_L g2500 ( 
.A(n_1520),
.B(n_466),
.Y(n_2500)
);

NOR3xp33_ASAP7_75t_L g2501 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2503)
);

NAND2x1p5_ASAP7_75t_L g2504 ( 
.A(n_1281),
.B(n_950),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2505)
);

OR2x2_ASAP7_75t_SL g2506 ( 
.A(n_1225),
.B(n_1106),
.Y(n_2506)
);

NAND2x1p5_ASAP7_75t_L g2507 ( 
.A(n_1281),
.B(n_950),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1221),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2509)
);

OAI22xp33_ASAP7_75t_L g2510 ( 
.A1(n_1240),
.A2(n_1587),
.B1(n_1892),
.B2(n_1845),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_1210),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1221),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1221),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1221),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2518)
);

NOR2xp33_ASAP7_75t_SL g2519 ( 
.A(n_1569),
.B(n_466),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2520)
);

OR2x6_ASAP7_75t_L g2521 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_1279),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1221),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_L g2527 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_1210),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_1220),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1221),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2532)
);

NOR2xp67_ASAP7_75t_L g2533 ( 
.A(n_1418),
.B(n_750),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2535)
);

O2A1O1Ixp5_ASAP7_75t_L g2536 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_L g2537 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_1210),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_1220),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2543)
);

BUFx8_ASAP7_75t_L g2544 ( 
.A(n_1229),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1221),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2548)
);

NOR2xp67_ASAP7_75t_SL g2549 ( 
.A(n_1220),
.B(n_378),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_1210),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_1210),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_SL g2562 ( 
.A(n_1569),
.B(n_466),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_1210),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2569)
);

NOR2xp67_ASAP7_75t_L g2570 ( 
.A(n_1418),
.B(n_750),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2571)
);

INVx2_ASAP7_75t_SL g2572 ( 
.A(n_1220),
.Y(n_2572)
);

OR2x6_ASAP7_75t_L g2573 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_1221),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1221),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_1210),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_1221),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_SL g2591 ( 
.A(n_1569),
.B(n_466),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_1221),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_1210),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_1569),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_1210),
.Y(n_2605)
);

INVx8_ASAP7_75t_L g2606 ( 
.A(n_1279),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_1210),
.Y(n_2608)
);

OR2x2_ASAP7_75t_L g2609 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2610)
);

AND3x1_ASAP7_75t_L g2611 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1221),
.Y(n_2612)
);

O2A1O1Ixp5_ASAP7_75t_L g2613 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1221),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_1569),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_R g2617 ( 
.A(n_1664),
.B(n_466),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_1210),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1221),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_1210),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2622)
);

INVx3_ASAP7_75t_L g2623 ( 
.A(n_1279),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_SL g2624 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_265),
.B2(n_288),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_1239),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_1210),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2630)
);

INVxp67_ASAP7_75t_SL g2631 ( 
.A(n_1240),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2635)
);

NOR3xp33_ASAP7_75t_L g2636 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2636)
);

NOR2xp67_ASAP7_75t_L g2637 ( 
.A(n_1418),
.B(n_750),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_1221),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2641)
);

INVx8_ASAP7_75t_L g2642 ( 
.A(n_1279),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2644)
);

BUFx6f_ASAP7_75t_L g2645 ( 
.A(n_1281),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2646)
);

INVx2_ASAP7_75t_SL g2647 ( 
.A(n_1220),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_1297),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_1210),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_1221),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_1221),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_1221),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_1210),
.Y(n_2659)
);

NAND3xp33_ASAP7_75t_L g2660 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2660)
);

BUFx3_ASAP7_75t_L g2661 ( 
.A(n_1220),
.Y(n_2661)
);

AND2x4_ASAP7_75t_SL g2662 ( 
.A(n_1297),
.B(n_750),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_SL g2664 ( 
.A(n_1276),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_1281),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_1221),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_1210),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_1221),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_1210),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2677)
);

HB1xp67_ASAP7_75t_L g2678 ( 
.A(n_1271),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2679)
);

BUFx3_ASAP7_75t_L g2680 ( 
.A(n_1220),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2683)
);

INVx3_ASAP7_75t_L g2684 ( 
.A(n_1279),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2686)
);

AND2x6_ASAP7_75t_L g2687 ( 
.A(n_1263),
.B(n_1264),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2688)
);

AND2x4_ASAP7_75t_L g2689 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2691)
);

AND2x6_ASAP7_75t_SL g2692 ( 
.A(n_1213),
.B(n_1218),
.Y(n_2692)
);

O2A1O1Ixp33_ASAP7_75t_L g2693 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1535),
.C(n_1226),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1221),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2697)
);

OR2x2_ASAP7_75t_L g2698 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_1221),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_1221),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2704)
);

INVxp67_ASAP7_75t_L g2705 ( 
.A(n_1239),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_1281),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2709)
);

OR2x6_ASAP7_75t_L g2710 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_1221),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_1220),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_SL g2716 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1845),
.B2(n_1587),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_1210),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_1221),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_1210),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2725)
);

AND3x2_ASAP7_75t_L g2726 ( 
.A(n_1249),
.B(n_844),
.C(n_1311),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_1221),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_1279),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2730)
);

INVxp67_ASAP7_75t_L g2731 ( 
.A(n_1239),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2733)
);

INVx4_ASAP7_75t_L g2734 ( 
.A(n_1308),
.Y(n_2734)
);

OR2x6_ASAP7_75t_L g2735 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_1210),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_1221),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_1210),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_1210),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2743)
);

O2A1O1Ixp5_ASAP7_75t_L g2744 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2744)
);

INVxp67_ASAP7_75t_SL g2745 ( 
.A(n_1240),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_1210),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2747)
);

A2O1A1Ixp33_ASAP7_75t_L g2748 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1249),
.C(n_1628),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_1221),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2754)
);

AND2x6_ASAP7_75t_SL g2755 ( 
.A(n_1213),
.B(n_1218),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_1279),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_1210),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_1210),
.Y(n_2766)
);

AOI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_1221),
.Y(n_2768)
);

BUFx2_ASAP7_75t_L g2769 ( 
.A(n_1361),
.Y(n_2769)
);

INVx5_ASAP7_75t_L g2770 ( 
.A(n_1279),
.Y(n_2770)
);

NOR2xp67_ASAP7_75t_L g2771 ( 
.A(n_1418),
.B(n_750),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_1271),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_SL g2774 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_1221),
.Y(n_2780)
);

AND2x4_ASAP7_75t_L g2781 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_1221),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_1221),
.Y(n_2787)
);

INVxp67_ASAP7_75t_SL g2788 ( 
.A(n_1240),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2789)
);

NOR2xp33_ASAP7_75t_L g2790 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2790)
);

NOR3xp33_ASAP7_75t_L g2791 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2795)
);

AOI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_1281),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2798)
);

AOI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1221),
.Y(n_2800)
);

INVx1_ASAP7_75t_SL g2801 ( 
.A(n_1635),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_1221),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_1210),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_1210),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_1271),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_1221),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_1220),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_SL g2810 ( 
.A(n_1747),
.B(n_1845),
.C(n_1587),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_1210),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_1210),
.Y(n_2815)
);

AND2x6_ASAP7_75t_L g2816 ( 
.A(n_1263),
.B(n_1264),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1221),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_1221),
.Y(n_2818)
);

AOI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_1210),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_1210),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_1221),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2825)
);

INVx1_ASAP7_75t_SL g2826 ( 
.A(n_1635),
.Y(n_2826)
);

OAI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_1240),
.A2(n_1587),
.B1(n_1892),
.B2(n_1845),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2829)
);

AOI22xp33_ASAP7_75t_L g2830 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_1221),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_1221),
.Y(n_2835)
);

OAI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_1240),
.A2(n_1587),
.B1(n_1892),
.B2(n_1845),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_2838)
);

O2A1O1Ixp5_ASAP7_75t_L g2839 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_1569),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_1221),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2845)
);

NAND2xp33_ASAP7_75t_L g2846 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2849)
);

CKINVDCx20_ASAP7_75t_R g2850 ( 
.A(n_1297),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_1220),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2852)
);

O2A1O1Ixp5_ASAP7_75t_L g2853 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2854)
);

NOR3xp33_ASAP7_75t_L g2855 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_1221),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2858)
);

A2O1A1Ixp33_ASAP7_75t_SL g2859 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1603),
.C(n_1517),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_1220),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_1210),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_SL g2865 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_1210),
.Y(n_2868)
);

AOI22xp33_ASAP7_75t_L g2869 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_1221),
.Y(n_2870)
);

O2A1O1Ixp5_ASAP7_75t_L g2871 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2871)
);

AOI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_SL g2873 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2874)
);

OR2x6_ASAP7_75t_L g2875 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2875)
);

INVx4_ASAP7_75t_L g2876 ( 
.A(n_1308),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_1569),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2878)
);

O2A1O1Ixp5_ASAP7_75t_L g2879 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_L g2880 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_1221),
.Y(n_2881)
);

AND2x4_ASAP7_75t_L g2882 ( 
.A(n_1281),
.B(n_1319),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2885)
);

INVx4_ASAP7_75t_L g2886 ( 
.A(n_1308),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_1221),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_1220),
.Y(n_2890)
);

INVx8_ASAP7_75t_L g2891 ( 
.A(n_1279),
.Y(n_2891)
);

AOI22xp33_ASAP7_75t_L g2892 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2892)
);

NAND2x1_ASAP7_75t_L g2893 ( 
.A(n_1231),
.B(n_889),
.Y(n_2893)
);

BUFx3_ASAP7_75t_L g2894 ( 
.A(n_1220),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_1210),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2897)
);

AOI22xp33_ASAP7_75t_L g2898 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_1221),
.Y(n_2900)
);

AOI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_1221),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2906)
);

AND2x6_ASAP7_75t_SL g2907 ( 
.A(n_1213),
.B(n_1218),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2908)
);

AOI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2909)
);

BUFx6f_ASAP7_75t_L g2910 ( 
.A(n_1281),
.Y(n_2910)
);

HB1xp67_ASAP7_75t_L g2911 ( 
.A(n_1271),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_1221),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_1210),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2916)
);

INVxp33_ASAP7_75t_L g2917 ( 
.A(n_1740),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_1210),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_1210),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_1554),
.B(n_1240),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_1210),
.Y(n_2923)
);

A2O1A1Ixp33_ASAP7_75t_L g2924 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1249),
.C(n_1628),
.Y(n_2924)
);

OAI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_1226),
.A2(n_1231),
.B(n_1344),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2927)
);

OR2x6_ASAP7_75t_L g2928 ( 
.A(n_1279),
.B(n_1289),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_1220),
.Y(n_2929)
);

O2A1O1Ixp33_ASAP7_75t_L g2930 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1535),
.C(n_1226),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_1220),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_1210),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_1221),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2937)
);

OAI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_1210),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2942)
);

INVx2_ASAP7_75t_SL g2943 ( 
.A(n_1220),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_1210),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_1210),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_1221),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_1210),
.Y(n_2953)
);

INVxp67_ASAP7_75t_L g2954 ( 
.A(n_1239),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_1257),
.B(n_1298),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_1220),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_1569),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2965)
);

NAND2xp33_ASAP7_75t_L g2966 ( 
.A(n_1240),
.B(n_1517),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_1210),
.Y(n_2969)
);

NOR2xp33_ASAP7_75t_SL g2970 ( 
.A(n_1569),
.B(n_466),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_1226),
.B(n_1293),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2979)
);

NAND3xp33_ASAP7_75t_SL g2980 ( 
.A(n_1747),
.B(n_1845),
.C(n_1587),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2982)
);

NOR2x2_ASAP7_75t_L g2983 ( 
.A(n_1496),
.B(n_1005),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_1554),
.B(n_1344),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_1221),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_1210),
.Y(n_2989)
);

INVx4_ASAP7_75t_L g2990 ( 
.A(n_1308),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_1210),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_1226),
.B(n_1344),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_1210),
.Y(n_2993)
);

INVx2_ASAP7_75t_SL g2994 ( 
.A(n_1220),
.Y(n_2994)
);

INVx1_ASAP7_75t_SL g2995 ( 
.A(n_1635),
.Y(n_2995)
);

O2A1O1Ixp5_ASAP7_75t_L g2996 ( 
.A1(n_1495),
.A2(n_1231),
.B(n_1240),
.C(n_1554),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_1226),
.B(n_1212),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_1281),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_1210),
.Y(n_3001)
);

INVx2_ASAP7_75t_SL g3002 ( 
.A(n_1220),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_1221),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_1221),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_1210),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3007)
);

AOI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_SL g3009 ( 
.A(n_1554),
.B(n_1344),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_1221),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_1554),
.B(n_1344),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_3013)
);

BUFx6f_ASAP7_75t_L g3014 ( 
.A(n_1281),
.Y(n_3014)
);

AND2x4_ASAP7_75t_SL g3015 ( 
.A(n_1297),
.B(n_750),
.Y(n_3015)
);

INVx4_ASAP7_75t_L g3016 ( 
.A(n_1308),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_SL g3020 ( 
.A(n_1554),
.B(n_1344),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_1240),
.A2(n_1554),
.B(n_1507),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3022)
);

INVxp67_ASAP7_75t_L g3023 ( 
.A(n_1239),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3024)
);

INVxp67_ASAP7_75t_L g3025 ( 
.A(n_1239),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_1221),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_1210),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_1210),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_1221),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_1226),
.B(n_1293),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_SL g3033 ( 
.A(n_1554),
.B(n_1240),
.Y(n_3033)
);

NAND3xp33_ASAP7_75t_SL g3034 ( 
.A(n_1747),
.B(n_1845),
.C(n_1587),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3035)
);

AOI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1226),
.B2(n_1747),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3039)
);

A2O1A1Ixp33_ASAP7_75t_L g3040 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1249),
.C(n_1628),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3041)
);

INVx4_ASAP7_75t_L g3042 ( 
.A(n_1308),
.Y(n_3042)
);

NOR3xp33_ASAP7_75t_L g3043 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_1226),
.B(n_1293),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_1554),
.B(n_1344),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_1281),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_1221),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_1240),
.A2(n_1226),
.B1(n_1845),
.B2(n_1587),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_1249),
.A2(n_844),
.B1(n_1246),
.B2(n_1244),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_1281),
.B(n_1319),
.Y(n_3052)
);

AND2x4_ASAP7_75t_L g3053 ( 
.A(n_1281),
.B(n_1319),
.Y(n_3053)
);

OAI22xp5_ASAP7_75t_SL g3054 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1845),
.B2(n_1587),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_1210),
.Y(n_3055)
);

A2O1A1Ixp33_ASAP7_75t_L g3056 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1249),
.C(n_1628),
.Y(n_3056)
);

NAND2xp33_ASAP7_75t_L g3057 ( 
.A(n_1240),
.B(n_1517),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3058)
);

INVx2_ASAP7_75t_SL g3059 ( 
.A(n_1220),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3061)
);

HB1xp67_ASAP7_75t_L g3062 ( 
.A(n_1271),
.Y(n_3062)
);

NOR3xp33_ASAP7_75t_L g3063 ( 
.A(n_1747),
.B(n_1218),
.C(n_1213),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_1210),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_1226),
.B(n_1344),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_1210),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_1226),
.B(n_1212),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_1221),
.Y(n_3070)
);

OR2x6_ASAP7_75t_L g3071 ( 
.A(n_1279),
.B(n_1289),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3074)
);

AO21x1_ASAP7_75t_L g3075 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3075)
);

OAI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_2005),
.B2(n_2084),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_SL g3078 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2631),
.Y(n_3079)
);

CKINVDCx20_ASAP7_75t_R g3080 ( 
.A(n_2257),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2745),
.B(n_2788),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2138),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2788),
.B(n_1936),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2584),
.A2(n_2779),
.B(n_2644),
.Y(n_3086)
);

AND2x2_ASAP7_75t_SL g3087 ( 
.A(n_1914),
.B(n_2041),
.Y(n_3087)
);

AOI21xp5_ASAP7_75t_L g3088 ( 
.A1(n_2786),
.A2(n_2838),
.B(n_2799),
.Y(n_3088)
);

AO22x1_ASAP7_75t_L g3089 ( 
.A1(n_2065),
.A2(n_2084),
.B1(n_2061),
.B2(n_2062),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_1936),
.B(n_1937),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2138),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_1937),
.B(n_2064),
.Y(n_3092)
);

NOR2x1_ASAP7_75t_L g3093 ( 
.A(n_2323),
.B(n_2334),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_SL g3094 ( 
.A(n_2836),
.B(n_2938),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_3021),
.A2(n_2518),
.B(n_2509),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2138),
.Y(n_3096)
);

AO22x1_ASAP7_75t_L g3097 ( 
.A1(n_2065),
.A2(n_2061),
.B1(n_2062),
.B2(n_2057),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2836),
.B(n_2952),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_SL g3099 ( 
.A(n_2040),
.B(n_2017),
.Y(n_3099)
);

NAND2x1p5_ASAP7_75t_L g3100 ( 
.A(n_2041),
.B(n_2893),
.Y(n_3100)
);

OAI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_3050),
.A2(n_2748),
.B(n_2455),
.Y(n_3101)
);

AND2x4_ASAP7_75t_L g3102 ( 
.A(n_2103),
.B(n_2252),
.Y(n_3102)
);

OAI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2924),
.A2(n_3056),
.B(n_3040),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2064),
.B(n_2518),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_1923),
.B(n_2311),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2525),
.A2(n_2675),
.B(n_2668),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2525),
.B(n_2668),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2675),
.B(n_2676),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_1918),
.A2(n_2369),
.B(n_2367),
.Y(n_3109)
);

AOI21x1_ASAP7_75t_L g3110 ( 
.A1(n_2676),
.A2(n_2683),
.B(n_2679),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_1914),
.B(n_2453),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2138),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2138),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2138),
.Y(n_3114)
);

AO21x1_ASAP7_75t_L g3115 ( 
.A1(n_2679),
.A2(n_2695),
.B(n_2683),
.Y(n_3115)
);

OAI321xp33_ASAP7_75t_L g3116 ( 
.A1(n_2373),
.A2(n_2414),
.A3(n_2406),
.B1(n_2425),
.B2(n_2412),
.C(n_2390),
.Y(n_3116)
);

BUFx6f_ASAP7_75t_L g3117 ( 
.A(n_2319),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_SL g3118 ( 
.A(n_2716),
.B(n_3054),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3119)
);

AOI21x1_ASAP7_75t_L g3120 ( 
.A1(n_2695),
.A2(n_2822),
.B(n_2774),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2774),
.A2(n_2899),
.B(n_2822),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2317),
.A2(n_2372),
.B1(n_2387),
.B2(n_2325),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2068),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2316),
.B(n_2329),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2899),
.B(n_2921),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2435),
.A2(n_2468),
.B1(n_2469),
.B2(n_2457),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2921),
.A2(n_3033),
.B(n_2922),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2558),
.A2(n_2576),
.B1(n_2587),
.B2(n_2571),
.Y(n_3128)
);

OAI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2434),
.A2(n_2494),
.B(n_2460),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2286),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_1944),
.B(n_2293),
.Y(n_3131)
);

AOI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_2922),
.A2(n_3033),
.B(n_2007),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_SL g3133 ( 
.A(n_1947),
.B(n_2052),
.Y(n_3133)
);

OAI321xp33_ASAP7_75t_L g3134 ( 
.A1(n_2495),
.A2(n_2496),
.A3(n_2561),
.B1(n_2648),
.B2(n_2635),
.C(n_2596),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2024),
.B(n_2054),
.Y(n_3135)
);

AOI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_2316),
.A2(n_2329),
.B1(n_2386),
.B2(n_2357),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2319),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2019),
.A2(n_1934),
.B(n_2536),
.Y(n_3138)
);

OAI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2649),
.A2(n_2667),
.B(n_2654),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2286),
.Y(n_3140)
);

O2A1O1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_2304),
.A2(n_2337),
.B(n_2980),
.C(n_2810),
.Y(n_3141)
);

AO21x1_ASAP7_75t_L g3142 ( 
.A1(n_2697),
.A2(n_2775),
.B(n_2712),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_1968),
.B(n_1969),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2536),
.A2(n_2744),
.B(n_2613),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2633),
.B(n_2704),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_2005),
.B2(n_2056),
.Y(n_3146)
);

AOI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_2613),
.A2(n_2839),
.B(n_2744),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_1968),
.B(n_1969),
.Y(n_3148)
);

AOI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2839),
.A2(n_2871),
.B(n_2853),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2853),
.A2(n_2879),
.B(n_2871),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_1952),
.B(n_2069),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2135),
.B(n_2202),
.Y(n_3152)
);

OR2x2_ASAP7_75t_L g3153 ( 
.A(n_2336),
.B(n_2338),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_2103),
.B(n_2252),
.Y(n_3154)
);

OAI21xp33_ASAP7_75t_L g3155 ( 
.A1(n_2720),
.A2(n_2819),
.B(n_2793),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2879),
.A2(n_2996),
.B(n_2034),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_1940),
.B(n_2028),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2996),
.A2(n_2035),
.B(n_1940),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2828),
.A2(n_2845),
.B(n_2843),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2733),
.B(n_2796),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_SL g3161 ( 
.A(n_2074),
.B(n_2878),
.Y(n_3161)
);

OAI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2847),
.A2(n_2858),
.B(n_2854),
.Y(n_3162)
);

OAI21xp33_ASAP7_75t_L g3163 ( 
.A1(n_2935),
.A2(n_2936),
.B(n_2909),
.Y(n_3163)
);

NOR2xp33_ASAP7_75t_L g3164 ( 
.A(n_2901),
.B(n_2974),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2863),
.A2(n_2873),
.B(n_2865),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_1952),
.B(n_1919),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_2068),
.Y(n_3167)
);

OAI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2874),
.A2(n_2948),
.B(n_2937),
.Y(n_3168)
);

CKINVDCx6p67_ASAP7_75t_R g3169 ( 
.A(n_2305),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2135),
.Y(n_3170)
);

AOI21x1_ASAP7_75t_L g3171 ( 
.A1(n_2043),
.A2(n_2105),
.B(n_2955),
.Y(n_3171)
);

AOI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_2961),
.A2(n_2978),
.B(n_2973),
.Y(n_3172)
);

A2O1A1Ixp33_ASAP7_75t_L g3173 ( 
.A1(n_2055),
.A2(n_1933),
.B(n_2693),
.C(n_2362),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_3036),
.B(n_3013),
.Y(n_3174)
);

O2A1O1Ixp33_ASAP7_75t_L g3175 ( 
.A1(n_3034),
.A2(n_2501),
.B(n_2636),
.C(n_2420),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2982),
.A2(n_3009),
.B(n_2984),
.Y(n_3176)
);

NOR2xp33_ASAP7_75t_L g3177 ( 
.A(n_2332),
.B(n_2660),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3012),
.B(n_3020),
.Y(n_3178)
);

OR2x6_ASAP7_75t_L g3179 ( 
.A(n_2224),
.B(n_2419),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3045),
.B(n_2289),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_2326),
.A2(n_2416),
.B(n_2400),
.Y(n_3181)
);

AOI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_2537),
.A2(n_2966),
.B(n_2846),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_3057),
.A2(n_2013),
.B(n_2043),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_1933),
.A2(n_2930),
.B(n_2037),
.Y(n_3184)
);

AOI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2357),
.A2(n_2407),
.B1(n_2437),
.B2(n_2386),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2289),
.B(n_2313),
.Y(n_3186)
);

OAI21xp33_ASAP7_75t_L g3187 ( 
.A1(n_2420),
.A2(n_2636),
.B(n_2501),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2202),
.Y(n_3188)
);

O2A1O1Ixp5_ASAP7_75t_L g3189 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2700),
.C(n_2018),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2454),
.A2(n_2925),
.B(n_2430),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2328),
.A2(n_2859),
.B(n_2430),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2328),
.A2(n_2859),
.B(n_2140),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_2407),
.A2(n_2443),
.B1(n_2473),
.B2(n_2437),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_2443),
.B(n_2473),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2032),
.A2(n_2036),
.B(n_1955),
.Y(n_3195)
);

INVxp67_ASAP7_75t_L g3196 ( 
.A(n_2004),
.Y(n_3196)
);

OAI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_2791),
.A2(n_3043),
.B(n_2855),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_1930),
.A2(n_1931),
.B(n_2015),
.Y(n_3198)
);

HB1xp67_ASAP7_75t_L g3199 ( 
.A(n_2356),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_2791),
.A2(n_3043),
.B(n_2855),
.Y(n_3200)
);

OR2x2_ASAP7_75t_L g3201 ( 
.A(n_2397),
.B(n_2594),
.Y(n_3201)
);

O2A1O1Ixp33_ASAP7_75t_SL g3202 ( 
.A1(n_1931),
.A2(n_2047),
.B(n_2053),
.C(n_2044),
.Y(n_3202)
);

NAND3xp33_ASAP7_75t_L g3203 ( 
.A(n_3063),
.B(n_2611),
.C(n_2488),
.Y(n_3203)
);

OR2x2_ASAP7_75t_L g3204 ( 
.A(n_2609),
.B(n_2628),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2313),
.B(n_2340),
.Y(n_3205)
);

BUFx3_ASAP7_75t_L g3206 ( 
.A(n_2068),
.Y(n_3206)
);

O2A1O1Ixp33_ASAP7_75t_L g3207 ( 
.A1(n_3063),
.A2(n_2063),
.B(n_2075),
.C(n_2071),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2340),
.B(n_2341),
.Y(n_3208)
);

O2A1O1Ixp33_ASAP7_75t_SL g3209 ( 
.A1(n_2077),
.A2(n_1941),
.B(n_2488),
.C(n_2476),
.Y(n_3209)
);

O2A1O1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2476),
.A2(n_2499),
.B(n_2505),
.C(n_2503),
.Y(n_3210)
);

OAI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2499),
.A2(n_2505),
.B(n_2503),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2341),
.B(n_2342),
.Y(n_3212)
);

NAND2x1p5_ASAP7_75t_L g3213 ( 
.A(n_2099),
.B(n_2120),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2342),
.B(n_2359),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_1922),
.B(n_2302),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_SL g3216 ( 
.A(n_2726),
.B(n_2057),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2728),
.A2(n_2772),
.B(n_2764),
.Y(n_3217)
);

A2O1A1Ixp33_ASAP7_75t_L g3218 ( 
.A1(n_2516),
.A2(n_2528),
.B(n_2560),
.C(n_2552),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2728),
.A2(n_2772),
.B(n_2764),
.Y(n_3219)
);

INVx4_ASAP7_75t_L g3220 ( 
.A(n_2319),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2234),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2359),
.B(n_2379),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_2308),
.B(n_2348),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2379),
.B(n_2441),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_2528),
.A2(n_2677),
.B(n_2656),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2656),
.A2(n_2913),
.B(n_2708),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2235),
.Y(n_3227)
);

A2O1A1Ixp33_ASAP7_75t_L g3228 ( 
.A1(n_2516),
.A2(n_2552),
.B(n_2564),
.C(n_2560),
.Y(n_3228)
);

O2A1O1Ixp33_ASAP7_75t_L g3229 ( 
.A1(n_2564),
.A2(n_2581),
.B(n_2626),
.C(n_2595),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2441),
.B(n_2449),
.Y(n_3230)
);

OAI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_2581),
.A2(n_2626),
.B(n_2595),
.Y(n_3231)
);

BUFx4f_ASAP7_75t_SL g3232 ( 
.A(n_2153),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_1929),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2867),
.A2(n_2941),
.B(n_2888),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_1939),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_2663),
.B(n_2677),
.Y(n_3236)
);

AND2x4_ASAP7_75t_L g3237 ( 
.A(n_2770),
.B(n_2319),
.Y(n_3237)
);

HB1xp67_ASAP7_75t_L g3238 ( 
.A(n_2356),
.Y(n_3238)
);

OAI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_2663),
.A2(n_2686),
.B(n_2681),
.Y(n_3239)
);

CKINVDCx20_ASAP7_75t_R g3240 ( 
.A(n_2349),
.Y(n_3240)
);

AOI21x1_ASAP7_75t_L g3241 ( 
.A1(n_2110),
.A2(n_2187),
.B(n_2149),
.Y(n_3241)
);

AO21x1_ASAP7_75t_L g3242 ( 
.A1(n_2066),
.A2(n_2081),
.B(n_2087),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2681),
.B(n_2686),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2696),
.A2(n_2743),
.B(n_2708),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2743),
.A2(n_3017),
.B(n_2913),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_2364),
.Y(n_3246)
);

AOI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_2926),
.A2(n_2761),
.B(n_2696),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2761),
.A2(n_2906),
.B(n_2867),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2888),
.A2(n_3067),
.B(n_3024),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_1942),
.Y(n_3250)
);

NOR2xp67_ASAP7_75t_L g3251 ( 
.A(n_2110),
.B(n_2288),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_2821),
.A2(n_2926),
.B(n_2848),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_SL g3253 ( 
.A(n_2789),
.B(n_2790),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2449),
.B(n_2479),
.Y(n_3254)
);

CKINVDCx8_ASAP7_75t_R g3255 ( 
.A(n_2107),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_2834),
.A2(n_2906),
.B(n_2790),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3024),
.A2(n_2821),
.B(n_2789),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2831),
.B(n_2834),
.Y(n_3258)
);

BUFx2_ASAP7_75t_L g3259 ( 
.A(n_2364),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2479),
.B(n_2527),
.Y(n_3260)
);

AOI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_2831),
.A2(n_2848),
.B1(n_2941),
.B2(n_2862),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2527),
.B(n_2547),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_2987),
.A2(n_3061),
.B(n_2965),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2987),
.A2(n_3061),
.B(n_2965),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2862),
.B(n_2976),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2320),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3007),
.A2(n_2992),
.B(n_2976),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_2992),
.A2(n_3017),
.B1(n_3018),
.B2(n_3007),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3018),
.A2(n_3048),
.B(n_3065),
.Y(n_3269)
);

AND2x2_ASAP7_75t_SL g3270 ( 
.A(n_2251),
.B(n_2006),
.Y(n_3270)
);

INVx3_ASAP7_75t_L g3271 ( 
.A(n_2068),
.Y(n_3271)
);

AO21x1_ASAP7_75t_L g3272 ( 
.A1(n_2066),
.A2(n_2188),
.B(n_2026),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_1946),
.Y(n_3273)
);

OAI22xp5_ASAP7_75t_L g3274 ( 
.A1(n_3048),
.A2(n_3067),
.B1(n_3065),
.B2(n_1935),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_2417),
.B(n_2482),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2547),
.B(n_2569),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_1917),
.A2(n_1928),
.B(n_1927),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_2079),
.A2(n_2296),
.B(n_1915),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2307),
.A2(n_2310),
.B(n_2309),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_1945),
.A2(n_1954),
.B(n_1950),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2569),
.B(n_2578),
.Y(n_3281)
);

OAI22xp33_ASAP7_75t_L g3282 ( 
.A1(n_2314),
.A2(n_2318),
.B1(n_2333),
.B2(n_2321),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_1957),
.A2(n_1960),
.B(n_1959),
.Y(n_3283)
);

OAI321xp33_ASAP7_75t_L g3284 ( 
.A1(n_2006),
.A2(n_2042),
.A3(n_2031),
.B1(n_2076),
.B2(n_2039),
.C(n_2578),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_1964),
.A2(n_1970),
.B(n_1967),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2597),
.B(n_2600),
.Y(n_3286)
);

AOI21x1_ASAP7_75t_L g3287 ( 
.A1(n_2164),
.A2(n_2209),
.B(n_3070),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2597),
.B(n_2600),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_1971),
.A2(n_1983),
.B(n_1973),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2602),
.B(n_2630),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2602),
.B(n_2630),
.Y(n_3291)
);

NAND2x1p5_ASAP7_75t_L g3292 ( 
.A(n_2320),
.B(n_2360),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_1935),
.B(n_1958),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2699),
.B(n_2751),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_1972),
.Y(n_3295)
);

O2A1O1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_2009),
.A2(n_1958),
.B(n_2346),
.C(n_2339),
.Y(n_3296)
);

NOR2xp33_ASAP7_75t_L g3297 ( 
.A(n_2692),
.B(n_2755),
.Y(n_3297)
);

A2O1A1Ixp33_ASAP7_75t_L g3298 ( 
.A1(n_2699),
.A2(n_2767),
.B(n_2785),
.C(n_2751),
.Y(n_3298)
);

OAI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_2350),
.A2(n_2354),
.B(n_2351),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_2907),
.B(n_2358),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_1985),
.A2(n_1991),
.B(n_1986),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_1992),
.A2(n_2010),
.B(n_1996),
.Y(n_3302)
);

NOR2x2_ASAP7_75t_L g3303 ( 
.A(n_2419),
.B(n_2521),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_2068),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_2012),
.A2(n_1982),
.B(n_1978),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2767),
.B(n_2785),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_L g3307 ( 
.A(n_2370),
.B(n_2375),
.Y(n_3307)
);

AO21x1_ASAP7_75t_L g3308 ( 
.A1(n_2106),
.A2(n_2275),
.B(n_2111),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2830),
.B(n_2841),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2830),
.B(n_2841),
.Y(n_3310)
);

O2A1O1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_2009),
.A2(n_2376),
.B(n_2380),
.C(n_2378),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_1916),
.Y(n_3312)
);

O2A1O1Ixp33_ASAP7_75t_L g3313 ( 
.A1(n_2381),
.A2(n_2382),
.B(n_2391),
.C(n_2389),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_1977),
.Y(n_3314)
);

NOR2x1p5_ASAP7_75t_L g3315 ( 
.A(n_2089),
.B(n_2320),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_2365),
.B(n_2371),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_1988),
.A2(n_1993),
.B(n_1989),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2398),
.B(n_2402),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2842),
.B(n_2869),
.Y(n_3319)
);

AOI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_2842),
.A2(n_2872),
.B1(n_2880),
.B2(n_2869),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2872),
.B(n_2880),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2887),
.B(n_2892),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_2368),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_1997),
.A2(n_2008),
.B(n_2001),
.Y(n_3324)
);

BUFx3_ASAP7_75t_L g3325 ( 
.A(n_2687),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_1984),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_2887),
.B(n_2892),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2404),
.B(n_2422),
.Y(n_3328)
);

INVx3_ASAP7_75t_L g3329 ( 
.A(n_2687),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_2423),
.B(n_2428),
.Y(n_3330)
);

HB1xp67_ASAP7_75t_L g3331 ( 
.A(n_2368),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2431),
.B(n_2433),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2436),
.B(n_2438),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_1990),
.Y(n_3334)
);

OAI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2440),
.A2(n_2445),
.B(n_2444),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2447),
.B(n_2451),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_1995),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2456),
.B(n_2458),
.Y(n_3338)
);

OR2x6_ASAP7_75t_L g3339 ( 
.A(n_2419),
.B(n_2521),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2461),
.B(n_2462),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_2403),
.B(n_2467),
.Y(n_3341)
);

AOI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2109),
.A2(n_2118),
.B(n_2116),
.Y(n_3342)
);

INVxp67_ASAP7_75t_L g3343 ( 
.A(n_1962),
.Y(n_3343)
);

A2O1A1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_2898),
.A2(n_2946),
.B(n_2958),
.C(n_2903),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_2122),
.A2(n_2124),
.B(n_2123),
.Y(n_3345)
);

O2A1O1Ixp5_ASAP7_75t_L g3346 ( 
.A1(n_2072),
.A2(n_2139),
.B(n_2137),
.C(n_2130),
.Y(n_3346)
);

NOR2xp33_ASAP7_75t_SL g3347 ( 
.A(n_2726),
.B(n_2770),
.Y(n_3347)
);

AOI21x1_ASAP7_75t_L g3348 ( 
.A1(n_1999),
.A2(n_2025),
.B(n_2014),
.Y(n_3348)
);

AND2x4_ASAP7_75t_L g3349 ( 
.A(n_2770),
.B(n_2320),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_2126),
.A2(n_2131),
.B(n_2129),
.Y(n_3350)
);

O2A1O1Ixp33_ASAP7_75t_L g3351 ( 
.A1(n_2474),
.A2(n_2477),
.B(n_2486),
.C(n_2484),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2493),
.A2(n_2502),
.B(n_2497),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2190),
.B(n_2515),
.Y(n_3353)
);

INVx4_ASAP7_75t_L g3354 ( 
.A(n_2360),
.Y(n_3354)
);

BUFx6f_ASAP7_75t_L g3355 ( 
.A(n_2360),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_2517),
.A2(n_2524),
.B(n_2520),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2048),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_2898),
.B(n_2903),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2946),
.B(n_2958),
.Y(n_3359)
);

BUFx4f_ASAP7_75t_L g3360 ( 
.A(n_2360),
.Y(n_3360)
);

INVx2_ASAP7_75t_SL g3361 ( 
.A(n_2448),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_2526),
.B(n_2532),
.Y(n_3362)
);

CKINVDCx10_ASAP7_75t_R g3363 ( 
.A(n_2664),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_2534),
.B(n_2535),
.Y(n_3364)
);

AOI21x1_ASAP7_75t_L g3365 ( 
.A1(n_2049),
.A2(n_2088),
.B(n_2070),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_2541),
.A2(n_2543),
.B(n_2542),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_2967),
.B(n_2975),
.Y(n_3367)
);

BUFx3_ASAP7_75t_L g3368 ( 
.A(n_2687),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_2546),
.B(n_2548),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_2550),
.B(n_2551),
.Y(n_3370)
);

NOR2x1p5_ASAP7_75t_L g3371 ( 
.A(n_2475),
.B(n_2645),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_2557),
.B(n_2559),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_2967),
.B(n_2975),
.Y(n_3373)
);

O2A1O1Ixp33_ASAP7_75t_L g3374 ( 
.A1(n_2553),
.A2(n_2555),
.B(n_2566),
.C(n_2565),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_2567),
.B(n_2568),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2986),
.B(n_3008),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2986),
.B(n_3008),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3046),
.B(n_3051),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3046),
.B(n_3051),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2574),
.B(n_2577),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_2580),
.A2(n_2586),
.B(n_2585),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2588),
.A2(n_2598),
.B(n_2592),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_2599),
.B(n_2607),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2610),
.B(n_2615),
.Y(n_3384)
);

NAND2x1p5_ASAP7_75t_L g3385 ( 
.A(n_2475),
.B(n_2645),
.Y(n_3385)
);

INVx3_ASAP7_75t_L g3386 ( 
.A(n_2687),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2622),
.B(n_2632),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_2634),
.A2(n_2640),
.B(n_2638),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_2448),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2641),
.A2(n_2646),
.B(n_2643),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_2042),
.A2(n_2039),
.B1(n_2076),
.B2(n_2031),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_1980),
.A2(n_2666),
.B1(n_2706),
.B2(n_2690),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_2652),
.B(n_2669),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_2682),
.A2(n_2688),
.B(n_2685),
.Y(n_3394)
);

AO22x1_ASAP7_75t_L g3395 ( 
.A1(n_2687),
.A2(n_2816),
.B1(n_2137),
.B2(n_2130),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_2691),
.B(n_2702),
.Y(n_3396)
);

OAI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2709),
.A2(n_2714),
.B(n_2713),
.Y(n_3397)
);

CKINVDCx20_ASAP7_75t_R g3398 ( 
.A(n_2650),
.Y(n_3398)
);

NAND2xp33_ASAP7_75t_L g3399 ( 
.A(n_2719),
.B(n_2721),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_2722),
.A2(n_2730),
.B(n_2725),
.Y(n_3400)
);

O2A1O1Ixp33_ASAP7_75t_SL g3401 ( 
.A1(n_2096),
.A2(n_2737),
.B(n_2752),
.C(n_2732),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_2753),
.B(n_2754),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2092),
.Y(n_3403)
);

O2A1O1Ixp33_ASAP7_75t_SL g3404 ( 
.A1(n_2096),
.A2(n_2759),
.B(n_2760),
.C(n_2757),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2094),
.Y(n_3405)
);

A2O1A1Ixp33_ASAP7_75t_L g3406 ( 
.A1(n_2762),
.A2(n_2763),
.B(n_2776),
.C(n_2765),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2777),
.B(n_2778),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_2782),
.B(n_2783),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2792),
.B(n_2794),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2795),
.A2(n_2808),
.B(n_2798),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_2575),
.B(n_2582),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2809),
.B(n_2811),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2812),
.A2(n_2829),
.B(n_2825),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_2832),
.A2(n_2849),
.B(n_2837),
.Y(n_3414)
);

OAI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_2852),
.A2(n_2864),
.B(n_2857),
.Y(n_3415)
);

O2A1O1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_2866),
.A2(n_2883),
.B(n_2885),
.C(n_2884),
.Y(n_3416)
);

A2O1A1Ixp33_ASAP7_75t_L g3417 ( 
.A1(n_2896),
.A2(n_2897),
.B(n_2905),
.C(n_2904),
.Y(n_3417)
);

AO21x1_ASAP7_75t_L g3418 ( 
.A1(n_2106),
.A2(n_2275),
.B(n_2022),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2908),
.B(n_2915),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2916),
.B(n_2927),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2100),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_2934),
.A2(n_2942),
.B(n_2939),
.Y(n_3422)
);

OAI321xp33_ASAP7_75t_L g3423 ( 
.A1(n_1965),
.A2(n_1980),
.A3(n_2951),
.B1(n_2956),
.B2(n_2950),
.C(n_2944),
.Y(n_3423)
);

INVx4_ASAP7_75t_L g3424 ( 
.A(n_2475),
.Y(n_3424)
);

A2O1A1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_2957),
.A2(n_2962),
.B(n_2968),
.C(n_2959),
.Y(n_3425)
);

BUFx4f_ASAP7_75t_L g3426 ( 
.A(n_2475),
.Y(n_3426)
);

OAI21xp33_ASAP7_75t_L g3427 ( 
.A1(n_3058),
.A2(n_3064),
.B(n_3060),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_2972),
.A2(n_2979),
.B(n_2977),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_2645),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2112),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_SL g3431 ( 
.A(n_2213),
.B(n_2098),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_2981),
.B(n_2985),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_2997),
.A2(n_2999),
.B(n_2998),
.Y(n_3433)
);

O2A1O1Ixp33_ASAP7_75t_L g3434 ( 
.A1(n_3005),
.A2(n_3011),
.B(n_3022),
.C(n_3019),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_3027),
.B(n_3030),
.Y(n_3435)
);

OAI21xp33_ASAP7_75t_L g3436 ( 
.A1(n_3069),
.A2(n_3037),
.B(n_3035),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3038),
.B(n_3039),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3041),
.A2(n_1975),
.B(n_2237),
.Y(n_3438)
);

OAI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_1965),
.A2(n_2086),
.B(n_2604),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_2238),
.A2(n_2276),
.B(n_2249),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2114),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_2150),
.A2(n_2161),
.B(n_2156),
.Y(n_3442)
);

HB1xp67_ASAP7_75t_L g3443 ( 
.A(n_2678),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2165),
.A2(n_2176),
.B(n_2170),
.Y(n_3444)
);

AO21x1_ASAP7_75t_L g3445 ( 
.A1(n_2022),
.A2(n_2180),
.B(n_2179),
.Y(n_3445)
);

A2O1A1Ixp33_ASAP7_75t_L g3446 ( 
.A1(n_2090),
.A2(n_2095),
.B(n_2113),
.C(n_2233),
.Y(n_3446)
);

INVxp67_ASAP7_75t_L g3447 ( 
.A(n_1963),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2185),
.A2(n_2197),
.B(n_2193),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_2201),
.A2(n_2208),
.B(n_2207),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_2217),
.A2(n_2218),
.B(n_2141),
.Y(n_3450)
);

HB1xp67_ASAP7_75t_L g3451 ( 
.A(n_2678),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2115),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2168),
.B(n_2134),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_2618),
.B(n_2655),
.Y(n_3454)
);

AOI21xp33_ASAP7_75t_L g3455 ( 
.A1(n_2168),
.A2(n_2917),
.B(n_1924),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_2223),
.A2(n_2227),
.B(n_2214),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_2223),
.A2(n_2214),
.B(n_2205),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_R g3458 ( 
.A(n_2850),
.B(n_2283),
.Y(n_3458)
);

INVx1_ASAP7_75t_SL g3459 ( 
.A(n_2093),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_2205),
.A2(n_2147),
.B(n_1951),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_1948),
.A2(n_1953),
.B(n_2671),
.Y(n_3461)
);

O2A1O1Ixp5_ASAP7_75t_L g3462 ( 
.A1(n_2167),
.A2(n_2219),
.B(n_2256),
.C(n_2233),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_2718),
.A2(n_2739),
.B1(n_2813),
.B2(n_2741),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2145),
.B(n_2146),
.Y(n_3464)
);

INVx3_ASAP7_75t_L g3465 ( 
.A(n_2816),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2918),
.A2(n_3032),
.B(n_2971),
.Y(n_3466)
);

BUFx12f_ASAP7_75t_L g3467 ( 
.A(n_2153),
.Y(n_3467)
);

CKINVDCx10_ASAP7_75t_R g3468 ( 
.A(n_2664),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_2155),
.B(n_2173),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3044),
.A2(n_2263),
.B(n_2203),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_1943),
.B(n_2177),
.Y(n_3471)
);

OAI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_2095),
.A2(n_1938),
.B(n_2256),
.Y(n_3472)
);

AOI22xp5_ASAP7_75t_L g3473 ( 
.A1(n_1974),
.A2(n_1981),
.B1(n_2030),
.B2(n_1994),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2194),
.A2(n_2101),
.B(n_2182),
.Y(n_3474)
);

A2O1A1Ixp33_ASAP7_75t_L g3475 ( 
.A1(n_2113),
.A2(n_2222),
.B(n_1956),
.C(n_2183),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2200),
.B(n_2290),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2298),
.B(n_2303),
.Y(n_3477)
);

INVx3_ASAP7_75t_L g3478 ( 
.A(n_2816),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2347),
.B(n_2353),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_2816),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_1938),
.B(n_2085),
.Y(n_3481)
);

CKINVDCx5p33_ASAP7_75t_R g3482 ( 
.A(n_2617),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_2361),
.A2(n_2388),
.B(n_2385),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_2216),
.B(n_2148),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_2216),
.B(n_2645),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_2665),
.B(n_2707),
.Y(n_3486)
);

AO21x1_ASAP7_75t_L g3487 ( 
.A1(n_2394),
.A2(n_2405),
.B(n_2395),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_2000),
.A2(n_2023),
.B1(n_2033),
.B2(n_2020),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2408),
.B(n_2410),
.Y(n_3489)
);

INVx2_ASAP7_75t_SL g3490 ( 
.A(n_2773),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_2222),
.A2(n_2091),
.B(n_2210),
.C(n_2098),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_2500),
.B(n_2698),
.Y(n_3492)
);

INVx3_ASAP7_75t_L g3493 ( 
.A(n_2816),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_2665),
.B(n_2707),
.Y(n_3494)
);

OAI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_2506),
.A2(n_2750),
.B1(n_2960),
.B2(n_2805),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_R g3496 ( 
.A(n_2519),
.B(n_2562),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2411),
.B(n_2415),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_2421),
.B(n_2427),
.Y(n_3498)
);

OAI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_2450),
.A2(n_2481),
.B(n_2480),
.Y(n_3499)
);

BUFx6f_ASAP7_75t_L g3500 ( 
.A(n_2665),
.Y(n_3500)
);

AOI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_2157),
.A2(n_2970),
.B1(n_2591),
.B2(n_2343),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2487),
.B(n_2489),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_2508),
.A2(n_2513),
.B(n_2512),
.Y(n_3503)
);

OAI21xp33_ASAP7_75t_L g3504 ( 
.A1(n_2773),
.A2(n_2911),
.B(n_2805),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_2514),
.B(n_2523),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_2050),
.B(n_2452),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_2531),
.A2(n_2579),
.B(n_2545),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_SL g3508 ( 
.A(n_2707),
.B(n_2797),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2583),
.A2(n_2593),
.B(n_2590),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_2707),
.B(n_2797),
.Y(n_3510)
);

OAI21xp33_ASAP7_75t_L g3511 ( 
.A1(n_2911),
.A2(n_3062),
.B(n_2240),
.Y(n_3511)
);

OAI22xp33_ASAP7_75t_L g3512 ( 
.A1(n_2119),
.A2(n_1998),
.B1(n_2226),
.B2(n_2221),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_L g3513 ( 
.A(n_2485),
.B(n_2769),
.Y(n_3513)
);

OAI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3062),
.A2(n_2614),
.B1(n_2620),
.B2(n_2612),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_2639),
.A2(n_2657),
.B(n_2653),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2658),
.B(n_2670),
.Y(n_3516)
);

AO21x1_ASAP7_75t_L g3517 ( 
.A1(n_2673),
.A2(n_2701),
.B(n_2694),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_2703),
.A2(n_2723),
.B(n_2711),
.Y(n_3518)
);

BUFx3_ASAP7_75t_L g3519 ( 
.A(n_1920),
.Y(n_3519)
);

OAI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_2727),
.A2(n_2749),
.B(n_2738),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2768),
.B(n_2780),
.Y(n_3521)
);

AOI21x1_ASAP7_75t_L g3522 ( 
.A1(n_2784),
.A2(n_2800),
.B(n_2787),
.Y(n_3522)
);

INVx5_ASAP7_75t_L g3523 ( 
.A(n_2797),
.Y(n_3523)
);

OR2x2_ASAP7_75t_L g3524 ( 
.A(n_1987),
.B(n_2343),
.Y(n_3524)
);

AOI22xp5_ASAP7_75t_L g3525 ( 
.A1(n_1987),
.A2(n_2625),
.B1(n_2705),
.B2(n_2345),
.Y(n_3525)
);

A2O1A1Ixp33_ASAP7_75t_L g3526 ( 
.A1(n_2195),
.A2(n_2215),
.B(n_2806),
.C(n_2802),
.Y(n_3526)
);

AOI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_2345),
.A2(n_2705),
.B1(n_2731),
.B2(n_2625),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_2817),
.A2(n_2824),
.B(n_2818),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2833),
.B(n_2835),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_2844),
.B(n_2856),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2870),
.A2(n_2889),
.B(n_2881),
.Y(n_3531)
);

INVxp67_ASAP7_75t_L g3532 ( 
.A(n_2801),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_2826),
.B(n_2995),
.Y(n_3533)
);

INVxp67_ASAP7_75t_L g3534 ( 
.A(n_2204),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_2900),
.A2(n_2912),
.B(n_2902),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_2933),
.A2(n_2988),
.B(n_2949),
.Y(n_3536)
);

NAND2x1p5_ASAP7_75t_L g3537 ( 
.A(n_2797),
.B(n_2910),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_2910),
.B(n_3000),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_2910),
.B(n_3000),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_2060),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_2082),
.A2(n_2104),
.B1(n_2125),
.B2(n_2102),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3003),
.B(n_3004),
.Y(n_3542)
);

AOI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3010),
.A2(n_3031),
.B(n_3026),
.Y(n_3543)
);

AOI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3049),
.A2(n_3000),
.B(n_2910),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3014),
.A2(n_3047),
.B(n_2255),
.Y(n_3545)
);

BUFx8_ASAP7_75t_L g3546 ( 
.A(n_2160),
.Y(n_3546)
);

INVx3_ASAP7_75t_L g3547 ( 
.A(n_3014),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_L g3548 ( 
.A(n_2163),
.B(n_2192),
.Y(n_3548)
);

NAND2xp33_ASAP7_75t_L g3549 ( 
.A(n_2045),
.B(n_2292),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3014),
.B(n_3047),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3014),
.A2(n_3047),
.B(n_2265),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3047),
.A2(n_2268),
.B(n_2247),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_2270),
.A2(n_2278),
.B(n_2273),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_2132),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_2128),
.B(n_2731),
.Y(n_3555)
);

BUFx4f_ASAP7_75t_L g3556 ( 
.A(n_2521),
.Y(n_3556)
);

AOI21x1_ASAP7_75t_L g3557 ( 
.A1(n_2021),
.A2(n_2174),
.B(n_2011),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_2231),
.B(n_2258),
.Y(n_3558)
);

OAI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_2954),
.A2(n_3025),
.B(n_3023),
.Y(n_3559)
);

INVx3_ASAP7_75t_L g3560 ( 
.A(n_1961),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_2021),
.A2(n_2191),
.B(n_1926),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_1920),
.A2(n_2322),
.B(n_1926),
.Y(n_3562)
);

BUFx2_ASAP7_75t_L g3563 ( 
.A(n_2954),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2163),
.B(n_2192),
.Y(n_3564)
);

INVx4_ASAP7_75t_L g3565 ( 
.A(n_2573),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3023),
.B(n_3025),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_2322),
.A2(n_2352),
.B(n_2324),
.Y(n_3567)
);

OAI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_2260),
.A2(n_2232),
.B(n_2504),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_2259),
.B(n_2262),
.Y(n_3569)
);

AOI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_2133),
.A2(n_2136),
.B1(n_2159),
.B2(n_2144),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_2266),
.B(n_2271),
.Y(n_3571)
);

AOI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_2324),
.A2(n_2363),
.B(n_2352),
.Y(n_3572)
);

O2A1O1Ixp33_ASAP7_75t_L g3573 ( 
.A1(n_2127),
.A2(n_2244),
.B(n_2245),
.C(n_2242),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_SL g3574 ( 
.A(n_2229),
.B(n_2617),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_2282),
.B(n_2172),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_2184),
.B(n_2186),
.Y(n_3576)
);

INVx1_ASAP7_75t_SL g3577 ( 
.A(n_1979),
.Y(n_3577)
);

O2A1O1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_2038),
.A2(n_2230),
.B(n_2143),
.C(n_2046),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_2189),
.B(n_2198),
.Y(n_3579)
);

O2A1O1Ixp33_ASAP7_75t_L g3580 ( 
.A1(n_2016),
.A2(n_2215),
.B(n_2171),
.C(n_1932),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_L g3581 ( 
.A(n_2374),
.B(n_2426),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_2363),
.A2(n_2429),
.B(n_2393),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_L g3583 ( 
.A1(n_2199),
.A2(n_2212),
.B1(n_2228),
.B2(n_2225),
.Y(n_3583)
);

AOI21x1_ASAP7_75t_L g3584 ( 
.A1(n_2151),
.A2(n_2243),
.B(n_2239),
.Y(n_3584)
);

INVx3_ASAP7_75t_L g3585 ( 
.A(n_1961),
.Y(n_3585)
);

OAI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_2003),
.A2(n_2051),
.B1(n_2330),
.B2(n_2027),
.Y(n_3586)
);

O2A1O1Ixp33_ASAP7_75t_L g3587 ( 
.A1(n_1921),
.A2(n_1925),
.B(n_2424),
.C(n_2399),
.Y(n_3587)
);

BUFx4f_ASAP7_75t_L g3588 ( 
.A(n_2573),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_2248),
.B(n_2299),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_2236),
.B(n_2281),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_SL g3591 ( 
.A(n_2236),
.B(n_2281),
.Y(n_3591)
);

AO21x1_ASAP7_75t_L g3592 ( 
.A1(n_2504),
.A2(n_2507),
.B(n_2344),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_2393),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_2429),
.A2(n_2538),
.B(n_2446),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2446),
.A2(n_2689),
.B(n_2538),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_2306),
.B(n_2366),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_2377),
.B(n_2383),
.Y(n_3597)
);

AOI21x1_ASAP7_75t_L g3598 ( 
.A1(n_2384),
.A2(n_2401),
.B(n_2396),
.Y(n_3598)
);

INVx3_ASAP7_75t_L g3599 ( 
.A(n_2003),
.Y(n_3599)
);

INVx2_ASAP7_75t_SL g3600 ( 
.A(n_2281),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_2281),
.B(n_2181),
.Y(n_3601)
);

AND2x4_ASAP7_75t_L g3602 ( 
.A(n_2573),
.B(n_2710),
.Y(n_3602)
);

A2O1A1Ixp33_ASAP7_75t_L g3603 ( 
.A1(n_2195),
.A2(n_2206),
.B(n_2355),
.C(n_2312),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_2413),
.B(n_2418),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_2442),
.B(n_2463),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_2689),
.A2(n_2781),
.B(n_2747),
.Y(n_3606)
);

OAI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2507),
.A2(n_2280),
.B(n_2246),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_2478),
.A2(n_2629),
.B1(n_3068),
.B2(n_3066),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_2181),
.B(n_2747),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_L g3610 ( 
.A(n_2459),
.B(n_2603),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2492),
.B(n_2511),
.Y(n_3611)
);

A2O1A1Ixp33_ASAP7_75t_L g3612 ( 
.A1(n_2472),
.A2(n_2637),
.B(n_2533),
.C(n_2570),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_2529),
.Y(n_3613)
);

OAI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_2246),
.A2(n_2280),
.B(n_2051),
.Y(n_3614)
);

OR2x2_ASAP7_75t_L g3615 ( 
.A(n_2539),
.B(n_2554),
.Y(n_3615)
);

INVx3_ASAP7_75t_L g3616 ( 
.A(n_2027),
.Y(n_3616)
);

AND2x4_ASAP7_75t_L g3617 ( 
.A(n_2710),
.B(n_2735),
.Y(n_3617)
);

OAI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2330),
.A2(n_2392),
.B(n_2335),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_2556),
.B(n_2563),
.Y(n_3619)
);

AO21x1_ASAP7_75t_L g3620 ( 
.A1(n_2589),
.A2(n_2605),
.B(n_2601),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_2616),
.B(n_2840),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_2608),
.B(n_2619),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_R g3623 ( 
.A(n_2877),
.B(n_2964),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_2781),
.A2(n_3052),
.B(n_2882),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_2181),
.B(n_2882),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3052),
.A2(n_3053),
.B(n_2735),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3053),
.A2(n_2735),
.B(n_2710),
.Y(n_3627)
);

BUFx2_ASAP7_75t_L g3628 ( 
.A(n_2029),
.Y(n_3628)
);

CKINVDCx5p33_ASAP7_75t_R g3629 ( 
.A(n_2253),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_2621),
.B(n_2651),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_SL g3631 ( 
.A(n_2181),
.B(n_2771),
.Y(n_3631)
);

INVx4_ASAP7_75t_L g3632 ( 
.A(n_3071),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_2335),
.A2(n_2522),
.B(n_2392),
.Y(n_3633)
);

AO21x1_ASAP7_75t_L g3634 ( 
.A1(n_2659),
.A2(n_2674),
.B(n_2672),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_2083),
.B(n_2178),
.Y(n_3635)
);

AND2x2_ASAP7_75t_L g3636 ( 
.A(n_2717),
.B(n_2724),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_2875),
.A2(n_3071),
.B(n_2928),
.Y(n_3637)
);

BUFx6f_ASAP7_75t_L g3638 ( 
.A(n_2083),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_L g3639 ( 
.A(n_2409),
.B(n_2662),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_2736),
.B(n_2740),
.Y(n_3640)
);

O2A1O1Ixp5_ASAP7_75t_L g3641 ( 
.A1(n_2549),
.A2(n_2623),
.B(n_2522),
.C(n_2684),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_2742),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_2875),
.A2(n_3071),
.B(n_2928),
.Y(n_3643)
);

OAI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2623),
.A2(n_2684),
.B(n_2729),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_2875),
.A2(n_2928),
.B(n_2923),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_2746),
.Y(n_3646)
);

AOI21x1_ASAP7_75t_L g3647 ( 
.A1(n_2758),
.A2(n_2766),
.B(n_3055),
.Y(n_3647)
);

INVxp67_ASAP7_75t_R g3648 ( 
.A(n_2295),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_2803),
.B(n_2804),
.Y(n_3649)
);

NOR2x1_ASAP7_75t_L g3650 ( 
.A(n_2097),
.B(n_2729),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2814),
.B(n_2815),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_2820),
.B(n_2823),
.Y(n_3652)
);

INVx1_ASAP7_75t_SL g3653 ( 
.A(n_2058),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_2861),
.B(n_2868),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_2083),
.B(n_2267),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3015),
.B(n_2465),
.Y(n_3656)
);

AOI21x1_ASAP7_75t_L g3657 ( 
.A1(n_2895),
.A2(n_2991),
.B(n_3029),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_2914),
.A2(n_2945),
.B(n_3028),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2919),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_2083),
.B(n_2756),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_2920),
.B(n_2932),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_2940),
.B(n_2947),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_2953),
.B(n_2969),
.Y(n_3663)
);

OAI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_2756),
.A2(n_3006),
.B(n_2989),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2993),
.B(n_3001),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_2067),
.A2(n_2439),
.B(n_2891),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_2067),
.A2(n_2439),
.B(n_2891),
.Y(n_3667)
);

INVx3_ASAP7_75t_L g3668 ( 
.A(n_2097),
.Y(n_3668)
);

O2A1O1Ixp5_ASAP7_75t_L g3669 ( 
.A1(n_2274),
.A2(n_2284),
.B(n_2287),
.C(n_2254),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_2983),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_2142),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_2067),
.A2(n_2439),
.B(n_2606),
.Y(n_3672)
);

OAI22xp5_ASAP7_75t_L g3673 ( 
.A1(n_2160),
.A2(n_2059),
.B1(n_3002),
.B2(n_2994),
.Y(n_3673)
);

NOR2xp67_ASAP7_75t_L g3674 ( 
.A(n_2241),
.B(n_2254),
.Y(n_3674)
);

NOR2xp67_ASAP7_75t_L g3675 ( 
.A(n_2241),
.B(n_2272),
.Y(n_3675)
);

OAI21xp5_ASAP7_75t_L g3676 ( 
.A1(n_2158),
.A2(n_2272),
.B(n_2002),
.Y(n_3676)
);

INVx3_ASAP7_75t_L g3677 ( 
.A(n_2606),
.Y(n_3677)
);

AOI33xp33_ASAP7_75t_L g3678 ( 
.A1(n_2490),
.A2(n_3059),
.A3(n_2963),
.B1(n_2530),
.B2(n_2540),
.B3(n_2572),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_2606),
.A2(n_2642),
.B(n_2891),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_1966),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_2642),
.A2(n_2166),
.B(n_2851),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_2642),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_2471),
.B(n_2860),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_2078),
.B(n_2175),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_2261),
.B(n_2277),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_1966),
.Y(n_3686)
);

AO21x1_ASAP7_75t_L g3687 ( 
.A1(n_2108),
.A2(n_2279),
.B(n_2196),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_2466),
.Y(n_3688)
);

BUFx8_ASAP7_75t_L g3689 ( 
.A(n_2491),
.Y(n_3689)
);

O2A1O1Ixp33_ASAP7_75t_L g3690 ( 
.A1(n_2647),
.A2(n_2929),
.B(n_2943),
.C(n_2931),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_2466),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_2269),
.A2(n_2211),
.B(n_2121),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2080),
.B(n_2117),
.Y(n_3693)
);

OAI22xp5_ASAP7_75t_L g3694 ( 
.A1(n_2470),
.A2(n_3042),
.B1(n_2734),
.B2(n_2876),
.Y(n_3694)
);

AOI21xp5_ASAP7_75t_L g3695 ( 
.A1(n_2269),
.A2(n_2470),
.B(n_3016),
.Y(n_3695)
);

A2O1A1Ixp33_ASAP7_75t_L g3696 ( 
.A1(n_1949),
.A2(n_2285),
.B(n_2162),
.C(n_2152),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3042),
.A2(n_3016),
.B(n_2990),
.Y(n_3697)
);

AOI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_2990),
.A2(n_2886),
.B(n_2876),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_SL g3699 ( 
.A(n_2734),
.B(n_2886),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_2108),
.B(n_2279),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_2073),
.A2(n_2196),
.B(n_2890),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_2661),
.B(n_2894),
.Y(n_3702)
);

AOI21x1_ASAP7_75t_L g3703 ( 
.A1(n_2464),
.A2(n_2807),
.B(n_2715),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_2680),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_2253),
.Y(n_3705)
);

INVx4_ASAP7_75t_L g3706 ( 
.A(n_2154),
.Y(n_3706)
);

NOR2xp67_ASAP7_75t_L g3707 ( 
.A(n_2169),
.B(n_2220),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_2483),
.Y(n_3708)
);

O2A1O1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_2483),
.A2(n_2544),
.B(n_2250),
.C(n_2264),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_2544),
.B(n_2631),
.Y(n_3710)
);

AOI21x1_ASAP7_75t_L g3711 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3711)
);

INVx2_ASAP7_75t_SL g3712 ( 
.A(n_2356),
.Y(n_3712)
);

NOR2xp67_ASAP7_75t_L g3713 ( 
.A(n_2007),
.B(n_2315),
.Y(n_3713)
);

INVxp67_ASAP7_75t_L g3714 ( 
.A(n_2004),
.Y(n_3714)
);

O2A1O1Ixp5_ASAP7_75t_L g3715 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_3715)
);

INVxp67_ASAP7_75t_SL g3716 ( 
.A(n_2631),
.Y(n_3716)
);

O2A1O1Ixp33_ASAP7_75t_L g3717 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3718)
);

A2O1A1Ixp33_ASAP7_75t_L g3719 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3719)
);

INVx1_ASAP7_75t_SL g3720 ( 
.A(n_2093),
.Y(n_3720)
);

BUFx2_ASAP7_75t_L g3721 ( 
.A(n_2631),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_2041),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3725)
);

INVx1_ASAP7_75t_SL g3726 ( 
.A(n_2093),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3728)
);

INVx3_ASAP7_75t_L g3729 ( 
.A(n_2893),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_2138),
.Y(n_3730)
);

AOI21x1_ASAP7_75t_L g3731 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3731)
);

AOI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3732)
);

INVx5_ASAP7_75t_L g3733 ( 
.A(n_2319),
.Y(n_3733)
);

NOR2x1_ASAP7_75t_L g3734 ( 
.A(n_2323),
.B(n_2334),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_2893),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3739)
);

AO21x1_ASAP7_75t_L g3740 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3740)
);

AO21x1_ASAP7_75t_L g3741 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3744)
);

CKINVDCx5p33_ASAP7_75t_R g3745 ( 
.A(n_2617),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_SL g3747 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3747)
);

AND2x4_ASAP7_75t_L g3748 ( 
.A(n_2103),
.B(n_2252),
.Y(n_3748)
);

OAI22xp5_ASAP7_75t_L g3749 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_L g3750 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3753)
);

OAI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3754)
);

OR2x2_ASAP7_75t_L g3755 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3756)
);

OAI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_L g3758 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3761)
);

INVx2_ASAP7_75t_SL g3762 ( 
.A(n_2356),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3767)
);

BUFx12f_ASAP7_75t_L g3768 ( 
.A(n_2283),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_SL g3772 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3772)
);

OAI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_2631),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3776)
);

OAI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3777)
);

OAI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3780)
);

OAI22xp5_ASAP7_75t_SL g3781 ( 
.A1(n_2611),
.A2(n_2304),
.B1(n_3054),
.B2(n_2716),
.Y(n_3781)
);

AND2x6_ASAP7_75t_SL g3782 ( 
.A(n_1923),
.B(n_1213),
.Y(n_3782)
);

INVx1_ASAP7_75t_SL g3783 ( 
.A(n_2093),
.Y(n_3783)
);

BUFx2_ASAP7_75t_L g3784 ( 
.A(n_2631),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3785)
);

OAI22xp5_ASAP7_75t_L g3786 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3788)
);

OAI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3792)
);

AOI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_2631),
.Y(n_3794)
);

NAND2x1_ASAP7_75t_L g3795 ( 
.A(n_2105),
.B(n_1494),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_2138),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3798)
);

AOI21x1_ASAP7_75t_L g3799 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3799)
);

NOR2xp67_ASAP7_75t_L g3800 ( 
.A(n_2007),
.B(n_2315),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3802)
);

AOI21x1_ASAP7_75t_L g3803 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_SL g3807 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3808)
);

BUFx4f_ASAP7_75t_L g3809 ( 
.A(n_2041),
.Y(n_3809)
);

A2O1A1Ixp33_ASAP7_75t_L g3810 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3811)
);

NOR3xp33_ASAP7_75t_L g3812 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3813)
);

HB1xp67_ASAP7_75t_L g3814 ( 
.A(n_2356),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3815)
);

A2O1A1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3816)
);

OAI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3818)
);

AOI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2294),
.B(n_2297),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3821)
);

O2A1O1Ixp33_ASAP7_75t_L g3822 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3823)
);

BUFx6f_ASAP7_75t_L g3824 ( 
.A(n_2041),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3825)
);

OAI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3835)
);

BUFx3_ASAP7_75t_L g3836 ( 
.A(n_2068),
.Y(n_3836)
);

INVx3_ASAP7_75t_L g3837 ( 
.A(n_2893),
.Y(n_3837)
);

NOR3xp33_ASAP7_75t_L g3838 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_3838)
);

AOI21xp33_ASAP7_75t_L g3839 ( 
.A1(n_2005),
.A2(n_2334),
.B(n_2323),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3843)
);

INVx1_ASAP7_75t_SL g3844 ( 
.A(n_2093),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3845)
);

OAI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_SL g3848 ( 
.A(n_2040),
.B(n_2017),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3850)
);

INVx1_ASAP7_75t_SL g3851 ( 
.A(n_2093),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_2138),
.Y(n_3856)
);

NOR3xp33_ASAP7_75t_L g3857 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_2138),
.Y(n_3858)
);

OAI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3859)
);

BUFx4f_ASAP7_75t_L g3860 ( 
.A(n_2041),
.Y(n_3860)
);

CKINVDCx20_ASAP7_75t_R g3861 ( 
.A(n_2257),
.Y(n_3861)
);

INVx4_ASAP7_75t_L g3862 ( 
.A(n_2041),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_2138),
.Y(n_3863)
);

O2A1O1Ixp5_ASAP7_75t_L g3864 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_3864)
);

BUFx3_ASAP7_75t_L g3865 ( 
.A(n_2068),
.Y(n_3865)
);

AND2x4_ASAP7_75t_L g3866 ( 
.A(n_2103),
.B(n_2252),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3868)
);

OAI22xp5_ASAP7_75t_L g3869 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3869)
);

O2A1O1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_2138),
.Y(n_3871)
);

O2A1O1Ixp33_ASAP7_75t_L g3872 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3872)
);

AOI21xp33_ASAP7_75t_L g3873 ( 
.A1(n_2005),
.A2(n_2334),
.B(n_2323),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3875)
);

O2A1O1Ixp33_ASAP7_75t_L g3876 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_SL g3879 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3879)
);

OR2x2_ASAP7_75t_SL g3880 ( 
.A(n_2337),
.B(n_2810),
.Y(n_3880)
);

BUFx12f_ASAP7_75t_L g3881 ( 
.A(n_2283),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3883)
);

INVx1_ASAP7_75t_SL g3884 ( 
.A(n_2093),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3885)
);

INVx2_ASAP7_75t_SL g3886 ( 
.A(n_2356),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_2893),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3889)
);

OAI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_L g3895 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3895)
);

O2A1O1Ixp5_ASAP7_75t_L g3896 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3899)
);

INVx3_ASAP7_75t_L g3900 ( 
.A(n_2893),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_2138),
.Y(n_3901)
);

NOR2xp33_ASAP7_75t_L g3902 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3907)
);

OAI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3909)
);

O2A1O1Ixp33_ASAP7_75t_L g3910 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_L g3913 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3913)
);

BUFx2_ASAP7_75t_L g3914 ( 
.A(n_2631),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3916)
);

OR2x6_ASAP7_75t_L g3917 ( 
.A(n_2069),
.B(n_2105),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3918)
);

NOR2xp67_ASAP7_75t_L g3919 ( 
.A(n_2007),
.B(n_2315),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_2138),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_2138),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3922)
);

NAND2x1_ASAP7_75t_L g3923 ( 
.A(n_2105),
.B(n_1494),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_2893),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3926)
);

OAI22xp5_ASAP7_75t_L g3927 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3927)
);

O2A1O1Ixp33_ASAP7_75t_L g3928 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3930)
);

NOR2xp67_ASAP7_75t_L g3931 ( 
.A(n_2007),
.B(n_2315),
.Y(n_3931)
);

AOI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3932)
);

AO21x1_ASAP7_75t_L g3933 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3933)
);

OR2x2_ASAP7_75t_L g3934 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3935)
);

HB1xp67_ASAP7_75t_L g3936 ( 
.A(n_2356),
.Y(n_3936)
);

AOI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3938)
);

NOR2x1_ASAP7_75t_L g3939 ( 
.A(n_2323),
.B(n_2334),
.Y(n_3939)
);

NOR2xp33_ASAP7_75t_L g3940 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3940)
);

CKINVDCx10_ASAP7_75t_R g3941 ( 
.A(n_2664),
.Y(n_3941)
);

A2O1A1Ixp33_ASAP7_75t_L g3942 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3942)
);

CKINVDCx5p33_ASAP7_75t_R g3943 ( 
.A(n_2617),
.Y(n_3943)
);

OAI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3944)
);

OAI21x1_ASAP7_75t_L g3945 ( 
.A1(n_2105),
.A2(n_1434),
.B(n_2043),
.Y(n_3945)
);

NOR2xp33_ASAP7_75t_SL g3946 ( 
.A(n_2040),
.B(n_2017),
.Y(n_3946)
);

O2A1O1Ixp5_ASAP7_75t_L g3947 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3949)
);

BUFx4f_ASAP7_75t_L g3950 ( 
.A(n_2041),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_2138),
.Y(n_3955)
);

AOI21x1_ASAP7_75t_L g3956 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3956)
);

AOI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3957)
);

INVx3_ASAP7_75t_L g3958 ( 
.A(n_2893),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3960)
);

OR2x2_ASAP7_75t_L g3961 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3961)
);

AOI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_844),
.B2(n_1249),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3964)
);

OAI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3966)
);

AOI21x1_ASAP7_75t_L g3967 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_2510),
.B(n_2827),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3971)
);

A2O1A1Ixp33_ASAP7_75t_L g3972 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3972)
);

INVxp67_ASAP7_75t_L g3973 ( 
.A(n_2004),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3974)
);

AND2x2_ASAP7_75t_SL g3975 ( 
.A(n_1914),
.B(n_2041),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_2138),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3978)
);

AO21x1_ASAP7_75t_L g3979 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_3979)
);

AOI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3980)
);

AOI21xp5_ASAP7_75t_SL g3981 ( 
.A1(n_2631),
.A2(n_2788),
.B(n_2745),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3982)
);

NAND3xp33_ASAP7_75t_SL g3983 ( 
.A(n_2453),
.B(n_2501),
.C(n_2420),
.Y(n_3983)
);

AO21x2_ASAP7_75t_L g3984 ( 
.A1(n_2069),
.A2(n_2745),
.B(n_2631),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3986)
);

OAI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3992)
);

A2O1A1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_3993)
);

OAI22xp5_ASAP7_75t_L g3994 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3995)
);

NOR2xp33_ASAP7_75t_L g3996 ( 
.A(n_1923),
.B(n_2300),
.Y(n_3996)
);

BUFx2_ASAP7_75t_L g3997 ( 
.A(n_2631),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_2631),
.B(n_2745),
.Y(n_3998)
);

NAND2xp33_ASAP7_75t_L g3999 ( 
.A(n_2065),
.B(n_2420),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_L g4000 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4000)
);

OR2x2_ASAP7_75t_L g4001 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4002)
);

O2A1O1Ixp5_ASAP7_75t_L g4003 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4004)
);

OAI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4007)
);

INVxp67_ASAP7_75t_SL g4008 ( 
.A(n_2631),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4009)
);

OAI321xp33_ASAP7_75t_L g4010 ( 
.A1(n_1918),
.A2(n_2373),
.A3(n_2369),
.B1(n_2406),
.B2(n_2390),
.C(n_2367),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4011)
);

OAI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4012)
);

INVx4_ASAP7_75t_L g4013 ( 
.A(n_2041),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4014)
);

OAI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4015)
);

AO21x2_ASAP7_75t_L g4016 ( 
.A1(n_2069),
.A2(n_2745),
.B(n_2631),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_2138),
.Y(n_4018)
);

OAI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4019)
);

INVx1_ASAP7_75t_SL g4020 ( 
.A(n_2093),
.Y(n_4020)
);

A2O1A1Ixp33_ASAP7_75t_L g4021 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4023)
);

AND2x4_ASAP7_75t_L g4024 ( 
.A(n_2103),
.B(n_2252),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4028)
);

O2A1O1Ixp33_ASAP7_75t_L g4029 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4029)
);

A2O1A1Ixp33_ASAP7_75t_L g4030 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4030)
);

AOI21xp5_ASAP7_75t_L g4031 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4031)
);

INVxp67_ASAP7_75t_L g4032 ( 
.A(n_2004),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_SL g4034 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4035)
);

AOI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4036)
);

OAI22xp5_ASAP7_75t_L g4037 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4037)
);

BUFx6f_ASAP7_75t_L g4038 ( 
.A(n_2041),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_2138),
.Y(n_4039)
);

BUFx2_ASAP7_75t_L g4040 ( 
.A(n_2631),
.Y(n_4040)
);

OAI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4041)
);

AOI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4042)
);

BUFx6f_ASAP7_75t_L g4043 ( 
.A(n_2041),
.Y(n_4043)
);

AOI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4045)
);

A2O1A1Ixp33_ASAP7_75t_L g4046 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4046)
);

CKINVDCx6p67_ASAP7_75t_R g4047 ( 
.A(n_2305),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4051)
);

NAND2x1p5_ASAP7_75t_L g4052 ( 
.A(n_2041),
.B(n_2893),
.Y(n_4052)
);

BUFx3_ASAP7_75t_L g4053 ( 
.A(n_2068),
.Y(n_4053)
);

BUFx8_ASAP7_75t_L g4054 ( 
.A(n_2664),
.Y(n_4054)
);

AOI33xp33_ASAP7_75t_L g4055 ( 
.A1(n_2300),
.A2(n_2372),
.A3(n_2317),
.B1(n_2387),
.B2(n_2325),
.B3(n_2311),
.Y(n_4055)
);

AOI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4056)
);

INVxp67_ASAP7_75t_L g4057 ( 
.A(n_2004),
.Y(n_4057)
);

NOR3xp33_ASAP7_75t_L g4058 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4058)
);

AO21x1_ASAP7_75t_L g4059 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4059)
);

A2O1A1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4062)
);

AOI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4063)
);

AOI21xp5_ASAP7_75t_L g4064 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4064)
);

AOI21xp5_ASAP7_75t_L g4065 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4065)
);

NAND2x1p5_ASAP7_75t_L g4066 ( 
.A(n_2041),
.B(n_2893),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4067)
);

AOI21xp5_ASAP7_75t_L g4068 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4068)
);

NOR2xp33_ASAP7_75t_L g4069 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4070)
);

AOI21xp5_ASAP7_75t_L g4071 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_844),
.B2(n_1249),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4073)
);

OR2x6_ASAP7_75t_L g4074 ( 
.A(n_2069),
.B(n_2105),
.Y(n_4074)
);

O2A1O1Ixp33_ASAP7_75t_L g4075 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_2138),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4080)
);

OAI21xp33_ASAP7_75t_L g4081 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2300),
.Y(n_4081)
);

BUFx3_ASAP7_75t_L g4082 ( 
.A(n_2068),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_844),
.B2(n_1249),
.Y(n_4083)
);

AOI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4084)
);

AOI33xp33_ASAP7_75t_L g4085 ( 
.A1(n_2300),
.A2(n_2372),
.A3(n_2317),
.B1(n_2387),
.B2(n_2325),
.B3(n_2311),
.Y(n_4085)
);

INVx11_ASAP7_75t_L g4086 ( 
.A(n_2153),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4089)
);

AOI21xp33_ASAP7_75t_L g4090 ( 
.A1(n_2005),
.A2(n_2334),
.B(n_2323),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_2138),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_SL g4093 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4094)
);

NOR2x2_ASAP7_75t_L g4095 ( 
.A(n_2419),
.B(n_1496),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4096)
);

BUFx4f_ASAP7_75t_L g4097 ( 
.A(n_2041),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_2041),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4099)
);

CKINVDCx5p33_ASAP7_75t_R g4100 ( 
.A(n_2617),
.Y(n_4100)
);

NOR3xp33_ASAP7_75t_L g4101 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4102)
);

NOR2xp33_ASAP7_75t_L g4103 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4103)
);

BUFx4f_ASAP7_75t_L g4104 ( 
.A(n_2041),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4105)
);

OAI21xp33_ASAP7_75t_L g4106 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2300),
.Y(n_4106)
);

INVxp67_ASAP7_75t_L g4107 ( 
.A(n_2004),
.Y(n_4107)
);

O2A1O1Ixp33_ASAP7_75t_L g4108 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4109)
);

AOI21x1_ASAP7_75t_L g4110 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4111)
);

AND2x4_ASAP7_75t_L g4112 ( 
.A(n_2103),
.B(n_2252),
.Y(n_4112)
);

AOI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4115)
);

NOR2xp67_ASAP7_75t_L g4116 ( 
.A(n_2007),
.B(n_2315),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_L g4117 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4118)
);

BUFx6f_ASAP7_75t_L g4119 ( 
.A(n_2041),
.Y(n_4119)
);

AND2x2_ASAP7_75t_SL g4120 ( 
.A(n_1914),
.B(n_2041),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4122)
);

O2A1O1Ixp33_ASAP7_75t_SL g4123 ( 
.A1(n_2040),
.A2(n_2430),
.B(n_2859),
.C(n_2328),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4125)
);

AOI22x1_ASAP7_75t_L g4126 ( 
.A1(n_2454),
.A2(n_2925),
.B1(n_2315),
.B2(n_2498),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4127)
);

OAI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4129)
);

BUFx8_ASAP7_75t_L g4130 ( 
.A(n_2664),
.Y(n_4130)
);

A2O1A1Ixp33_ASAP7_75t_L g4131 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4135)
);

A2O1A1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4137)
);

NOR2xp33_ASAP7_75t_L g4138 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4138)
);

OAI21xp33_ASAP7_75t_L g4139 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2300),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4141)
);

O2A1O1Ixp33_ASAP7_75t_L g4142 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4142)
);

INVx11_ASAP7_75t_L g4143 ( 
.A(n_2153),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4145)
);

NOR3xp33_ASAP7_75t_L g4146 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4149)
);

INVx3_ASAP7_75t_L g4150 ( 
.A(n_2893),
.Y(n_4150)
);

O2A1O1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4151)
);

AOI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4153)
);

AOI21xp5_ASAP7_75t_L g4154 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4154)
);

NOR3xp33_ASAP7_75t_L g4155 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4155)
);

HB1xp67_ASAP7_75t_L g4156 ( 
.A(n_2356),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4157)
);

BUFx8_ASAP7_75t_L g4158 ( 
.A(n_2664),
.Y(n_4158)
);

A2O1A1Ixp33_ASAP7_75t_L g4159 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4159)
);

AOI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4161)
);

NAND2x1p5_ASAP7_75t_L g4162 ( 
.A(n_2041),
.B(n_2893),
.Y(n_4162)
);

AOI21xp5_ASAP7_75t_L g4163 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4164)
);

O2A1O1Ixp33_ASAP7_75t_L g4165 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4166)
);

A2O1A1Ixp33_ASAP7_75t_L g4167 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4168)
);

INVx4_ASAP7_75t_L g4169 ( 
.A(n_2041),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_2138),
.Y(n_4170)
);

HB1xp67_ASAP7_75t_L g4171 ( 
.A(n_2356),
.Y(n_4171)
);

NOR2xp33_ASAP7_75t_L g4172 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4173)
);

NOR2x1p5_ASAP7_75t_L g4174 ( 
.A(n_2893),
.B(n_2337),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_L g4175 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4176)
);

OAI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4177)
);

BUFx4f_ASAP7_75t_L g4178 ( 
.A(n_2041),
.Y(n_4178)
);

AOI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_4179)
);

AOI21xp5_ASAP7_75t_L g4180 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_2138),
.Y(n_4181)
);

AOI21xp5_ASAP7_75t_L g4182 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4182)
);

NOR2xp33_ASAP7_75t_L g4183 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4184)
);

AND2x2_ASAP7_75t_L g4185 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_R g4186 ( 
.A(n_2650),
.B(n_466),
.Y(n_4186)
);

INVxp67_ASAP7_75t_L g4187 ( 
.A(n_2004),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4188)
);

AOI21xp5_ASAP7_75t_L g4189 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_2138),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4192)
);

AOI21xp33_ASAP7_75t_L g4193 ( 
.A1(n_2005),
.A2(n_2334),
.B(n_2323),
.Y(n_4193)
);

NOR2xp33_ASAP7_75t_L g4194 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4197)
);

CKINVDCx10_ASAP7_75t_R g4198 ( 
.A(n_2664),
.Y(n_4198)
);

BUFx6f_ASAP7_75t_L g4199 ( 
.A(n_2041),
.Y(n_4199)
);

INVxp67_ASAP7_75t_L g4200 ( 
.A(n_2004),
.Y(n_4200)
);

AND2x6_ASAP7_75t_L g4201 ( 
.A(n_2103),
.B(n_2319),
.Y(n_4201)
);

AOI21xp5_ASAP7_75t_L g4202 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_2138),
.Y(n_4203)
);

NAND3xp33_ASAP7_75t_L g4204 ( 
.A(n_2420),
.B(n_2636),
.C(n_2501),
.Y(n_4204)
);

AOI21xp5_ASAP7_75t_L g4205 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_2068),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_SL g4207 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_2138),
.Y(n_4209)
);

A2O1A1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4210)
);

NOR3xp33_ASAP7_75t_L g4211 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4217)
);

AO21x1_ASAP7_75t_L g4218 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4218)
);

AOI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4220)
);

AOI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4223)
);

A2O1A1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4224)
);

AOI21xp5_ASAP7_75t_L g4225 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4225)
);

O2A1O1Ixp33_ASAP7_75t_SL g4226 ( 
.A1(n_2040),
.A2(n_2430),
.B(n_2859),
.C(n_2328),
.Y(n_4226)
);

INVx3_ASAP7_75t_L g4227 ( 
.A(n_2893),
.Y(n_4227)
);

OAI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4229)
);

AOI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4230)
);

NAND3xp33_ASAP7_75t_SL g4231 ( 
.A(n_2453),
.B(n_2501),
.C(n_2420),
.Y(n_4231)
);

BUFx8_ASAP7_75t_L g4232 ( 
.A(n_2664),
.Y(n_4232)
);

AOI21xp33_ASAP7_75t_L g4233 ( 
.A1(n_2005),
.A2(n_2334),
.B(n_2323),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4234)
);

O2A1O1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_2138),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4241)
);

OAI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4242)
);

OAI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_2631),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_2631),
.Y(n_4245)
);

INVx4_ASAP7_75t_L g4246 ( 
.A(n_2041),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4247)
);

INVx2_ASAP7_75t_SL g4248 ( 
.A(n_2356),
.Y(n_4248)
);

NOR3xp33_ASAP7_75t_L g4249 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_2138),
.Y(n_4250)
);

NOR2xp67_ASAP7_75t_L g4251 ( 
.A(n_2007),
.B(n_2315),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_2138),
.Y(n_4252)
);

AO21x1_ASAP7_75t_L g4253 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_2631),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4256)
);

NOR2xp33_ASAP7_75t_L g4257 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_SL g4258 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4258)
);

AO21x1_ASAP7_75t_L g4259 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_2631),
.Y(n_4260)
);

NOR3xp33_ASAP7_75t_L g4261 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4261)
);

NOR2xp33_ASAP7_75t_L g4262 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4262)
);

INVx4_ASAP7_75t_L g4263 ( 
.A(n_2041),
.Y(n_4263)
);

AO21x1_ASAP7_75t_L g4264 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4264)
);

A2O1A1Ixp33_ASAP7_75t_L g4265 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_2631),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4268)
);

NOR2xp33_ASAP7_75t_L g4269 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_SL g4270 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_SL g4271 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_2631),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_SL g4273 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4274)
);

INVx2_ASAP7_75t_SL g4275 ( 
.A(n_2356),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_2631),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_2631),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4278)
);

AOI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_4279)
);

INVx1_ASAP7_75t_SL g4280 ( 
.A(n_2093),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_SL g4282 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4282)
);

INVx2_ASAP7_75t_SL g4283 ( 
.A(n_2356),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_SL g4285 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_2138),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4287)
);

INVx2_ASAP7_75t_SL g4288 ( 
.A(n_2356),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_SL g4292 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_SL g4293 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4294)
);

OAI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4295)
);

INVx3_ASAP7_75t_L g4296 ( 
.A(n_2893),
.Y(n_4296)
);

INVx3_ASAP7_75t_L g4297 ( 
.A(n_2893),
.Y(n_4297)
);

NOR2x1p5_ASAP7_75t_SL g4298 ( 
.A(n_2138),
.B(n_1470),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_SL g4299 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4300)
);

OAI22xp5_ASAP7_75t_L g4301 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_2041),
.Y(n_4303)
);

O2A1O1Ixp33_ASAP7_75t_L g4304 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4304)
);

OAI321xp33_ASAP7_75t_L g4305 ( 
.A1(n_1918),
.A2(n_2373),
.A3(n_2369),
.B1(n_2406),
.B2(n_2390),
.C(n_2367),
.Y(n_4305)
);

AOI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_2138),
.Y(n_4307)
);

HB1xp67_ASAP7_75t_L g4308 ( 
.A(n_2356),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_2631),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_2138),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4313)
);

CKINVDCx10_ASAP7_75t_R g4314 ( 
.A(n_2664),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4315)
);

O2A1O1Ixp33_ASAP7_75t_SL g4316 ( 
.A1(n_2040),
.A2(n_2430),
.B(n_2859),
.C(n_2328),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4317)
);

BUFx12f_ASAP7_75t_L g4318 ( 
.A(n_2283),
.Y(n_4318)
);

A2O1A1Ixp33_ASAP7_75t_L g4319 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_L g4320 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4321)
);

INVx3_ASAP7_75t_L g4322 ( 
.A(n_2893),
.Y(n_4322)
);

OAI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4323)
);

NOR3xp33_ASAP7_75t_L g4324 ( 
.A(n_2453),
.B(n_2810),
.C(n_2337),
.Y(n_4324)
);

AOI21x1_ASAP7_75t_L g4325 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4325)
);

OR2x6_ASAP7_75t_L g4326 ( 
.A(n_2069),
.B(n_2105),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4327)
);

NAND2xp33_ASAP7_75t_L g4328 ( 
.A(n_2065),
.B(n_2420),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4329)
);

AOI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4331)
);

O2A1O1Ixp5_ASAP7_75t_L g4332 ( 
.A1(n_2291),
.A2(n_2331),
.B(n_2040),
.C(n_1923),
.Y(n_4332)
);

NOR2x1_ASAP7_75t_R g4333 ( 
.A(n_2305),
.B(n_378),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_2631),
.Y(n_4336)
);

NOR2xp33_ASAP7_75t_L g4337 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_2138),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4340)
);

OAI21xp33_ASAP7_75t_SL g4341 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4345)
);

AO21x1_ASAP7_75t_L g4346 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_2138),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_SL g4349 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4349)
);

INVx11_ASAP7_75t_L g4350 ( 
.A(n_2153),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_2631),
.Y(n_4351)
);

AOI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_2294),
.A2(n_2297),
.B1(n_2329),
.B2(n_2316),
.Y(n_4352)
);

AO21x1_ASAP7_75t_L g4353 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_2631),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4355)
);

A2O1A1Ixp33_ASAP7_75t_L g4356 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4356)
);

A2O1A1Ixp33_ASAP7_75t_L g4357 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4357)
);

A2O1A1Ixp33_ASAP7_75t_L g4358 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4358)
);

BUFx3_ASAP7_75t_L g4359 ( 
.A(n_2068),
.Y(n_4359)
);

AND2x6_ASAP7_75t_L g4360 ( 
.A(n_2103),
.B(n_2319),
.Y(n_4360)
);

CKINVDCx5p33_ASAP7_75t_R g4361 ( 
.A(n_2617),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4363)
);

NOR2xp33_ASAP7_75t_L g4364 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4364)
);

AOI22xp33_ASAP7_75t_L g4365 ( 
.A1(n_2624),
.A2(n_1976),
.B1(n_844),
.B2(n_1249),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_2356),
.Y(n_4367)
);

AOI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4368)
);

AOI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4369)
);

BUFx6f_ASAP7_75t_L g4370 ( 
.A(n_2041),
.Y(n_4370)
);

OAI21x1_ASAP7_75t_L g4371 ( 
.A1(n_2105),
.A2(n_1434),
.B(n_2043),
.Y(n_4371)
);

INVxp67_ASAP7_75t_L g4372 ( 
.A(n_2004),
.Y(n_4372)
);

AOI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4373)
);

BUFx4f_ASAP7_75t_L g4374 ( 
.A(n_2041),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_2138),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4376)
);

AOI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4377)
);

AOI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_2631),
.Y(n_4379)
);

AOI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4382)
);

INVx1_ASAP7_75t_SL g4383 ( 
.A(n_2093),
.Y(n_4383)
);

A2O1A1Ixp33_ASAP7_75t_L g4384 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4387)
);

OAI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_2631),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4390)
);

OAI22xp5_ASAP7_75t_L g4391 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4392)
);

AO21x2_ASAP7_75t_L g4393 ( 
.A1(n_2069),
.A2(n_2745),
.B(n_2631),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4394)
);

AOI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_SL g4398 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4399)
);

AOI21xp5_ASAP7_75t_L g4400 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4400)
);

A2O1A1Ixp33_ASAP7_75t_L g4401 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_2631),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4404)
);

AOI21xp5_ASAP7_75t_L g4405 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_2631),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_L g4409 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4410)
);

NOR2xp33_ASAP7_75t_L g4411 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4412)
);

INVx11_ASAP7_75t_L g4413 ( 
.A(n_2153),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_2631),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4415)
);

NOR2xp67_ASAP7_75t_L g4416 ( 
.A(n_2007),
.B(n_2315),
.Y(n_4416)
);

A2O1A1Ixp33_ASAP7_75t_L g4417 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4419)
);

HB1xp67_ASAP7_75t_L g4420 ( 
.A(n_2356),
.Y(n_4420)
);

AOI21xp5_ASAP7_75t_L g4421 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_2631),
.Y(n_4422)
);

AOI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_2631),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4426)
);

O2A1O1Ixp33_ASAP7_75t_L g4427 ( 
.A1(n_2040),
.A2(n_2304),
.B(n_2810),
.C(n_2337),
.Y(n_4427)
);

BUFx6f_ASAP7_75t_L g4428 ( 
.A(n_2041),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_2631),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_SL g4430 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_2631),
.Y(n_4431)
);

OAI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4432)
);

OAI21xp5_ASAP7_75t_L g4433 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4433)
);

AOI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4434)
);

AOI21xp5_ASAP7_75t_L g4435 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4435)
);

AOI21xp5_ASAP7_75t_L g4436 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4436)
);

AOI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4439)
);

AOI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4440)
);

AOI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4441)
);

CKINVDCx6p67_ASAP7_75t_R g4442 ( 
.A(n_2305),
.Y(n_4442)
);

BUFx2_ASAP7_75t_L g4443 ( 
.A(n_2631),
.Y(n_4443)
);

NOR2xp33_ASAP7_75t_L g4444 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4444)
);

HB1xp67_ASAP7_75t_L g4445 ( 
.A(n_2356),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_2631),
.Y(n_4446)
);

AND2x2_ASAP7_75t_L g4447 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4447)
);

BUFx12f_ASAP7_75t_L g4448 ( 
.A(n_2283),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4449)
);

AND2x4_ASAP7_75t_L g4450 ( 
.A(n_2103),
.B(n_2252),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_SL g4451 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4451)
);

AOI21x1_ASAP7_75t_L g4452 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4452)
);

OAI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_2301),
.A2(n_2627),
.B(n_2432),
.Y(n_4453)
);

AOI21xp5_ASAP7_75t_L g4454 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4455)
);

AOI21x1_ASAP7_75t_L g4456 ( 
.A1(n_2323),
.A2(n_2509),
.B(n_2334),
.Y(n_4456)
);

BUFx4f_ASAP7_75t_L g4457 ( 
.A(n_2041),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4459)
);

INVx3_ASAP7_75t_L g4460 ( 
.A(n_2893),
.Y(n_4460)
);

AOI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4461)
);

A2O1A1Ixp33_ASAP7_75t_L g4462 ( 
.A1(n_2040),
.A2(n_2453),
.B(n_2017),
.C(n_2055),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_SL g4463 ( 
.A(n_2510),
.B(n_2827),
.Y(n_4463)
);

AO22x1_ASAP7_75t_L g4464 ( 
.A1(n_2065),
.A2(n_2084),
.B1(n_1249),
.B2(n_2061),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_2631),
.B(n_2745),
.Y(n_4465)
);

OAI21xp33_ASAP7_75t_L g4466 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2300),
.Y(n_4466)
);

INVx3_ASAP7_75t_L g4467 ( 
.A(n_2893),
.Y(n_4467)
);

AOI21xp5_ASAP7_75t_L g4468 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4468)
);

NOR2xp33_ASAP7_75t_L g4469 ( 
.A(n_1923),
.B(n_2300),
.Y(n_4469)
);

AOI21xp5_ASAP7_75t_L g4470 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_2138),
.Y(n_4472)
);

OAI22xp5_ASAP7_75t_L g4473 ( 
.A1(n_2300),
.A2(n_2317),
.B1(n_2325),
.B2(n_2311),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_2294),
.B(n_2297),
.Y(n_4474)
);

AOI21xp5_ASAP7_75t_L g4475 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_2315),
.A2(n_2498),
.B(n_2327),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_3076),
.B(n_3757),
.Y(n_4477)
);

AND2x6_ASAP7_75t_L g4478 ( 
.A(n_3722),
.B(n_3824),
.Y(n_4478)
);

OAI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_3145),
.A2(n_3164),
.B1(n_3160),
.B2(n_3126),
.Y(n_4479)
);

OR2x6_ASAP7_75t_L g4480 ( 
.A(n_3981),
.B(n_3795),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_SL g4481 ( 
.A(n_3076),
.B(n_3757),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_3074),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3074),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_3081),
.Y(n_4484)
);

BUFx6f_ASAP7_75t_L g4485 ( 
.A(n_3123),
.Y(n_4485)
);

AND2x4_ASAP7_75t_L g4486 ( 
.A(n_3123),
.B(n_3206),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_3081),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_3130),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_3130),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_3724),
.Y(n_4490)
);

INVx3_ASAP7_75t_L g4491 ( 
.A(n_3167),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_3130),
.Y(n_4492)
);

A2O1A1Ixp33_ASAP7_75t_L g4493 ( 
.A1(n_4341),
.A2(n_3717),
.B(n_3870),
.C(n_3822),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_3140),
.Y(n_4494)
);

INVx3_ASAP7_75t_L g4495 ( 
.A(n_3167),
.Y(n_4495)
);

INVx2_ASAP7_75t_SL g4496 ( 
.A(n_3123),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_3140),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_3083),
.B(n_3090),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_3083),
.B(n_3090),
.Y(n_4499)
);

BUFx3_ASAP7_75t_L g4500 ( 
.A(n_3206),
.Y(n_4500)
);

OR2x2_ASAP7_75t_SL g4501 ( 
.A(n_3092),
.B(n_3104),
.Y(n_4501)
);

BUFx2_ASAP7_75t_L g4502 ( 
.A(n_3721),
.Y(n_4502)
);

INVx2_ASAP7_75t_SL g4503 ( 
.A(n_3206),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3092),
.B(n_3342),
.Y(n_4504)
);

AND2x4_ASAP7_75t_L g4505 ( 
.A(n_3325),
.B(n_3368),
.Y(n_4505)
);

BUFx3_ASAP7_75t_L g4506 ( 
.A(n_3325),
.Y(n_4506)
);

BUFx6f_ASAP7_75t_L g4507 ( 
.A(n_3325),
.Y(n_4507)
);

BUFx6f_ASAP7_75t_L g4508 ( 
.A(n_3368),
.Y(n_4508)
);

BUFx2_ASAP7_75t_L g4509 ( 
.A(n_3721),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_3345),
.B(n_3350),
.Y(n_4510)
);

BUFx4f_ASAP7_75t_L g4511 ( 
.A(n_4201),
.Y(n_4511)
);

BUFx3_ASAP7_75t_L g4512 ( 
.A(n_3368),
.Y(n_4512)
);

NOR2x1_ASAP7_75t_L g4513 ( 
.A(n_3093),
.B(n_3734),
.Y(n_4513)
);

OAI31xp33_ASAP7_75t_SL g4514 ( 
.A1(n_3777),
.A2(n_3817),
.A3(n_3846),
.B(n_3778),
.Y(n_4514)
);

OR2x6_ASAP7_75t_L g4515 ( 
.A(n_3981),
.B(n_3795),
.Y(n_4515)
);

INVx3_ASAP7_75t_L g4516 ( 
.A(n_3271),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_3271),
.Y(n_4517)
);

BUFx6f_ASAP7_75t_L g4518 ( 
.A(n_3480),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_SL g4519 ( 
.A(n_3777),
.B(n_3778),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_3104),
.B(n_3817),
.Y(n_4520)
);

BUFx12f_ASAP7_75t_L g4521 ( 
.A(n_4054),
.Y(n_4521)
);

AND2x4_ASAP7_75t_L g4522 ( 
.A(n_3480),
.B(n_3836),
.Y(n_4522)
);

BUFx2_ASAP7_75t_L g4523 ( 
.A(n_3784),
.Y(n_4523)
);

AND2x2_ASAP7_75t_SL g4524 ( 
.A(n_3809),
.B(n_3860),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3724),
.Y(n_4525)
);

BUFx4f_ASAP7_75t_L g4526 ( 
.A(n_4201),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_3846),
.B(n_3890),
.Y(n_4527)
);

AND2x4_ASAP7_75t_L g4528 ( 
.A(n_3480),
.B(n_3836),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_3725),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3725),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_3784),
.Y(n_4531)
);

BUFx6f_ASAP7_75t_L g4532 ( 
.A(n_3836),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_SL g4533 ( 
.A(n_3890),
.B(n_3905),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_3079),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3728),
.Y(n_4535)
);

BUFx2_ASAP7_75t_L g4536 ( 
.A(n_3914),
.Y(n_4536)
);

CKINVDCx5p33_ASAP7_75t_R g4537 ( 
.A(n_4186),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3905),
.B(n_3908),
.Y(n_4538)
);

OAI22xp5_ASAP7_75t_L g4539 ( 
.A1(n_3122),
.A2(n_3128),
.B1(n_3727),
.B2(n_3126),
.Y(n_4539)
);

BUFx6f_ASAP7_75t_L g4540 ( 
.A(n_3865),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_3908),
.B(n_3909),
.Y(n_4541)
);

AOI22xp33_ASAP7_75t_L g4542 ( 
.A1(n_3155),
.A2(n_3163),
.B1(n_4106),
.B2(n_4081),
.Y(n_4542)
);

BUFx2_ASAP7_75t_L g4543 ( 
.A(n_3914),
.Y(n_4543)
);

AOI21xp5_ASAP7_75t_L g4544 ( 
.A1(n_3072),
.A2(n_3088),
.B(n_3086),
.Y(n_4544)
);

BUFx3_ASAP7_75t_L g4545 ( 
.A(n_3865),
.Y(n_4545)
);

BUFx2_ASAP7_75t_L g4546 ( 
.A(n_3997),
.Y(n_4546)
);

NOR2xp67_ASAP7_75t_L g4547 ( 
.A(n_3181),
.B(n_3182),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3909),
.B(n_3965),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_3965),
.B(n_3987),
.Y(n_4549)
);

BUFx3_ASAP7_75t_L g4550 ( 
.A(n_3865),
.Y(n_4550)
);

BUFx3_ASAP7_75t_L g4551 ( 
.A(n_4053),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_3188),
.B(n_3718),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_3728),
.Y(n_4553)
);

A2O1A1Ixp33_ASAP7_75t_L g4554 ( 
.A1(n_4341),
.A2(n_3876),
.B(n_3910),
.C(n_3872),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_3987),
.B(n_4009),
.Y(n_4555)
);

AND2x4_ASAP7_75t_L g4556 ( 
.A(n_4053),
.B(n_4082),
.Y(n_4556)
);

NAND2x1p5_ASAP7_75t_L g4557 ( 
.A(n_3923),
.B(n_3093),
.Y(n_4557)
);

CKINVDCx20_ASAP7_75t_R g4558 ( 
.A(n_3080),
.Y(n_4558)
);

BUFx12f_ASAP7_75t_L g4559 ( 
.A(n_4054),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4009),
.B(n_4012),
.Y(n_4560)
);

NAND2x1p5_ASAP7_75t_L g4561 ( 
.A(n_3923),
.B(n_3734),
.Y(n_4561)
);

INVxp67_ASAP7_75t_L g4562 ( 
.A(n_3736),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_4012),
.B(n_4015),
.Y(n_4563)
);

INVxp67_ASAP7_75t_L g4564 ( 
.A(n_3736),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4015),
.B(n_4041),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_SL g4566 ( 
.A(n_4041),
.B(n_4128),
.Y(n_4566)
);

AND3x1_ASAP7_75t_SL g4567 ( 
.A(n_3781),
.B(n_3118),
.C(n_4055),
.Y(n_4567)
);

HB1xp67_ASAP7_75t_L g4568 ( 
.A(n_3997),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4128),
.B(n_4177),
.Y(n_4569)
);

BUFx4f_ASAP7_75t_L g4570 ( 
.A(n_4201),
.Y(n_4570)
);

INVx4_ASAP7_75t_L g4571 ( 
.A(n_3809),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_3737),
.Y(n_4572)
);

NOR2xp33_ASAP7_75t_L g4573 ( 
.A(n_3133),
.B(n_3135),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4177),
.B(n_4228),
.Y(n_4574)
);

BUFx3_ASAP7_75t_L g4575 ( 
.A(n_4053),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_3737),
.Y(n_4576)
);

AND3x1_ASAP7_75t_SL g4577 ( 
.A(n_3781),
.B(n_4085),
.C(n_3810),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_3746),
.Y(n_4578)
);

INVx4_ASAP7_75t_L g4579 ( 
.A(n_3809),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_4040),
.Y(n_4580)
);

BUFx6f_ASAP7_75t_L g4581 ( 
.A(n_4082),
.Y(n_4581)
);

NOR2xp33_ASAP7_75t_L g4582 ( 
.A(n_3155),
.B(n_3163),
.Y(n_4582)
);

BUFx3_ASAP7_75t_L g4583 ( 
.A(n_4082),
.Y(n_4583)
);

INVxp67_ASAP7_75t_L g4584 ( 
.A(n_3746),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4228),
.B(n_4242),
.Y(n_4585)
);

BUFx2_ASAP7_75t_L g4586 ( 
.A(n_4040),
.Y(n_4586)
);

INVx4_ASAP7_75t_L g4587 ( 
.A(n_3809),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_3759),
.Y(n_4588)
);

OAI22xp5_ASAP7_75t_SL g4589 ( 
.A1(n_4473),
.A2(n_3128),
.B1(n_3727),
.B2(n_3122),
.Y(n_4589)
);

INVx1_ASAP7_75t_SL g4590 ( 
.A(n_3710),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4242),
.B(n_4243),
.Y(n_4591)
);

INVx2_ASAP7_75t_SL g4592 ( 
.A(n_4206),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4243),
.B(n_4295),
.Y(n_4593)
);

AOI22xp5_ASAP7_75t_L g4594 ( 
.A1(n_4081),
.A2(n_4139),
.B1(n_4466),
.B2(n_4106),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_3759),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_SL g4596 ( 
.A(n_4295),
.B(n_4323),
.Y(n_4596)
);

A2O1A1Ixp33_ASAP7_75t_L g4597 ( 
.A1(n_3928),
.A2(n_4075),
.B(n_4108),
.C(n_4029),
.Y(n_4597)
);

INVx4_ASAP7_75t_L g4598 ( 
.A(n_3860),
.Y(n_4598)
);

INVx2_ASAP7_75t_SL g4599 ( 
.A(n_4206),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4323),
.B(n_4343),
.Y(n_4600)
);

BUFx2_ASAP7_75t_L g4601 ( 
.A(n_4443),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4343),
.B(n_4388),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4388),
.B(n_4412),
.Y(n_4603)
);

AND2x4_ASAP7_75t_L g4604 ( 
.A(n_4206),
.B(n_4359),
.Y(n_4604)
);

OR2x6_ASAP7_75t_L g4605 ( 
.A(n_3917),
.B(n_4326),
.Y(n_4605)
);

INVx1_ASAP7_75t_SL g4606 ( 
.A(n_3710),
.Y(n_4606)
);

BUFx2_ASAP7_75t_L g4607 ( 
.A(n_4443),
.Y(n_4607)
);

BUFx12f_ASAP7_75t_L g4608 ( 
.A(n_4054),
.Y(n_4608)
);

CKINVDCx5p33_ASAP7_75t_R g4609 ( 
.A(n_3363),
.Y(n_4609)
);

BUFx2_ASAP7_75t_L g4610 ( 
.A(n_3716),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4412),
.B(n_4432),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4432),
.B(n_4433),
.Y(n_4612)
);

INVx1_ASAP7_75t_SL g4613 ( 
.A(n_3563),
.Y(n_4613)
);

BUFx6f_ASAP7_75t_L g4614 ( 
.A(n_4359),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_3760),
.Y(n_4615)
);

OR2x4_ASAP7_75t_L g4616 ( 
.A(n_3722),
.B(n_3824),
.Y(n_4616)
);

INVxp67_ASAP7_75t_L g4617 ( 
.A(n_3760),
.Y(n_4617)
);

BUFx6f_ASAP7_75t_L g4618 ( 
.A(n_4359),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4433),
.B(n_4453),
.Y(n_4619)
);

BUFx6f_ASAP7_75t_L g4620 ( 
.A(n_3917),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_3775),
.Y(n_4621)
);

NOR2x2_ASAP7_75t_L g4622 ( 
.A(n_3339),
.B(n_3179),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_SL g4623 ( 
.A(n_4453),
.B(n_3101),
.Y(n_4623)
);

INVx2_ASAP7_75t_SL g4624 ( 
.A(n_3304),
.Y(n_4624)
);

NOR2xp33_ASAP7_75t_L g4625 ( 
.A(n_4139),
.B(n_4466),
.Y(n_4625)
);

INVx4_ASAP7_75t_L g4626 ( 
.A(n_3860),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_3107),
.B(n_3108),
.Y(n_4627)
);

BUFx4f_ASAP7_75t_L g4628 ( 
.A(n_4201),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_3794),
.Y(n_4629)
);

AOI221xp5_ASAP7_75t_L g4630 ( 
.A1(n_3749),
.A2(n_3754),
.B1(n_3789),
.B2(n_3786),
.C(n_3773),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_3821),
.Y(n_4631)
);

A2O1A1Ixp33_ASAP7_75t_L g4632 ( 
.A1(n_4142),
.A2(n_4165),
.B(n_4235),
.C(n_4151),
.Y(n_4632)
);

OR2x2_ASAP7_75t_L g4633 ( 
.A(n_3188),
.B(n_3755),
.Y(n_4633)
);

AOI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_3812),
.A2(n_3857),
.B1(n_4058),
.B2(n_3838),
.Y(n_4634)
);

NOR2xp33_ASAP7_75t_L g4635 ( 
.A(n_3099),
.B(n_3848),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_SL g4636 ( 
.A(n_3101),
.B(n_3075),
.Y(n_4636)
);

CKINVDCx20_ASAP7_75t_R g4637 ( 
.A(n_3861),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_3821),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_3107),
.B(n_3108),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_3304),
.B(n_3329),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_3363),
.Y(n_4641)
);

BUFx2_ASAP7_75t_L g4642 ( 
.A(n_4008),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_3125),
.B(n_3282),
.Y(n_4643)
);

AND2x4_ASAP7_75t_L g4644 ( 
.A(n_3329),
.B(n_3386),
.Y(n_4644)
);

AND2x4_ASAP7_75t_L g4645 ( 
.A(n_3329),
.B(n_3386),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_3125),
.B(n_3939),
.Y(n_4646)
);

NOR2xp33_ASAP7_75t_L g4647 ( 
.A(n_3099),
.B(n_3848),
.Y(n_4647)
);

HB1xp67_ASAP7_75t_L g4648 ( 
.A(n_3830),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_3939),
.B(n_3106),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_3121),
.B(n_3127),
.Y(n_4650)
);

AOI22xp5_ASAP7_75t_L g4651 ( 
.A1(n_4101),
.A2(n_4155),
.B1(n_4211),
.B2(n_4146),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_3188),
.B(n_3718),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_3742),
.B(n_3743),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_3830),
.Y(n_4654)
);

CKINVDCx16_ASAP7_75t_R g4655 ( 
.A(n_3946),
.Y(n_4655)
);

BUFx4f_ASAP7_75t_L g4656 ( 
.A(n_4201),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_3742),
.B(n_3743),
.Y(n_4657)
);

INVx2_ASAP7_75t_SL g4658 ( 
.A(n_3329),
.Y(n_4658)
);

INVx1_ASAP7_75t_SL g4659 ( 
.A(n_3563),
.Y(n_4659)
);

AND2x6_ASAP7_75t_L g4660 ( 
.A(n_3722),
.B(n_3824),
.Y(n_4660)
);

NAND2x1_ASAP7_75t_L g4661 ( 
.A(n_3713),
.B(n_3800),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_3833),
.Y(n_4662)
);

AND2x4_ASAP7_75t_L g4663 ( 
.A(n_3386),
.B(n_3465),
.Y(n_4663)
);

BUFx6f_ASAP7_75t_L g4664 ( 
.A(n_4074),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_3756),
.B(n_3763),
.Y(n_4665)
);

AND2x6_ASAP7_75t_L g4666 ( 
.A(n_3722),
.B(n_3824),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_3468),
.Y(n_4667)
);

INVx4_ASAP7_75t_L g4668 ( 
.A(n_3860),
.Y(n_4668)
);

NAND2x2_ASAP7_75t_L g4669 ( 
.A(n_4174),
.B(n_3323),
.Y(n_4669)
);

BUFx2_ASAP7_75t_L g4670 ( 
.A(n_3152),
.Y(n_4670)
);

AND2x4_ASAP7_75t_L g4671 ( 
.A(n_3386),
.B(n_3465),
.Y(n_4671)
);

AOI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4249),
.A2(n_4324),
.B1(n_4261),
.B2(n_3749),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_3833),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_3465),
.B(n_3478),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_3841),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_3756),
.B(n_3763),
.Y(n_4676)
);

OAI22xp5_ASAP7_75t_L g4677 ( 
.A1(n_3754),
.A2(n_3786),
.B1(n_3789),
.B2(n_3773),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_3788),
.B(n_3808),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_3841),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_3788),
.B(n_3808),
.Y(n_4680)
);

BUFx2_ASAP7_75t_L g4681 ( 
.A(n_3152),
.Y(n_4681)
);

INVx1_ASAP7_75t_SL g4682 ( 
.A(n_3259),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_3843),
.Y(n_4683)
);

CKINVDCx20_ASAP7_75t_R g4684 ( 
.A(n_3398),
.Y(n_4684)
);

CKINVDCx20_ASAP7_75t_R g4685 ( 
.A(n_3240),
.Y(n_4685)
);

INVxp67_ASAP7_75t_SL g4686 ( 
.A(n_3755),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_3843),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_3823),
.B(n_3966),
.Y(n_4688)
);

BUFx2_ASAP7_75t_L g4689 ( 
.A(n_3082),
.Y(n_4689)
);

NOR2xp33_ASAP7_75t_L g4690 ( 
.A(n_3946),
.B(n_3161),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_3823),
.B(n_3966),
.Y(n_4691)
);

NOR2xp33_ASAP7_75t_R g4692 ( 
.A(n_3431),
.B(n_3950),
.Y(n_4692)
);

HB1xp67_ASAP7_75t_L g4693 ( 
.A(n_3845),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4017),
.B(n_4048),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4017),
.B(n_4048),
.Y(n_4695)
);

NOR2xp33_ASAP7_75t_L g4696 ( 
.A(n_3826),
.B(n_3832),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_3845),
.Y(n_4697)
);

OR2x6_ASAP7_75t_L g4698 ( 
.A(n_4326),
.B(n_3395),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_3849),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4067),
.B(n_4080),
.Y(n_4700)
);

NOR2x1_ASAP7_75t_L g4701 ( 
.A(n_3157),
.B(n_3095),
.Y(n_4701)
);

AOI22xp5_ASAP7_75t_L g4702 ( 
.A1(n_3826),
.A2(n_3832),
.B1(n_3869),
.B2(n_3859),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4067),
.B(n_4080),
.Y(n_4703)
);

BUFx6f_ASAP7_75t_L g4704 ( 
.A(n_4326),
.Y(n_4704)
);

BUFx6f_ASAP7_75t_L g4705 ( 
.A(n_4326),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_3849),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_3850),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4111),
.B(n_4115),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_3850),
.Y(n_4709)
);

CKINVDCx5p33_ASAP7_75t_R g4710 ( 
.A(n_3468),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_3082),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_3852),
.Y(n_4712)
);

BUFx8_ASAP7_75t_L g4713 ( 
.A(n_3722),
.Y(n_4713)
);

INVx1_ASAP7_75t_SL g4714 ( 
.A(n_3259),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4111),
.B(n_4115),
.Y(n_4715)
);

AOI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_3859),
.A2(n_3869),
.B1(n_3927),
.B2(n_3904),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_3075),
.B(n_3115),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4137),
.B(n_4157),
.Y(n_4718)
);

AOI21xp5_ASAP7_75t_L g4719 ( 
.A1(n_3732),
.A2(n_3739),
.B(n_3735),
.Y(n_4719)
);

INVx2_ASAP7_75t_SL g4720 ( 
.A(n_3493),
.Y(n_4720)
);

AOI22x1_ASAP7_75t_L g4721 ( 
.A1(n_3192),
.A2(n_3198),
.B1(n_3190),
.B2(n_3197),
.Y(n_4721)
);

BUFx3_ASAP7_75t_L g4722 ( 
.A(n_3493),
.Y(n_4722)
);

AOI22xp33_ASAP7_75t_L g4723 ( 
.A1(n_3962),
.A2(n_4083),
.B1(n_4365),
.B2(n_4072),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_L g4724 ( 
.A(n_4137),
.B(n_4157),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4185),
.B(n_4192),
.Y(n_4725)
);

OAI22xp5_ASAP7_75t_L g4726 ( 
.A1(n_3904),
.A2(n_3944),
.B1(n_3994),
.B2(n_3927),
.Y(n_4726)
);

BUFx6f_ASAP7_75t_L g4727 ( 
.A(n_3171),
.Y(n_4727)
);

NAND2x1p5_ASAP7_75t_L g4728 ( 
.A(n_3713),
.B(n_3800),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_3852),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4185),
.B(n_4192),
.Y(n_4730)
);

CKINVDCx5p33_ASAP7_75t_R g4731 ( 
.A(n_3941),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4213),
.B(n_4284),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4213),
.B(n_4284),
.Y(n_4733)
);

BUFx3_ASAP7_75t_L g4734 ( 
.A(n_3179),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4290),
.B(n_4294),
.Y(n_4735)
);

CKINVDCx5p33_ASAP7_75t_R g4736 ( 
.A(n_3941),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_3853),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4290),
.B(n_4294),
.Y(n_4738)
);

BUFx2_ASAP7_75t_L g4739 ( 
.A(n_3112),
.Y(n_4739)
);

AOI22xp5_ASAP7_75t_L g4740 ( 
.A1(n_3944),
.A2(n_3994),
.B1(n_4019),
.B2(n_4005),
.Y(n_4740)
);

BUFx6f_ASAP7_75t_L g4741 ( 
.A(n_3171),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_3853),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_3867),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_3867),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4311),
.B(n_4329),
.Y(n_4745)
);

OAI22xp5_ASAP7_75t_L g4746 ( 
.A1(n_4005),
.A2(n_4037),
.B1(n_4087),
.B2(n_4019),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4311),
.B(n_4329),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4396),
.B(n_4397),
.Y(n_4748)
);

O2A1O1Ixp33_ASAP7_75t_L g4749 ( 
.A1(n_3719),
.A2(n_3816),
.B(n_3972),
.C(n_3942),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4396),
.B(n_4397),
.Y(n_4750)
);

CKINVDCx14_ASAP7_75t_R g4751 ( 
.A(n_3458),
.Y(n_4751)
);

OR2x6_ASAP7_75t_L g4752 ( 
.A(n_3395),
.B(n_4298),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_3878),
.Y(n_4753)
);

BUFx3_ASAP7_75t_L g4754 ( 
.A(n_3179),
.Y(n_4754)
);

AOI22xp33_ASAP7_75t_L g4755 ( 
.A1(n_3146),
.A2(n_4231),
.B1(n_3983),
.B2(n_3174),
.Y(n_4755)
);

NOR2xp33_ASAP7_75t_R g4756 ( 
.A(n_3431),
.B(n_3950),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4447),
.B(n_3184),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4298),
.B(n_3114),
.Y(n_4758)
);

CKINVDCx20_ASAP7_75t_R g4759 ( 
.A(n_3232),
.Y(n_4759)
);

OR2x6_ASAP7_75t_L g4760 ( 
.A(n_3179),
.B(n_3744),
.Y(n_4760)
);

A2O1A1Ixp33_ASAP7_75t_L g4761 ( 
.A1(n_4304),
.A2(n_4427),
.B(n_4021),
.C(n_4030),
.Y(n_4761)
);

CKINVDCx5p33_ASAP7_75t_R g4762 ( 
.A(n_4198),
.Y(n_4762)
);

INVx2_ASAP7_75t_SL g4763 ( 
.A(n_3934),
.Y(n_4763)
);

A2O1A1Ixp33_ASAP7_75t_L g4764 ( 
.A1(n_3993),
.A2(n_4060),
.B(n_4131),
.C(n_4046),
.Y(n_4764)
);

BUFx3_ASAP7_75t_L g4765 ( 
.A(n_3179),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4447),
.B(n_3277),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_3280),
.B(n_3283),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_3285),
.B(n_3289),
.Y(n_4768)
);

BUFx2_ASAP7_75t_L g4769 ( 
.A(n_3114),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_3878),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_3301),
.B(n_3302),
.Y(n_4771)
);

BUFx6f_ASAP7_75t_L g4772 ( 
.A(n_3950),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_3882),
.Y(n_4773)
);

BUFx2_ASAP7_75t_L g4774 ( 
.A(n_3730),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_SL g4775 ( 
.A(n_3115),
.B(n_3740),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_3882),
.Y(n_4776)
);

OAI22xp5_ASAP7_75t_L g4777 ( 
.A1(n_4037),
.A2(n_4217),
.B1(n_4301),
.B2(n_4087),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_3143),
.B(n_3148),
.Y(n_4778)
);

BUFx8_ASAP7_75t_L g4779 ( 
.A(n_3824),
.Y(n_4779)
);

CKINVDCx20_ASAP7_75t_R g4780 ( 
.A(n_3169),
.Y(n_4780)
);

NOR2xp33_ASAP7_75t_L g4781 ( 
.A(n_4217),
.B(n_4301),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_3883),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_3883),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_3143),
.B(n_3148),
.Y(n_4784)
);

INVxp67_ASAP7_75t_L g4785 ( 
.A(n_3888),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_3888),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_3740),
.B(n_3741),
.Y(n_4787)
);

INVx2_ASAP7_75t_SL g4788 ( 
.A(n_3934),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_SL g4789 ( 
.A(n_3741),
.B(n_3933),
.Y(n_4789)
);

INVx2_ASAP7_75t_SL g4790 ( 
.A(n_3961),
.Y(n_4790)
);

BUFx2_ASAP7_75t_L g4791 ( 
.A(n_3797),
.Y(n_4791)
);

OR2x6_ASAP7_75t_L g4792 ( 
.A(n_4476),
.B(n_3796),
.Y(n_4792)
);

INVx6_ASAP7_75t_L g4793 ( 
.A(n_3862),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_3889),
.Y(n_4794)
);

AOI22xp33_ASAP7_75t_L g4795 ( 
.A1(n_4345),
.A2(n_4473),
.B1(n_4391),
.B2(n_3177),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_3889),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4345),
.B(n_4391),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_3907),
.Y(n_4798)
);

OR2x4_ASAP7_75t_L g4799 ( 
.A(n_4038),
.B(n_4043),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_3907),
.Y(n_4800)
);

NOR2xp33_ASAP7_75t_L g4801 ( 
.A(n_3084),
.B(n_3105),
.Y(n_4801)
);

INVxp67_ASAP7_75t_L g4802 ( 
.A(n_3911),
.Y(n_4802)
);

AND3x2_ASAP7_75t_SL g4803 ( 
.A(n_3308),
.B(n_3284),
.C(n_3418),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_3911),
.Y(n_4804)
);

BUFx2_ASAP7_75t_L g4805 ( 
.A(n_3856),
.Y(n_4805)
);

CKINVDCx20_ASAP7_75t_R g4806 ( 
.A(n_3169),
.Y(n_4806)
);

AND2x6_ASAP7_75t_L g4807 ( 
.A(n_4038),
.B(n_4043),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_3916),
.Y(n_4808)
);

AO21x2_ASAP7_75t_L g4809 ( 
.A1(n_3308),
.A2(n_3440),
.B(n_3839),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_R g4810 ( 
.A(n_3950),
.B(n_4097),
.Y(n_4810)
);

BUFx2_ASAP7_75t_L g4811 ( 
.A(n_3858),
.Y(n_4811)
);

AO22x1_ASAP7_75t_L g4812 ( 
.A1(n_3103),
.A2(n_3186),
.B1(n_3208),
.B2(n_3205),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_3933),
.B(n_3979),
.Y(n_4813)
);

BUFx6f_ASAP7_75t_L g4814 ( 
.A(n_4097),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_3916),
.Y(n_4815)
);

BUFx2_ASAP7_75t_L g4816 ( 
.A(n_3858),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_3979),
.B(n_4059),
.Y(n_4817)
);

INVx2_ASAP7_75t_SL g4818 ( 
.A(n_3961),
.Y(n_4818)
);

AO22x1_ASAP7_75t_L g4819 ( 
.A1(n_3103),
.A2(n_3186),
.B1(n_3208),
.B2(n_3205),
.Y(n_4819)
);

AOI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_3723),
.A2(n_3902),
.B1(n_4103),
.B2(n_3750),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_SL g4821 ( 
.A(n_4059),
.B(n_4218),
.Y(n_4821)
);

BUFx2_ASAP7_75t_L g4822 ( 
.A(n_3863),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_3929),
.Y(n_4823)
);

BUFx2_ASAP7_75t_L g4824 ( 
.A(n_3871),
.Y(n_4824)
);

NOR2xp67_ASAP7_75t_L g4825 ( 
.A(n_3132),
.B(n_3158),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_3929),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4218),
.B(n_4253),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_3752),
.A2(n_3780),
.B1(n_3828),
.B2(n_3758),
.Y(n_4828)
);

BUFx2_ASAP7_75t_L g4829 ( 
.A(n_3871),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4253),
.B(n_4259),
.Y(n_4830)
);

BUFx2_ASAP7_75t_L g4831 ( 
.A(n_3901),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4259),
.B(n_4264),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4264),
.B(n_4346),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_3935),
.Y(n_4834)
);

INVxp67_ASAP7_75t_L g4835 ( 
.A(n_3935),
.Y(n_4835)
);

INVxp67_ASAP7_75t_SL g4836 ( 
.A(n_4001),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4346),
.B(n_4353),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_3938),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_3938),
.Y(n_4839)
);

INVx2_ASAP7_75t_SL g4840 ( 
.A(n_4001),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4353),
.B(n_4469),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_3948),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_3855),
.B(n_3895),
.Y(n_4843)
);

BUFx2_ASAP7_75t_L g4844 ( 
.A(n_3901),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_3897),
.B(n_3906),
.Y(n_4845)
);

CKINVDCx5p33_ASAP7_75t_R g4846 ( 
.A(n_4198),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_3913),
.B(n_3915),
.Y(n_4847)
);

BUFx2_ASAP7_75t_L g4848 ( 
.A(n_3901),
.Y(n_4848)
);

INVx4_ASAP7_75t_L g4849 ( 
.A(n_4097),
.Y(n_4849)
);

INVx2_ASAP7_75t_SL g4850 ( 
.A(n_3948),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_3940),
.B(n_3968),
.Y(n_4851)
);

NOR2xp67_ASAP7_75t_L g4852 ( 
.A(n_3751),
.B(n_3761),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_3992),
.B(n_3996),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_3949),
.Y(n_4854)
);

AOI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_3764),
.A2(n_3771),
.B(n_3766),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4000),
.B(n_4025),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_3949),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4069),
.B(n_4117),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_SL g4859 ( 
.A(n_4097),
.B(n_4104),
.Y(n_4859)
);

INVx4_ASAP7_75t_L g4860 ( 
.A(n_4104),
.Y(n_4860)
);

BUFx2_ASAP7_75t_L g4861 ( 
.A(n_3920),
.Y(n_4861)
);

AOI21x1_ASAP7_75t_L g4862 ( 
.A1(n_3779),
.A2(n_3811),
.B(n_3804),
.Y(n_4862)
);

BUFx8_ASAP7_75t_L g4863 ( 
.A(n_4043),
.Y(n_4863)
);

NOR2xp67_ASAP7_75t_L g4864 ( 
.A(n_3813),
.B(n_3815),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4138),
.B(n_4166),
.Y(n_4865)
);

CKINVDCx5p33_ASAP7_75t_R g4866 ( 
.A(n_4314),
.Y(n_4866)
);

NOR2xp33_ASAP7_75t_L g4867 ( 
.A(n_4172),
.B(n_4183),
.Y(n_4867)
);

INVx4_ASAP7_75t_L g4868 ( 
.A(n_4104),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_3952),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_3921),
.B(n_3955),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_3952),
.Y(n_4871)
);

INVxp67_ASAP7_75t_SL g4872 ( 
.A(n_3954),
.Y(n_4872)
);

HB1xp67_ASAP7_75t_L g4873 ( 
.A(n_3954),
.Y(n_4873)
);

HB1xp67_ASAP7_75t_L g4874 ( 
.A(n_3959),
.Y(n_4874)
);

INVx5_ASAP7_75t_L g4875 ( 
.A(n_4098),
.Y(n_4875)
);

BUFx2_ASAP7_75t_L g4876 ( 
.A(n_3955),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_3959),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_3971),
.Y(n_4878)
);

BUFx2_ASAP7_75t_L g4879 ( 
.A(n_3976),
.Y(n_4879)
);

CKINVDCx5p33_ASAP7_75t_R g4880 ( 
.A(n_4314),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_3971),
.Y(n_4881)
);

INVx3_ASAP7_75t_SL g4882 ( 
.A(n_3087),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4194),
.B(n_4223),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4257),
.B(n_4262),
.Y(n_4884)
);

AND3x1_ASAP7_75t_SL g4885 ( 
.A(n_4136),
.B(n_4159),
.C(n_4147),
.Y(n_4885)
);

NAND2x1p5_ASAP7_75t_L g4886 ( 
.A(n_3919),
.B(n_3931),
.Y(n_4886)
);

HB1xp67_ASAP7_75t_L g4887 ( 
.A(n_3977),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4269),
.B(n_4320),
.Y(n_4888)
);

HB1xp67_ASAP7_75t_L g4889 ( 
.A(n_3977),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_3982),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_SL g4891 ( 
.A(n_4104),
.B(n_4178),
.Y(n_4891)
);

HB1xp67_ASAP7_75t_L g4892 ( 
.A(n_3982),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4337),
.B(n_4459),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_3985),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4364),
.B(n_4409),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4411),
.B(n_4444),
.Y(n_4896)
);

OR2x2_ASAP7_75t_L g4897 ( 
.A(n_4465),
.B(n_3985),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_3986),
.Y(n_4898)
);

INVx4_ASAP7_75t_L g4899 ( 
.A(n_4178),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_3986),
.Y(n_4900)
);

INVx4_ASAP7_75t_L g4901 ( 
.A(n_4178),
.Y(n_4901)
);

AND3x1_ASAP7_75t_SL g4902 ( 
.A(n_4167),
.B(n_4224),
.C(n_4210),
.Y(n_4902)
);

NOR2xp33_ASAP7_75t_L g4903 ( 
.A(n_3274),
.B(n_4265),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_3988),
.Y(n_4904)
);

BUFx2_ASAP7_75t_L g4905 ( 
.A(n_4018),
.Y(n_4905)
);

CKINVDCx5p33_ASAP7_75t_R g4906 ( 
.A(n_4086),
.Y(n_4906)
);

INVxp67_ASAP7_75t_L g4907 ( 
.A(n_3988),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_3274),
.B(n_3217),
.Y(n_4908)
);

OR2x2_ASAP7_75t_L g4909 ( 
.A(n_3990),
.B(n_4458),
.Y(n_4909)
);

BUFx4f_ASAP7_75t_SL g4910 ( 
.A(n_3467),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_3990),
.Y(n_4911)
);

INVx2_ASAP7_75t_SL g4912 ( 
.A(n_3991),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_3219),
.B(n_3225),
.Y(n_4913)
);

AOI221xp5_ASAP7_75t_L g4914 ( 
.A1(n_3187),
.A2(n_3175),
.B1(n_3141),
.B2(n_3200),
.C(n_3197),
.Y(n_4914)
);

BUFx4f_ASAP7_75t_L g4915 ( 
.A(n_4201),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_SL g4916 ( 
.A(n_4178),
.B(n_4374),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_3991),
.Y(n_4917)
);

INVx6_ASAP7_75t_L g4918 ( 
.A(n_3862),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_3226),
.B(n_3234),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_3245),
.B(n_3247),
.Y(n_4920)
);

AOI22xp5_ASAP7_75t_L g4921 ( 
.A1(n_3320),
.A2(n_3391),
.B1(n_3111),
.B2(n_3078),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_3248),
.B(n_3249),
.Y(n_4922)
);

BUFx2_ASAP7_75t_L g4923 ( 
.A(n_4018),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_3995),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_3995),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_3252),
.B(n_3256),
.Y(n_4926)
);

BUFx2_ASAP7_75t_L g4927 ( 
.A(n_4039),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_3257),
.B(n_3263),
.Y(n_4928)
);

OR2x6_ASAP7_75t_L g4929 ( 
.A(n_4468),
.B(n_4470),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4374),
.B(n_4457),
.Y(n_4930)
);

INVxp67_ASAP7_75t_L g4931 ( 
.A(n_3998),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_3998),
.Y(n_4932)
);

NOR2xp33_ASAP7_75t_L g4933 ( 
.A(n_4319),
.B(n_4356),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4002),
.Y(n_4934)
);

BUFx2_ASAP7_75t_L g4935 ( 
.A(n_4039),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4039),
.B(n_4079),
.Y(n_4936)
);

AOI22xp33_ASAP7_75t_L g4937 ( 
.A1(n_3203),
.A2(n_3085),
.B1(n_3753),
.B2(n_3747),
.Y(n_4937)
);

BUFx4f_ASAP7_75t_L g4938 ( 
.A(n_4201),
.Y(n_4938)
);

OR2x6_ASAP7_75t_L g4939 ( 
.A(n_4471),
.B(n_3831),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4002),
.Y(n_4940)
);

AOI22xp5_ASAP7_75t_L g4941 ( 
.A1(n_3320),
.A2(n_3774),
.B1(n_3791),
.B2(n_3772),
.Y(n_4941)
);

AOI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_3802),
.A2(n_3827),
.B1(n_3879),
.B2(n_3807),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_L g4943 ( 
.A(n_4357),
.B(n_4358),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_3264),
.B(n_3267),
.Y(n_4944)
);

AND2x6_ASAP7_75t_L g4945 ( 
.A(n_4119),
.B(n_4199),
.Y(n_4945)
);

AND3x1_ASAP7_75t_SL g4946 ( 
.A(n_4384),
.B(n_4417),
.C(n_4401),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_3269),
.B(n_3442),
.Y(n_4947)
);

OAI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4462),
.A2(n_4204),
.B1(n_3185),
.B2(n_3193),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_3444),
.B(n_3448),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4014),
.Y(n_4950)
);

HB1xp67_ASAP7_75t_L g4951 ( 
.A(n_4014),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_3449),
.B(n_3278),
.Y(n_4952)
);

HB1xp67_ASAP7_75t_L g4953 ( 
.A(n_4023),
.Y(n_4953)
);

AND2x6_ASAP7_75t_L g4954 ( 
.A(n_4199),
.B(n_4303),
.Y(n_4954)
);

INVx2_ASAP7_75t_SL g4955 ( 
.A(n_4023),
.Y(n_4955)
);

BUFx2_ASAP7_75t_L g4956 ( 
.A(n_4092),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_3278),
.B(n_3157),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4033),
.Y(n_4958)
);

AOI22x1_ASAP7_75t_L g4959 ( 
.A1(n_3200),
.A2(n_3191),
.B1(n_3819),
.B2(n_3818),
.Y(n_4959)
);

BUFx2_ASAP7_75t_L g4960 ( 
.A(n_4092),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4033),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4045),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_3825),
.A2(n_3834),
.B(n_3829),
.Y(n_4963)
);

INVx4_ASAP7_75t_L g4964 ( 
.A(n_4374),
.Y(n_4964)
);

INVx4_ASAP7_75t_L g4965 ( 
.A(n_4374),
.Y(n_4965)
);

O2A1O1Ixp5_ASAP7_75t_L g4966 ( 
.A1(n_3885),
.A2(n_3922),
.B(n_3924),
.C(n_3892),
.Y(n_4966)
);

AOI22xp33_ASAP7_75t_L g4967 ( 
.A1(n_3203),
.A2(n_3953),
.B1(n_4004),
.B2(n_3969),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_SL g4968 ( 
.A(n_4457),
.B(n_3142),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4045),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4050),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4050),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4061),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_SL g4973 ( 
.A(n_4457),
.B(n_3142),
.Y(n_4973)
);

INVx1_ASAP7_75t_SL g4974 ( 
.A(n_3459),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4061),
.Y(n_4975)
);

NOR2xp67_ASAP7_75t_L g4976 ( 
.A(n_3835),
.B(n_3840),
.Y(n_4976)
);

NOR2xp33_ASAP7_75t_L g4977 ( 
.A(n_3268),
.B(n_3880),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_4086),
.Y(n_4978)
);

HB1xp67_ASAP7_75t_L g4979 ( 
.A(n_4070),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_3392),
.B(n_3353),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_3392),
.B(n_4070),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4073),
.Y(n_4982)
);

INVx1_ASAP7_75t_SL g4983 ( 
.A(n_3459),
.Y(n_4983)
);

INVxp67_ASAP7_75t_L g4984 ( 
.A(n_4073),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4076),
.B(n_4077),
.Y(n_4985)
);

AOI22xp33_ASAP7_75t_L g4986 ( 
.A1(n_4007),
.A2(n_4034),
.B1(n_4049),
.B2(n_4035),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4076),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4077),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4088),
.Y(n_4989)
);

AOI21xp5_ASAP7_75t_L g4990 ( 
.A1(n_3842),
.A2(n_3868),
.B(n_3854),
.Y(n_4990)
);

HB1xp67_ASAP7_75t_L g4991 ( 
.A(n_4088),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4094),
.B(n_4099),
.Y(n_4992)
);

NOR2xp33_ASAP7_75t_L g4993 ( 
.A(n_3268),
.B(n_3880),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4094),
.Y(n_4994)
);

AND2x4_ASAP7_75t_L g4995 ( 
.A(n_4170),
.B(n_4181),
.Y(n_4995)
);

HB1xp67_ASAP7_75t_L g4996 ( 
.A(n_4099),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4102),
.B(n_4105),
.Y(n_4997)
);

AND2x4_ASAP7_75t_L g4998 ( 
.A(n_4181),
.B(n_4191),
.Y(n_4998)
);

NAND3xp33_ASAP7_75t_L g4999 ( 
.A(n_3999),
.B(n_4328),
.C(n_3173),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_SL g5000 ( 
.A(n_4457),
.B(n_3138),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4102),
.B(n_4105),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4118),
.Y(n_5002)
);

INVx4_ASAP7_75t_L g5003 ( 
.A(n_3862),
.Y(n_5003)
);

OR2x2_ASAP7_75t_L g5004 ( 
.A(n_4118),
.B(n_4121),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4121),
.Y(n_5005)
);

NAND2x1p5_ASAP7_75t_L g5006 ( 
.A(n_3919),
.B(n_3931),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4122),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4122),
.Y(n_5008)
);

OR2x6_ASAP7_75t_L g5009 ( 
.A(n_4011),
.B(n_4031),
.Y(n_5009)
);

AOI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4051),
.A2(n_4133),
.B1(n_4134),
.B2(n_4093),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4125),
.Y(n_5011)
);

HB1xp67_ASAP7_75t_L g5012 ( 
.A(n_4125),
.Y(n_5012)
);

INVx2_ASAP7_75t_SL g5013 ( 
.A(n_4135),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4135),
.B(n_4141),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4141),
.B(n_4144),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4144),
.B(n_4145),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_SL g5017 ( 
.A(n_3087),
.B(n_3975),
.Y(n_5017)
);

INVxp67_ASAP7_75t_SL g5018 ( 
.A(n_4145),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4153),
.Y(n_5019)
);

OR2x2_ASAP7_75t_L g5020 ( 
.A(n_4153),
.B(n_4164),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4164),
.Y(n_5021)
);

INVxp67_ASAP7_75t_SL g5022 ( 
.A(n_4168),
.Y(n_5022)
);

INVx2_ASAP7_75t_SL g5023 ( 
.A(n_4168),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4203),
.B(n_4209),
.Y(n_5024)
);

NAND2xp33_ASAP7_75t_SL g5025 ( 
.A(n_3094),
.B(n_3098),
.Y(n_5025)
);

INVxp67_ASAP7_75t_SL g5026 ( 
.A(n_4176),
.Y(n_5026)
);

HB1xp67_ASAP7_75t_L g5027 ( 
.A(n_4176),
.Y(n_5027)
);

CKINVDCx8_ASAP7_75t_R g5028 ( 
.A(n_4303),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4184),
.B(n_4188),
.Y(n_5029)
);

HB1xp67_ASAP7_75t_L g5030 ( 
.A(n_4184),
.Y(n_5030)
);

INVx4_ASAP7_75t_L g5031 ( 
.A(n_3862),
.Y(n_5031)
);

CKINVDCx5p33_ASAP7_75t_R g5032 ( 
.A(n_4143),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4188),
.B(n_4190),
.Y(n_5033)
);

OR2x6_ASAP7_75t_L g5034 ( 
.A(n_3874),
.B(n_3875),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4190),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_4197),
.B(n_4208),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4197),
.B(n_4208),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4214),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4214),
.Y(n_5039)
);

NOR2xp67_ASAP7_75t_L g5040 ( 
.A(n_3877),
.B(n_3891),
.Y(n_5040)
);

HB1xp67_ASAP7_75t_L g5041 ( 
.A(n_4222),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4222),
.Y(n_5042)
);

INVx3_ASAP7_75t_SL g5043 ( 
.A(n_3087),
.Y(n_5043)
);

NOR2x1_ASAP7_75t_L g5044 ( 
.A(n_3156),
.B(n_4465),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4238),
.Y(n_5045)
);

OAI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4161),
.A2(n_4216),
.B(n_4207),
.Y(n_5046)
);

AOI22xp33_ASAP7_75t_L g5047 ( 
.A1(n_4258),
.A2(n_4270),
.B1(n_4273),
.B2(n_4271),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4238),
.B(n_4239),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4239),
.B(n_4241),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4241),
.Y(n_5050)
);

INVx5_ASAP7_75t_L g5051 ( 
.A(n_4370),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4266),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4266),
.B(n_4268),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4268),
.B(n_4274),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4274),
.B(n_4281),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4281),
.Y(n_5056)
);

OAI221xp5_ASAP7_75t_L g5057 ( 
.A1(n_3187),
.A2(n_3189),
.B1(n_3109),
.B2(n_3162),
.C(n_3139),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4287),
.B(n_4291),
.Y(n_5058)
);

NOR2xp33_ASAP7_75t_L g5059 ( 
.A(n_3136),
.B(n_3185),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4287),
.Y(n_5060)
);

AND2x2_ASAP7_75t_SL g5061 ( 
.A(n_3975),
.B(n_4120),
.Y(n_5061)
);

INVx2_ASAP7_75t_SL g5062 ( 
.A(n_4291),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4300),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4300),
.B(n_4313),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4313),
.B(n_4317),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_SL g5066 ( 
.A(n_3975),
.B(n_4120),
.Y(n_5066)
);

INVx4_ASAP7_75t_L g5067 ( 
.A(n_4013),
.Y(n_5067)
);

INVx2_ASAP7_75t_SL g5068 ( 
.A(n_4317),
.Y(n_5068)
);

AOI22xp33_ASAP7_75t_L g5069 ( 
.A1(n_4282),
.A2(n_4285),
.B1(n_4293),
.B2(n_4292),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4321),
.B(n_4331),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_SL g5071 ( 
.A(n_4120),
.B(n_3116),
.Y(n_5071)
);

HB1xp67_ASAP7_75t_L g5072 ( 
.A(n_4321),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4331),
.Y(n_5073)
);

INVxp67_ASAP7_75t_L g5074 ( 
.A(n_4339),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4339),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_4342),
.B(n_4344),
.Y(n_5076)
);

CKINVDCx20_ASAP7_75t_R g5077 ( 
.A(n_4047),
.Y(n_5077)
);

HB1xp67_ASAP7_75t_L g5078 ( 
.A(n_4342),
.Y(n_5078)
);

BUFx2_ASAP7_75t_R g5079 ( 
.A(n_3255),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_SL g5080 ( 
.A(n_3116),
.B(n_3134),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4344),
.Y(n_5081)
);

BUFx2_ASAP7_75t_L g5082 ( 
.A(n_4237),
.Y(n_5082)
);

AND3x1_ASAP7_75t_SL g5083 ( 
.A(n_4174),
.B(n_3782),
.C(n_4204),
.Y(n_5083)
);

NAND3xp33_ASAP7_75t_SL g5084 ( 
.A(n_3715),
.B(n_3896),
.C(n_3864),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_4362),
.B(n_4381),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4362),
.B(n_4381),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4382),
.Y(n_5087)
);

BUFx2_ASAP7_75t_L g5088 ( 
.A(n_4237),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4382),
.B(n_4385),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_3893),
.A2(n_3898),
.B(n_3894),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_SL g5091 ( 
.A(n_3134),
.B(n_4010),
.Y(n_5091)
);

INVxp67_ASAP7_75t_L g5092 ( 
.A(n_4385),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4386),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4386),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4387),
.B(n_4392),
.Y(n_5095)
);

NAND2xp5_ASAP7_75t_SL g5096 ( 
.A(n_4010),
.B(n_4305),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4387),
.Y(n_5097)
);

O2A1O1Ixp33_ASAP7_75t_L g5098 ( 
.A1(n_4299),
.A2(n_4340),
.B(n_4349),
.C(n_4315),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4392),
.Y(n_5099)
);

INVxp67_ASAP7_75t_L g5100 ( 
.A(n_4402),
.Y(n_5100)
);

OR2x2_ASAP7_75t_L g5101 ( 
.A(n_4402),
.B(n_4404),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_L g5102 ( 
.A(n_4404),
.B(n_4406),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4406),
.B(n_4410),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4410),
.B(n_4415),
.Y(n_5104)
);

AOI22xp5_ASAP7_75t_L g5105 ( 
.A1(n_4398),
.A2(n_4418),
.B1(n_4430),
.B2(n_4407),
.Y(n_5105)
);

AOI22xp33_ASAP7_75t_L g5106 ( 
.A1(n_4451),
.A2(n_4463),
.B1(n_3077),
.B2(n_3214),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_4415),
.B(n_4419),
.Y(n_5107)
);

AND2x4_ASAP7_75t_SL g5108 ( 
.A(n_4013),
.B(n_4169),
.Y(n_5108)
);

INVx4_ASAP7_75t_L g5109 ( 
.A(n_4013),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4419),
.Y(n_5110)
);

BUFx2_ASAP7_75t_L g5111 ( 
.A(n_4250),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_4424),
.B(n_4426),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4424),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_4426),
.B(n_4439),
.Y(n_5114)
);

NOR2xp33_ASAP7_75t_L g5115 ( 
.A(n_3136),
.B(n_3193),
.Y(n_5115)
);

AOI22xp33_ASAP7_75t_L g5116 ( 
.A1(n_3212),
.A2(n_3214),
.B1(n_3224),
.B2(n_3222),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_SL g5117 ( 
.A(n_4305),
.B(n_3947),
.Y(n_5117)
);

CKINVDCx20_ASAP7_75t_R g5118 ( 
.A(n_4047),
.Y(n_5118)
);

NOR2xp33_ASAP7_75t_L g5119 ( 
.A(n_3261),
.B(n_3793),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_3261),
.B(n_3793),
.Y(n_5120)
);

O2A1O1Ixp33_ASAP7_75t_L g5121 ( 
.A1(n_3209),
.A2(n_3218),
.B(n_3228),
.C(n_4003),
.Y(n_5121)
);

NOR2xp33_ASAP7_75t_L g5122 ( 
.A(n_3847),
.B(n_4113),
.Y(n_5122)
);

NAND2xp5_ASAP7_75t_L g5123 ( 
.A(n_4439),
.B(n_4449),
.Y(n_5123)
);

INVx5_ASAP7_75t_L g5124 ( 
.A(n_4428),
.Y(n_5124)
);

INVx1_ASAP7_75t_SL g5125 ( 
.A(n_3720),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_4449),
.B(n_4455),
.Y(n_5126)
);

NOR2xp33_ASAP7_75t_L g5127 ( 
.A(n_3847),
.B(n_4113),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_4455),
.B(n_4458),
.Y(n_5128)
);

OAI22xp5_ASAP7_75t_SL g5129 ( 
.A1(n_4179),
.A2(n_4352),
.B1(n_4279),
.B2(n_3297),
.Y(n_5129)
);

BUFx2_ASAP7_75t_L g5130 ( 
.A(n_4250),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_3899),
.A2(n_3912),
.B(n_3903),
.Y(n_5131)
);

AOI22xp33_ASAP7_75t_L g5132 ( 
.A1(n_3212),
.A2(n_3222),
.B1(n_3230),
.B2(n_3224),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_3166),
.B(n_4244),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_3166),
.B(n_4245),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_3487),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_SL g5136 ( 
.A(n_4332),
.B(n_3270),
.Y(n_5136)
);

NOR2xp33_ASAP7_75t_L g5137 ( 
.A(n_4179),
.B(n_4279),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_4254),
.B(n_4260),
.Y(n_5138)
);

BUFx2_ASAP7_75t_L g5139 ( 
.A(n_4252),
.Y(n_5139)
);

OR2x2_ASAP7_75t_L g5140 ( 
.A(n_4260),
.B(n_4267),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_3487),
.Y(n_5141)
);

INVxp67_ASAP7_75t_L g5142 ( 
.A(n_4267),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_4272),
.B(n_4276),
.Y(n_5143)
);

AOI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_3180),
.A2(n_3243),
.B1(n_3265),
.B2(n_3236),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_4276),
.B(n_4277),
.Y(n_5145)
);

HB1xp67_ASAP7_75t_L g5146 ( 
.A(n_3984),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_SL g5147 ( 
.A(n_3270),
.B(n_3144),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_4277),
.B(n_4309),
.Y(n_5148)
);

NOR4xp25_ASAP7_75t_SL g5149 ( 
.A(n_3423),
.B(n_3284),
.C(n_3873),
.D(n_3839),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_3517),
.Y(n_5150)
);

NAND2xp33_ASAP7_75t_L g5151 ( 
.A(n_4126),
.B(n_4352),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_4336),
.B(n_4351),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_3517),
.Y(n_5153)
);

INVx2_ASAP7_75t_SL g5154 ( 
.A(n_4351),
.Y(n_5154)
);

A2O1A1Ixp33_ASAP7_75t_L g5155 ( 
.A1(n_3873),
.A2(n_4193),
.B(n_4233),
.C(n_4090),
.Y(n_5155)
);

NAND3xp33_ASAP7_75t_L g5156 ( 
.A(n_3109),
.B(n_3139),
.C(n_3129),
.Y(n_5156)
);

AO22x1_ASAP7_75t_L g5157 ( 
.A1(n_3230),
.A2(n_3254),
.B1(n_3262),
.B2(n_3260),
.Y(n_5157)
);

INVxp67_ASAP7_75t_SL g5158 ( 
.A(n_4354),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4379),
.B(n_4389),
.Y(n_5159)
);

HB1xp67_ASAP7_75t_L g5160 ( 
.A(n_3984),
.Y(n_5160)
);

INVx2_ASAP7_75t_SL g5161 ( 
.A(n_4403),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4403),
.Y(n_5162)
);

NOR2xp33_ASAP7_75t_L g5163 ( 
.A(n_3782),
.B(n_4464),
.Y(n_5163)
);

AOI22xp33_ASAP7_75t_L g5164 ( 
.A1(n_3254),
.A2(n_3260),
.B1(n_3276),
.B2(n_3262),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_4408),
.B(n_4414),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_SL g5166 ( 
.A(n_3270),
.B(n_3147),
.Y(n_5166)
);

BUFx6f_ASAP7_75t_L g5167 ( 
.A(n_3110),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_L g5168 ( 
.A(n_4414),
.B(n_4422),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4422),
.Y(n_5169)
);

NOR2xp33_ASAP7_75t_L g5170 ( 
.A(n_4464),
.B(n_3293),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_SL g5171 ( 
.A(n_3149),
.B(n_3150),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_4425),
.B(n_4429),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_4429),
.B(n_4431),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4431),
.Y(n_5174)
);

INVx5_ASAP7_75t_L g5175 ( 
.A(n_4201),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4446),
.Y(n_5176)
);

BUFx6f_ASAP7_75t_L g5177 ( 
.A(n_3110),
.Y(n_5177)
);

BUFx6f_ASAP7_75t_L g5178 ( 
.A(n_3120),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4446),
.Y(n_5179)
);

INVx5_ASAP7_75t_L g5180 ( 
.A(n_4360),
.Y(n_5180)
);

OR2x6_ASAP7_75t_L g5181 ( 
.A(n_3951),
.B(n_4036),
.Y(n_5181)
);

AOI22xp33_ASAP7_75t_L g5182 ( 
.A1(n_3276),
.A2(n_3281),
.B1(n_3288),
.B2(n_3286),
.Y(n_5182)
);

INVx2_ASAP7_75t_SL g5183 ( 
.A(n_3102),
.Y(n_5183)
);

AOI22xp5_ASAP7_75t_L g5184 ( 
.A1(n_3180),
.A2(n_3216),
.B1(n_3286),
.B2(n_3281),
.Y(n_5184)
);

AOI21xp33_ASAP7_75t_L g5185 ( 
.A1(n_3423),
.A2(n_3290),
.B(n_3288),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_3352),
.B(n_3356),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_3366),
.B(n_3381),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_3382),
.B(n_3388),
.Y(n_5188)
);

NOR2xp33_ASAP7_75t_L g5189 ( 
.A(n_3211),
.B(n_3231),
.Y(n_5189)
);

BUFx3_ASAP7_75t_L g5190 ( 
.A(n_3339),
.Y(n_5190)
);

BUFx12f_ASAP7_75t_L g5191 ( 
.A(n_4054),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_3348),
.Y(n_5192)
);

HB1xp67_ASAP7_75t_L g5193 ( 
.A(n_3984),
.Y(n_5193)
);

OR2x6_ASAP7_75t_L g5194 ( 
.A(n_4461),
.B(n_3963),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_3348),
.Y(n_5195)
);

AND3x1_ASAP7_75t_SL g5196 ( 
.A(n_3705),
.B(n_3708),
.C(n_4123),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_3390),
.B(n_3394),
.Y(n_5197)
);

BUFx4f_ASAP7_75t_L g5198 ( 
.A(n_4360),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_3211),
.B(n_3231),
.Y(n_5199)
);

OR2x6_ASAP7_75t_L g5200 ( 
.A(n_3930),
.B(n_3932),
.Y(n_5200)
);

INVxp67_ASAP7_75t_SL g5201 ( 
.A(n_3151),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_3365),
.Y(n_5202)
);

AOI221x1_ASAP7_75t_L g5203 ( 
.A1(n_3918),
.A2(n_3926),
.B1(n_3960),
.B2(n_3957),
.C(n_3937),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_3400),
.B(n_3410),
.Y(n_5204)
);

BUFx2_ASAP7_75t_L g5205 ( 
.A(n_4286),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_3413),
.B(n_3414),
.Y(n_5206)
);

AND2x6_ASAP7_75t_L g5207 ( 
.A(n_3602),
.B(n_3617),
.Y(n_5207)
);

BUFx2_ASAP7_75t_L g5208 ( 
.A(n_4286),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_3365),
.Y(n_5209)
);

NOR2xp33_ASAP7_75t_L g5210 ( 
.A(n_3239),
.B(n_3244),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_3522),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_3221),
.Y(n_5212)
);

OAI22xp5_ASAP7_75t_L g5213 ( 
.A1(n_3298),
.A2(n_3344),
.B1(n_3239),
.B2(n_3244),
.Y(n_5213)
);

BUFx4f_ASAP7_75t_L g5214 ( 
.A(n_4360),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_L g5215 ( 
.A(n_3422),
.B(n_3428),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_3221),
.Y(n_5216)
);

NOR2xp33_ASAP7_75t_L g5217 ( 
.A(n_3089),
.B(n_3210),
.Y(n_5217)
);

NOR2xp33_ASAP7_75t_L g5218 ( 
.A(n_3089),
.B(n_3229),
.Y(n_5218)
);

HB1xp67_ASAP7_75t_L g5219 ( 
.A(n_3984),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_3522),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_3433),
.B(n_3456),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_3227),
.Y(n_5222)
);

HB1xp67_ASAP7_75t_L g5223 ( 
.A(n_4016),
.Y(n_5223)
);

INVx4_ASAP7_75t_L g5224 ( 
.A(n_4013),
.Y(n_5224)
);

INVx4_ASAP7_75t_L g5225 ( 
.A(n_4169),
.Y(n_5225)
);

NOR2x1_ASAP7_75t_L g5226 ( 
.A(n_4116),
.B(n_4251),
.Y(n_5226)
);

HB1xp67_ASAP7_75t_L g5227 ( 
.A(n_4016),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_3543),
.Y(n_5228)
);

NAND2xp5_ASAP7_75t_L g5229 ( 
.A(n_3474),
.B(n_3450),
.Y(n_5229)
);

BUFx2_ASAP7_75t_L g5230 ( 
.A(n_4307),
.Y(n_5230)
);

OAI22xp5_ASAP7_75t_L g5231 ( 
.A1(n_3178),
.A2(n_3119),
.B1(n_3124),
.B2(n_3073),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_3170),
.B(n_3097),
.Y(n_5232)
);

BUFx12f_ASAP7_75t_L g5233 ( 
.A(n_4130),
.Y(n_5233)
);

BUFx2_ASAP7_75t_L g5234 ( 
.A(n_4307),
.Y(n_5234)
);

AOI22xp5_ASAP7_75t_L g5235 ( 
.A1(n_3216),
.A2(n_3290),
.B1(n_3294),
.B2(n_3291),
.Y(n_5235)
);

NAND2xp5_ASAP7_75t_SL g5236 ( 
.A(n_4126),
.B(n_4090),
.Y(n_5236)
);

CKINVDCx20_ASAP7_75t_R g5237 ( 
.A(n_4442),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_3170),
.B(n_3097),
.Y(n_5238)
);

INVxp67_ASAP7_75t_SL g5239 ( 
.A(n_3151),
.Y(n_5239)
);

OAI22xp5_ASAP7_75t_L g5240 ( 
.A1(n_3178),
.A2(n_3767),
.B1(n_3769),
.B2(n_3765),
.Y(n_5240)
);

INVx5_ASAP7_75t_L g5241 ( 
.A(n_4360),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_3543),
.Y(n_5242)
);

BUFx3_ASAP7_75t_L g5243 ( 
.A(n_3339),
.Y(n_5243)
);

BUFx6f_ASAP7_75t_L g5244 ( 
.A(n_3120),
.Y(n_5244)
);

BUFx3_ASAP7_75t_L g5245 ( 
.A(n_3339),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_3504),
.B(n_3453),
.Y(n_5246)
);

A2O1A1Ixp33_ASAP7_75t_L g5247 ( 
.A1(n_4193),
.A2(n_4233),
.B(n_3159),
.C(n_3172),
.Y(n_5247)
);

AND2x2_ASAP7_75t_L g5248 ( 
.A(n_4307),
.B(n_4312),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_3233),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_SL g5250 ( 
.A(n_3195),
.B(n_3242),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_3227),
.Y(n_5251)
);

BUFx6f_ASAP7_75t_L g5252 ( 
.A(n_3711),
.Y(n_5252)
);

BUFx4f_ASAP7_75t_L g5253 ( 
.A(n_4360),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_3504),
.B(n_3453),
.Y(n_5254)
);

BUFx6f_ASAP7_75t_L g5255 ( 
.A(n_3711),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_4312),
.B(n_4338),
.Y(n_5256)
);

AOI22xp5_ASAP7_75t_L g5257 ( 
.A1(n_3291),
.A2(n_3306),
.B1(n_3309),
.B2(n_3294),
.Y(n_5257)
);

BUFx6f_ASAP7_75t_L g5258 ( 
.A(n_3731),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_3233),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_3457),
.B(n_3427),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_3427),
.B(n_3436),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_3436),
.B(n_3165),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_3176),
.B(n_3323),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_3361),
.B(n_3490),
.Y(n_5264)
);

BUFx2_ASAP7_75t_L g5265 ( 
.A(n_4338),
.Y(n_5265)
);

BUFx6f_ASAP7_75t_L g5266 ( 
.A(n_3731),
.Y(n_5266)
);

OR2x2_ASAP7_75t_L g5267 ( 
.A(n_4016),
.B(n_4393),
.Y(n_5267)
);

OAI21xp33_ASAP7_75t_L g5268 ( 
.A1(n_3129),
.A2(n_3168),
.B(n_3162),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_3361),
.B(n_3490),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_3712),
.B(n_3762),
.Y(n_5270)
);

AOI22xp33_ASAP7_75t_L g5271 ( 
.A1(n_3306),
.A2(n_3309),
.B1(n_3319),
.B2(n_3310),
.Y(n_5271)
);

BUFx2_ASAP7_75t_L g5272 ( 
.A(n_4348),
.Y(n_5272)
);

AND3x1_ASAP7_75t_SL g5273 ( 
.A(n_3705),
.B(n_3708),
.C(n_4226),
.Y(n_5273)
);

CKINVDCx20_ASAP7_75t_R g5274 ( 
.A(n_4442),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_3235),
.Y(n_5275)
);

INVx4_ASAP7_75t_L g5276 ( 
.A(n_4169),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_3712),
.B(n_3762),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_3235),
.Y(n_5278)
);

AND2x6_ASAP7_75t_L g5279 ( 
.A(n_3602),
.B(n_3617),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_3886),
.B(n_4248),
.Y(n_5280)
);

CKINVDCx8_ASAP7_75t_R g5281 ( 
.A(n_3339),
.Y(n_5281)
);

BUFx4f_ASAP7_75t_L g5282 ( 
.A(n_4360),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_3886),
.B(n_4248),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_4143),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_4275),
.B(n_4283),
.Y(n_5285)
);

INVx2_ASAP7_75t_L g5286 ( 
.A(n_3227),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_3250),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_3250),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_3273),
.Y(n_5289)
);

INVx2_ASAP7_75t_L g5290 ( 
.A(n_4016),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_4275),
.B(n_4283),
.Y(n_5291)
);

INVx4_ASAP7_75t_L g5292 ( 
.A(n_4169),
.Y(n_5292)
);

AOI211xp5_ASAP7_75t_L g5293 ( 
.A1(n_3168),
.A2(n_4316),
.B(n_3202),
.C(n_3495),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_4393),
.Y(n_5294)
);

AOI22xp33_ASAP7_75t_L g5295 ( 
.A1(n_3310),
.A2(n_3319),
.B1(n_3322),
.B2(n_3321),
.Y(n_5295)
);

NOR2xp33_ASAP7_75t_L g5296 ( 
.A(n_3194),
.B(n_3253),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_3273),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_4393),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_4393),
.Y(n_5299)
);

BUFx6f_ASAP7_75t_L g5300 ( 
.A(n_3799),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_3514),
.Y(n_5301)
);

AOI22x1_ASAP7_75t_L g5302 ( 
.A1(n_3964),
.A2(n_3970),
.B1(n_3978),
.B2(n_3974),
.Y(n_5302)
);

HB1xp67_ASAP7_75t_L g5303 ( 
.A(n_3514),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_4288),
.B(n_3321),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_4288),
.B(n_3322),
.Y(n_5305)
);

HB1xp67_ASAP7_75t_L g5306 ( 
.A(n_3199),
.Y(n_5306)
);

BUFx2_ASAP7_75t_L g5307 ( 
.A(n_4375),
.Y(n_5307)
);

INVx4_ASAP7_75t_L g5308 ( 
.A(n_4246),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_SL g5309 ( 
.A(n_3242),
.B(n_3980),
.Y(n_5309)
);

OR2x2_ASAP7_75t_L g5310 ( 
.A(n_3327),
.B(n_3358),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_3327),
.B(n_3358),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_3359),
.B(n_3367),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_3359),
.B(n_3367),
.Y(n_5313)
);

HB1xp67_ASAP7_75t_L g5314 ( 
.A(n_3238),
.Y(n_5314)
);

BUFx2_ASAP7_75t_L g5315 ( 
.A(n_4472),
.Y(n_5315)
);

AOI221xp5_ASAP7_75t_L g5316 ( 
.A1(n_3296),
.A2(n_3207),
.B1(n_3311),
.B2(n_3376),
.C(n_3373),
.Y(n_5316)
);

AND2x4_ASAP7_75t_L g5317 ( 
.A(n_4472),
.B(n_4450),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_4472),
.Y(n_5318)
);

CKINVDCx5p33_ASAP7_75t_R g5319 ( 
.A(n_4350),
.Y(n_5319)
);

INVx3_ASAP7_75t_L g5320 ( 
.A(n_3945),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_3373),
.B(n_3377),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_3295),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_3376),
.B(n_3377),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_3378),
.B(n_3379),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_3378),
.B(n_3379),
.Y(n_5325)
);

BUFx6f_ASAP7_75t_L g5326 ( 
.A(n_3799),
.Y(n_5326)
);

INVx2_ASAP7_75t_L g5327 ( 
.A(n_3314),
.Y(n_5327)
);

AOI22xp5_ASAP7_75t_SL g5328 ( 
.A1(n_3495),
.A2(n_3275),
.B1(n_3628),
.B2(n_3300),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_3406),
.B(n_3417),
.Y(n_5329)
);

AND2x2_ASAP7_75t_L g5330 ( 
.A(n_3471),
.B(n_3326),
.Y(n_5330)
);

HB1xp67_ASAP7_75t_L g5331 ( 
.A(n_3246),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_3425),
.B(n_3307),
.Y(n_5332)
);

INVx4_ASAP7_75t_SL g5333 ( 
.A(n_4360),
.Y(n_5333)
);

BUFx3_ASAP7_75t_L g5334 ( 
.A(n_3100),
.Y(n_5334)
);

OR2x6_ASAP7_75t_L g5335 ( 
.A(n_4441),
.B(n_4026),
.Y(n_5335)
);

OAI22xp5_ASAP7_75t_L g5336 ( 
.A1(n_3770),
.A2(n_3785),
.B1(n_3787),
.B2(n_3776),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_SL g5337 ( 
.A(n_3989),
.B(n_4006),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_3334),
.Y(n_5338)
);

INVx2_ASAP7_75t_L g5339 ( 
.A(n_3337),
.Y(n_5339)
);

BUFx2_ASAP7_75t_L g5340 ( 
.A(n_3091),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_3318),
.B(n_3338),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_3362),
.B(n_3370),
.Y(n_5342)
);

AOI22xp33_ASAP7_75t_L g5343 ( 
.A1(n_3439),
.A2(n_3272),
.B1(n_3258),
.B2(n_3790),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_3337),
.Y(n_5344)
);

AO22x1_ASAP7_75t_L g5345 ( 
.A1(n_4130),
.A2(n_4158),
.B1(n_4232),
.B2(n_4246),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_SL g5346 ( 
.A(n_4022),
.B(n_4027),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_SL g5347 ( 
.A(n_4028),
.B(n_4042),
.Y(n_5347)
);

NOR2xp33_ASAP7_75t_L g5348 ( 
.A(n_3792),
.B(n_3798),
.Y(n_5348)
);

BUFx12f_ASAP7_75t_L g5349 ( 
.A(n_4130),
.Y(n_5349)
);

BUFx2_ASAP7_75t_L g5350 ( 
.A(n_3091),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_3402),
.B(n_3432),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_3460),
.B(n_3183),
.Y(n_5352)
);

INVxp67_ASAP7_75t_SL g5353 ( 
.A(n_3445),
.Y(n_5353)
);

INVx3_ASAP7_75t_L g5354 ( 
.A(n_3945),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_3357),
.Y(n_5355)
);

AND2x4_ASAP7_75t_L g5356 ( 
.A(n_4450),
.B(n_3102),
.Y(n_5356)
);

AND3x1_ASAP7_75t_SL g5357 ( 
.A(n_3682),
.B(n_3648),
.C(n_4350),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_3403),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_3720),
.B(n_3726),
.Y(n_5359)
);

AOI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_3399),
.A2(n_3484),
.B1(n_3439),
.B2(n_3801),
.Y(n_5360)
);

AND2x2_ASAP7_75t_L g5361 ( 
.A(n_3471),
.B(n_3405),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_3421),
.Y(n_5362)
);

INVx2_ASAP7_75t_L g5363 ( 
.A(n_3421),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_3726),
.B(n_3783),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_L g5365 ( 
.A(n_3783),
.B(n_3844),
.Y(n_5365)
);

AND2x6_ASAP7_75t_L g5366 ( 
.A(n_3602),
.B(n_3617),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_3844),
.B(n_3851),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_3851),
.B(n_3884),
.Y(n_5368)
);

INVx4_ASAP7_75t_L g5369 ( 
.A(n_4246),
.Y(n_5369)
);

OAI22xp33_ASAP7_75t_L g5370 ( 
.A1(n_3805),
.A2(n_3820),
.B1(n_4474),
.B2(n_3806),
.Y(n_5370)
);

HB1xp67_ASAP7_75t_L g5371 ( 
.A(n_3331),
.Y(n_5371)
);

AND2x2_ASAP7_75t_L g5372 ( 
.A(n_3430),
.B(n_3441),
.Y(n_5372)
);

BUFx2_ASAP7_75t_L g5373 ( 
.A(n_3096),
.Y(n_5373)
);

BUFx6f_ASAP7_75t_L g5374 ( 
.A(n_3803),
.Y(n_5374)
);

BUFx3_ASAP7_75t_L g5375 ( 
.A(n_3100),
.Y(n_5375)
);

AOI21xp5_ASAP7_75t_L g5376 ( 
.A1(n_4044),
.A2(n_4062),
.B(n_4056),
.Y(n_5376)
);

INVx2_ASAP7_75t_L g5377 ( 
.A(n_3430),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_3884),
.B(n_4020),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_4020),
.B(n_4280),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_3441),
.Y(n_5380)
);

INVx2_ASAP7_75t_SL g5381 ( 
.A(n_3102),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_3452),
.Y(n_5382)
);

HB1xp67_ASAP7_75t_L g5383 ( 
.A(n_3389),
.Y(n_5383)
);

NOR2xp33_ASAP7_75t_L g5384 ( 
.A(n_3446),
.B(n_3401),
.Y(n_5384)
);

HB1xp67_ASAP7_75t_L g5385 ( 
.A(n_3443),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_4280),
.B(n_4383),
.Y(n_5386)
);

NOR2xp33_ASAP7_75t_L g5387 ( 
.A(n_3404),
.B(n_3511),
.Y(n_5387)
);

BUFx6f_ASAP7_75t_L g5388 ( 
.A(n_3803),
.Y(n_5388)
);

CKINVDCx5p33_ASAP7_75t_R g5389 ( 
.A(n_4413),
.Y(n_5389)
);

NOR4xp25_ASAP7_75t_SL g5390 ( 
.A(n_3628),
.B(n_3511),
.C(n_3745),
.D(n_3482),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_3452),
.Y(n_5391)
);

OAI22xp5_ASAP7_75t_L g5392 ( 
.A1(n_3473),
.A2(n_3472),
.B1(n_3447),
.B2(n_3343),
.Y(n_5392)
);

BUFx3_ASAP7_75t_L g5393 ( 
.A(n_3100),
.Y(n_5393)
);

BUFx4f_ASAP7_75t_L g5394 ( 
.A(n_4360),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_3096),
.Y(n_5395)
);

INVx2_ASAP7_75t_L g5396 ( 
.A(n_3113),
.Y(n_5396)
);

AND2x2_ASAP7_75t_SL g5397 ( 
.A(n_3556),
.B(n_3588),
.Y(n_5397)
);

AND2x4_ASAP7_75t_L g5398 ( 
.A(n_3102),
.B(n_3154),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_3113),
.Y(n_5399)
);

NAND2xp5_ASAP7_75t_L g5400 ( 
.A(n_4383),
.B(n_3956),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_3241),
.Y(n_5401)
);

BUFx3_ASAP7_75t_L g5402 ( 
.A(n_4052),
.Y(n_5402)
);

NAND2xp5_ASAP7_75t_L g5403 ( 
.A(n_3956),
.B(n_3967),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_3241),
.Y(n_5404)
);

INVx3_ASAP7_75t_L g5405 ( 
.A(n_4371),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_3598),
.Y(n_5406)
);

BUFx6f_ASAP7_75t_L g5407 ( 
.A(n_3967),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_3464),
.Y(n_5408)
);

HB1xp67_ASAP7_75t_L g5409 ( 
.A(n_3451),
.Y(n_5409)
);

HB1xp67_ASAP7_75t_L g5410 ( 
.A(n_3814),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_3464),
.Y(n_5411)
);

AND2x2_ASAP7_75t_L g5412 ( 
.A(n_3498),
.B(n_3215),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_4110),
.B(n_4325),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_4110),
.B(n_4325),
.Y(n_5414)
);

AND2x2_ASAP7_75t_L g5415 ( 
.A(n_3498),
.B(n_3215),
.Y(n_5415)
);

INVx2_ASAP7_75t_L g5416 ( 
.A(n_3598),
.Y(n_5416)
);

INVx3_ASAP7_75t_L g5417 ( 
.A(n_4371),
.Y(n_5417)
);

INVx4_ASAP7_75t_L g5418 ( 
.A(n_4246),
.Y(n_5418)
);

AOI22xp5_ASAP7_75t_L g5419 ( 
.A1(n_3481),
.A2(n_3512),
.B1(n_3418),
.B2(n_3272),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_4452),
.B(n_4456),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_3469),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_3647),
.Y(n_5422)
);

AND2x2_ASAP7_75t_L g5423 ( 
.A(n_3499),
.B(n_3520),
.Y(n_5423)
);

NAND2xp5_ASAP7_75t_SL g5424 ( 
.A(n_4063),
.B(n_4064),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_3469),
.Y(n_5425)
);

INVx2_ASAP7_75t_SL g5426 ( 
.A(n_3154),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_SL g5427 ( 
.A(n_4065),
.B(n_4068),
.Y(n_5427)
);

NAND2x1p5_ASAP7_75t_L g5428 ( 
.A(n_4116),
.B(n_4251),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_3647),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_4452),
.B(n_4456),
.Y(n_5430)
);

BUFx6f_ASAP7_75t_L g5431 ( 
.A(n_4263),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_3657),
.Y(n_5432)
);

AOI21xp5_ASAP7_75t_L g5433 ( 
.A1(n_4071),
.A2(n_4084),
.B(n_4078),
.Y(n_5433)
);

OR2x2_ASAP7_75t_L g5434 ( 
.A(n_3936),
.B(n_4156),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_3476),
.Y(n_5435)
);

CKINVDCx5p33_ASAP7_75t_R g5436 ( 
.A(n_4413),
.Y(n_5436)
);

AOI22x1_ASAP7_75t_L g5437 ( 
.A1(n_4089),
.A2(n_4091),
.B1(n_4109),
.B2(n_4096),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_3279),
.B(n_3299),
.Y(n_5438)
);

HB1xp67_ASAP7_75t_L g5439 ( 
.A(n_4171),
.Y(n_5439)
);

BUFx3_ASAP7_75t_L g5440 ( 
.A(n_4052),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_3657),
.Y(n_5441)
);

INVx2_ASAP7_75t_L g5442 ( 
.A(n_3312),
.Y(n_5442)
);

NOR2xp33_ASAP7_75t_L g5443 ( 
.A(n_3384),
.B(n_3387),
.Y(n_5443)
);

CKINVDCx20_ASAP7_75t_R g5444 ( 
.A(n_4130),
.Y(n_5444)
);

AOI21xp5_ASAP7_75t_L g5445 ( 
.A1(n_4114),
.A2(n_4127),
.B(n_4124),
.Y(n_5445)
);

AOI22xp5_ASAP7_75t_L g5446 ( 
.A1(n_3473),
.A2(n_3466),
.B1(n_3369),
.B2(n_3375),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_3279),
.B(n_3299),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_3476),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_3477),
.Y(n_5449)
);

HB1xp67_ASAP7_75t_L g5450 ( 
.A(n_4308),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_3335),
.B(n_3397),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_3477),
.Y(n_5452)
);

NOR2xp33_ASAP7_75t_L g5453 ( 
.A(n_3384),
.B(n_3387),
.Y(n_5453)
);

AND3x1_ASAP7_75t_SL g5454 ( 
.A(n_3682),
.B(n_3648),
.C(n_3546),
.Y(n_5454)
);

AOI22xp5_ASAP7_75t_L g5455 ( 
.A1(n_3364),
.A2(n_3383),
.B1(n_3396),
.B2(n_3380),
.Y(n_5455)
);

BUFx3_ASAP7_75t_L g5456 ( 
.A(n_4052),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_3479),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_3335),
.B(n_3397),
.Y(n_5458)
);

NAND2xp5_ASAP7_75t_L g5459 ( 
.A(n_3415),
.B(n_4367),
.Y(n_5459)
);

OR2x4_ASAP7_75t_L g5460 ( 
.A(n_3524),
.B(n_3638),
.Y(n_5460)
);

INVx2_ASAP7_75t_L g5461 ( 
.A(n_3312),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_3479),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_3467),
.Y(n_5463)
);

OAI22xp5_ASAP7_75t_SL g5464 ( 
.A1(n_3472),
.A2(n_3255),
.B1(n_4263),
.B2(n_3501),
.Y(n_5464)
);

AOI22x1_ASAP7_75t_L g5465 ( 
.A1(n_4129),
.A2(n_4140),
.B1(n_4148),
.B2(n_4132),
.Y(n_5465)
);

INVx1_ASAP7_75t_SL g5466 ( 
.A(n_3524),
.Y(n_5466)
);

AOI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_3408),
.A2(n_3435),
.B1(n_3223),
.B2(n_3341),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_3154),
.Y(n_5468)
);

INVx2_ASAP7_75t_SL g5469 ( 
.A(n_3154),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_3489),
.Y(n_5470)
);

CKINVDCx5p33_ASAP7_75t_R g5471 ( 
.A(n_3467),
.Y(n_5471)
);

BUFx3_ASAP7_75t_L g5472 ( 
.A(n_4066),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_3393),
.B(n_3409),
.Y(n_5473)
);

AND2x2_ASAP7_75t_SL g5474 ( 
.A(n_3556),
.B(n_3588),
.Y(n_5474)
);

OR2x6_ASAP7_75t_L g5475 ( 
.A(n_4149),
.B(n_4152),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_3489),
.Y(n_5476)
);

AOI22xp5_ASAP7_75t_L g5477 ( 
.A1(n_3223),
.A2(n_3341),
.B1(n_3372),
.B2(n_3316),
.Y(n_5477)
);

AND2x4_ASAP7_75t_L g5478 ( 
.A(n_3748),
.B(n_3866),
.Y(n_5478)
);

HB1xp67_ASAP7_75t_L g5479 ( 
.A(n_4420),
.Y(n_5479)
);

O2A1O1Ixp33_ASAP7_75t_L g5480 ( 
.A1(n_3346),
.A2(n_4160),
.B(n_4163),
.C(n_4154),
.Y(n_5480)
);

AOI22xp5_ASAP7_75t_L g5481 ( 
.A1(n_3316),
.A2(n_3411),
.B1(n_3454),
.B2(n_3372),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_3497),
.Y(n_5482)
);

AND2x4_ASAP7_75t_L g5483 ( 
.A(n_3748),
.B(n_3866),
.Y(n_5483)
);

AND2x2_ASAP7_75t_L g5484 ( 
.A(n_3499),
.B(n_3520),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_L g5485 ( 
.A(n_3415),
.B(n_4445),
.Y(n_5485)
);

CKINVDCx5p33_ASAP7_75t_R g5486 ( 
.A(n_3768),
.Y(n_5486)
);

BUFx3_ASAP7_75t_L g5487 ( 
.A(n_4066),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_3497),
.Y(n_5488)
);

AOI22xp5_ASAP7_75t_L g5489 ( 
.A1(n_3411),
.A2(n_3454),
.B1(n_3409),
.B2(n_3412),
.Y(n_5489)
);

AND2x2_ASAP7_75t_L g5490 ( 
.A(n_4263),
.B(n_3748),
.Y(n_5490)
);

NAND2xp5_ASAP7_75t_L g5491 ( 
.A(n_3313),
.B(n_3351),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_3374),
.B(n_3416),
.Y(n_5492)
);

INVxp67_ASAP7_75t_L g5493 ( 
.A(n_4416),
.Y(n_5493)
);

CKINVDCx8_ASAP7_75t_R g5494 ( 
.A(n_3602),
.Y(n_5494)
);

AND2x2_ASAP7_75t_L g5495 ( 
.A(n_4263),
.B(n_3748),
.Y(n_5495)
);

CKINVDCx5p33_ASAP7_75t_R g5496 ( 
.A(n_3768),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_3434),
.B(n_4173),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_4175),
.B(n_4180),
.Y(n_5498)
);

AOI22xp33_ASAP7_75t_L g5499 ( 
.A1(n_3438),
.A2(n_3455),
.B1(n_3463),
.B2(n_3412),
.Y(n_5499)
);

NOR2xp33_ASAP7_75t_L g5500 ( 
.A(n_3393),
.B(n_3419),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_4182),
.B(n_4189),
.Y(n_5501)
);

HB1xp67_ASAP7_75t_L g5502 ( 
.A(n_4416),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_3502),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_4195),
.B(n_4196),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_3502),
.Y(n_5505)
);

OAI22xp5_ASAP7_75t_SL g5506 ( 
.A1(n_3501),
.A2(n_4100),
.B1(n_4361),
.B2(n_3943),
.Y(n_5506)
);

AND2x2_ASAP7_75t_L g5507 ( 
.A(n_3866),
.B(n_4024),
.Y(n_5507)
);

HB1xp67_ASAP7_75t_L g5508 ( 
.A(n_3445),
.Y(n_5508)
);

NOR2x1_ASAP7_75t_L g5509 ( 
.A(n_4202),
.B(n_4205),
.Y(n_5509)
);

AND3x1_ASAP7_75t_SL g5510 ( 
.A(n_3546),
.B(n_4232),
.C(n_4158),
.Y(n_5510)
);

AND2x2_ASAP7_75t_L g5511 ( 
.A(n_3866),
.B(n_4024),
.Y(n_5511)
);

BUFx6f_ASAP7_75t_L g5512 ( 
.A(n_4066),
.Y(n_5512)
);

BUFx6f_ASAP7_75t_L g5513 ( 
.A(n_4162),
.Y(n_5513)
);

NAND2xp33_ASAP7_75t_L g5514 ( 
.A(n_4212),
.B(n_4215),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_4219),
.B(n_4220),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_L g5516 ( 
.A(n_4221),
.B(n_4225),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_3505),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_3505),
.Y(n_5518)
);

A2O1A1Ixp33_ASAP7_75t_L g5519 ( 
.A1(n_4229),
.A2(n_4475),
.B(n_4230),
.C(n_4236),
.Y(n_5519)
);

INVxp67_ASAP7_75t_SL g5520 ( 
.A(n_4234),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_3516),
.Y(n_5521)
);

NOR2xp33_ASAP7_75t_L g5522 ( 
.A(n_3419),
.B(n_3420),
.Y(n_5522)
);

AOI22x1_ASAP7_75t_L g5523 ( 
.A1(n_4240),
.A2(n_4247),
.B1(n_4256),
.B2(n_4255),
.Y(n_5523)
);

AOI22xp33_ASAP7_75t_L g5524 ( 
.A1(n_3455),
.A2(n_3437),
.B1(n_3420),
.B2(n_3330),
.Y(n_5524)
);

A2O1A1Ixp33_ASAP7_75t_L g5525 ( 
.A1(n_4278),
.A2(n_4289),
.B(n_4306),
.C(n_4302),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_3516),
.Y(n_5526)
);

AND2x4_ASAP7_75t_L g5527 ( 
.A(n_4024),
.B(n_4112),
.Y(n_5527)
);

NAND2xp33_ASAP7_75t_L g5528 ( 
.A(n_4310),
.B(n_4327),
.Y(n_5528)
);

INVx2_ASAP7_75t_SL g5529 ( 
.A(n_4024),
.Y(n_5529)
);

NAND2xp5_ASAP7_75t_L g5530 ( 
.A(n_4330),
.B(n_4334),
.Y(n_5530)
);

AND2x2_ASAP7_75t_L g5531 ( 
.A(n_4112),
.B(n_4450),
.Y(n_5531)
);

BUFx3_ASAP7_75t_L g5532 ( 
.A(n_4162),
.Y(n_5532)
);

HB1xp67_ASAP7_75t_L g5533 ( 
.A(n_3287),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_3521),
.Y(n_5534)
);

INVx1_ASAP7_75t_SL g5535 ( 
.A(n_3131),
.Y(n_5535)
);

OAI22xp5_ASAP7_75t_L g5536 ( 
.A1(n_4335),
.A2(n_4347),
.B1(n_4363),
.B2(n_4355),
.Y(n_5536)
);

INVx1_ASAP7_75t_SL g5537 ( 
.A(n_3131),
.Y(n_5537)
);

BUFx4f_ASAP7_75t_L g5538 ( 
.A(n_4162),
.Y(n_5538)
);

CKINVDCx5p33_ASAP7_75t_R g5539 ( 
.A(n_3768),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_SL g5540 ( 
.A(n_4366),
.B(n_4368),
.Y(n_5540)
);

NOR2xp33_ASAP7_75t_L g5541 ( 
.A(n_3437),
.B(n_3475),
.Y(n_5541)
);

INVx4_ASAP7_75t_L g5542 ( 
.A(n_3729),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_3521),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_3529),
.Y(n_5544)
);

BUFx6f_ASAP7_75t_L g5545 ( 
.A(n_3117),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_4369),
.B(n_4373),
.Y(n_5546)
);

CKINVDCx8_ASAP7_75t_R g5547 ( 
.A(n_3617),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_3529),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_4376),
.B(n_4377),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_3530),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_3530),
.Y(n_5551)
);

NAND2xp5_ASAP7_75t_SL g5552 ( 
.A(n_4378),
.B(n_4380),
.Y(n_5552)
);

CKINVDCx5p33_ASAP7_75t_R g5553 ( 
.A(n_3881),
.Y(n_5553)
);

INVx3_ASAP7_75t_L g5554 ( 
.A(n_4112),
.Y(n_5554)
);

BUFx3_ASAP7_75t_L g5555 ( 
.A(n_3556),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_4112),
.B(n_4450),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_3542),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_3556),
.Y(n_5558)
);

AOI22xp33_ASAP7_75t_L g5559 ( 
.A1(n_3328),
.A2(n_3333),
.B1(n_3336),
.B2(n_3332),
.Y(n_5559)
);

CKINVDCx5p33_ASAP7_75t_R g5560 ( 
.A(n_3881),
.Y(n_5560)
);

INVxp67_ASAP7_75t_L g5561 ( 
.A(n_3542),
.Y(n_5561)
);

BUFx2_ASAP7_75t_L g5562 ( 
.A(n_3729),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_4390),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_4394),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_4395),
.B(n_4399),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_SL g5566 ( 
.A(n_4400),
.B(n_4405),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_4421),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_4423),
.Y(n_5568)
);

NAND2xp5_ASAP7_75t_L g5569 ( 
.A(n_4434),
.B(n_4435),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_4436),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_SL g5571 ( 
.A(n_4437),
.B(n_4438),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_4440),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_4454),
.B(n_3305),
.Y(n_5573)
);

AND2x2_ASAP7_75t_L g5574 ( 
.A(n_3559),
.B(n_3738),
.Y(n_5574)
);

BUFx4f_ASAP7_75t_SL g5575 ( 
.A(n_3881),
.Y(n_5575)
);

INVx3_ASAP7_75t_L g5576 ( 
.A(n_3738),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_3340),
.B(n_3407),
.Y(n_5577)
);

BUFx2_ASAP7_75t_L g5578 ( 
.A(n_3738),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_3287),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_3483),
.B(n_3503),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_3507),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_SL g5582 ( 
.A(n_3525),
.B(n_3527),
.Y(n_5582)
);

INVx3_ASAP7_75t_L g5583 ( 
.A(n_3738),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_3509),
.B(n_3515),
.Y(n_5584)
);

BUFx3_ASAP7_75t_L g5585 ( 
.A(n_3588),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_3518),
.Y(n_5586)
);

CKINVDCx8_ASAP7_75t_R g5587 ( 
.A(n_3523),
.Y(n_5587)
);

CKINVDCx5p33_ASAP7_75t_R g5588 ( 
.A(n_4318),
.Y(n_5588)
);

INVxp67_ASAP7_75t_L g5589 ( 
.A(n_3559),
.Y(n_5589)
);

NOR2xp33_ASAP7_75t_L g5590 ( 
.A(n_3548),
.B(n_3564),
.Y(n_5590)
);

NAND2xp5_ASAP7_75t_L g5591 ( 
.A(n_3528),
.B(n_3531),
.Y(n_5591)
);

NAND2xp5_ASAP7_75t_L g5592 ( 
.A(n_3535),
.B(n_3536),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_3620),
.Y(n_5593)
);

CKINVDCx5p33_ASAP7_75t_R g5594 ( 
.A(n_4318),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_3620),
.Y(n_5595)
);

BUFx4f_ASAP7_75t_L g5596 ( 
.A(n_3117),
.Y(n_5596)
);

INVx5_ASAP7_75t_L g5597 ( 
.A(n_3837),
.Y(n_5597)
);

BUFx2_ASAP7_75t_L g5598 ( 
.A(n_4467),
.Y(n_5598)
);

AOI22xp5_ASAP7_75t_L g5599 ( 
.A1(n_3555),
.A2(n_3492),
.B1(n_3347),
.B2(n_3461),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_3634),
.Y(n_5600)
);

HB1xp67_ASAP7_75t_L g5601 ( 
.A(n_3213),
.Y(n_5601)
);

NAND2xp5_ASAP7_75t_L g5602 ( 
.A(n_3317),
.B(n_3324),
.Y(n_5602)
);

AND2x2_ASAP7_75t_L g5603 ( 
.A(n_3837),
.B(n_3887),
.Y(n_5603)
);

NOR2xp67_ASAP7_75t_L g5604 ( 
.A(n_3544),
.B(n_3565),
.Y(n_5604)
);

BUFx6f_ASAP7_75t_L g5605 ( 
.A(n_3117),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_3634),
.Y(n_5606)
);

AO22x1_ASAP7_75t_L g5607 ( 
.A1(n_4158),
.A2(n_4232),
.B1(n_3670),
.B2(n_3614),
.Y(n_5607)
);

BUFx6f_ASAP7_75t_L g5608 ( 
.A(n_3117),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_3470),
.B(n_3526),
.Y(n_5609)
);

INVx1_ASAP7_75t_SL g5610 ( 
.A(n_3153),
.Y(n_5610)
);

INVx3_ASAP7_75t_L g5611 ( 
.A(n_3837),
.Y(n_5611)
);

AND2x2_ASAP7_75t_L g5612 ( 
.A(n_3837),
.B(n_3887),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_L g5613 ( 
.A(n_3525),
.B(n_3527),
.Y(n_5613)
);

INVx3_ASAP7_75t_L g5614 ( 
.A(n_3887),
.Y(n_5614)
);

NOR2xp67_ASAP7_75t_L g5615 ( 
.A(n_3565),
.B(n_3632),
.Y(n_5615)
);

BUFx3_ASAP7_75t_L g5616 ( 
.A(n_3588),
.Y(n_5616)
);

BUFx3_ASAP7_75t_L g5617 ( 
.A(n_3213),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_SL g5618 ( 
.A(n_3347),
.B(n_3462),
.Y(n_5618)
);

NOR3xp33_ASAP7_75t_L g5619 ( 
.A(n_3641),
.B(n_3568),
.C(n_3586),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_SL g5620 ( 
.A(n_3568),
.B(n_3900),
.Y(n_5620)
);

BUFx6f_ASAP7_75t_L g5621 ( 
.A(n_3117),
.Y(n_5621)
);

AND2x2_ASAP7_75t_L g5622 ( 
.A(n_3900),
.B(n_3925),
.Y(n_5622)
);

BUFx3_ASAP7_75t_L g5623 ( 
.A(n_3213),
.Y(n_5623)
);

NAND2xp5_ASAP7_75t_L g5624 ( 
.A(n_3153),
.B(n_3201),
.Y(n_5624)
);

NAND2xp5_ASAP7_75t_SL g5625 ( 
.A(n_3925),
.B(n_3958),
.Y(n_5625)
);

AOI22xp5_ASAP7_75t_L g5626 ( 
.A1(n_3574),
.A2(n_3534),
.B1(n_3714),
.B2(n_3196),
.Y(n_5626)
);

BUFx3_ASAP7_75t_L g5627 ( 
.A(n_3925),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_3201),
.B(n_3204),
.Y(n_5628)
);

BUFx6f_ASAP7_75t_L g5629 ( 
.A(n_3117),
.Y(n_5629)
);

AND2x4_ASAP7_75t_L g5630 ( 
.A(n_3925),
.B(n_3958),
.Y(n_5630)
);

INVxp67_ASAP7_75t_SL g5631 ( 
.A(n_3566),
.Y(n_5631)
);

AND2x4_ASAP7_75t_L g5632 ( 
.A(n_3958),
.B(n_4150),
.Y(n_5632)
);

A2O1A1Ixp33_ASAP7_75t_L g5633 ( 
.A1(n_3614),
.A2(n_3491),
.B(n_3607),
.C(n_3561),
.Y(n_5633)
);

AND2x2_ASAP7_75t_L g5634 ( 
.A(n_4150),
.B(n_4227),
.Y(n_5634)
);

NAND2xp5_ASAP7_75t_L g5635 ( 
.A(n_3204),
.B(n_3251),
.Y(n_5635)
);

AOI21xp5_ASAP7_75t_L g5636 ( 
.A1(n_4150),
.A2(n_4296),
.B(n_4227),
.Y(n_5636)
);

NOR2xp33_ASAP7_75t_L g5637 ( 
.A(n_3485),
.B(n_3586),
.Y(n_5637)
);

AOI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_4150),
.A2(n_4296),
.B(n_4227),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_3251),
.B(n_3558),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_3558),
.B(n_3315),
.Y(n_5640)
);

INVx4_ASAP7_75t_L g5641 ( 
.A(n_4227),
.Y(n_5641)
);

NOR2xp33_ASAP7_75t_L g5642 ( 
.A(n_3573),
.B(n_3673),
.Y(n_5642)
);

CKINVDCx16_ASAP7_75t_R g5643 ( 
.A(n_3565),
.Y(n_5643)
);

NAND2xp33_ASAP7_75t_L g5644 ( 
.A(n_4296),
.B(n_4297),
.Y(n_5644)
);

BUFx2_ASAP7_75t_L g5645 ( 
.A(n_4296),
.Y(n_5645)
);

AOI22xp33_ASAP7_75t_L g5646 ( 
.A1(n_3496),
.A2(n_3671),
.B1(n_3670),
.B2(n_3653),
.Y(n_5646)
);

OR2x2_ASAP7_75t_L g5647 ( 
.A(n_3973),
.B(n_4032),
.Y(n_5647)
);

INVxp67_ASAP7_75t_SL g5648 ( 
.A(n_4297),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_3315),
.B(n_4297),
.Y(n_5649)
);

NAND2xp5_ASAP7_75t_SL g5650 ( 
.A(n_4297),
.B(n_4322),
.Y(n_5650)
);

INVx2_ASAP7_75t_SL g5651 ( 
.A(n_4322),
.Y(n_5651)
);

AND2x2_ASAP7_75t_L g5652 ( 
.A(n_4322),
.B(n_4460),
.Y(n_5652)
);

NAND2xp5_ASAP7_75t_L g5653 ( 
.A(n_4322),
.B(n_4460),
.Y(n_5653)
);

INVxp67_ASAP7_75t_SL g5654 ( 
.A(n_4460),
.Y(n_5654)
);

NOR2xp33_ASAP7_75t_L g5655 ( 
.A(n_3673),
.B(n_3668),
.Y(n_5655)
);

INVx2_ASAP7_75t_SL g5656 ( 
.A(n_4460),
.Y(n_5656)
);

NAND2xp5_ASAP7_75t_L g5657 ( 
.A(n_4467),
.B(n_3553),
.Y(n_5657)
);

NOR2xp33_ASAP7_75t_L g5658 ( 
.A(n_3668),
.B(n_3638),
.Y(n_5658)
);

NAND2xp5_ASAP7_75t_L g5659 ( 
.A(n_3664),
.B(n_3540),
.Y(n_5659)
);

NAND2xp5_ASAP7_75t_SL g5660 ( 
.A(n_3137),
.B(n_3266),
.Y(n_5660)
);

BUFx6f_ASAP7_75t_L g5661 ( 
.A(n_3137),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_3664),
.B(n_3554),
.Y(n_5662)
);

NOR2xp33_ASAP7_75t_L g5663 ( 
.A(n_3668),
.B(n_3638),
.Y(n_5663)
);

NOR2xp33_ASAP7_75t_L g5664 ( 
.A(n_3668),
.B(n_3638),
.Y(n_5664)
);

AND3x1_ASAP7_75t_SL g5665 ( 
.A(n_3546),
.B(n_4232),
.C(n_4158),
.Y(n_5665)
);

INVx5_ASAP7_75t_L g5666 ( 
.A(n_3523),
.Y(n_5666)
);

NAND2xp5_ASAP7_75t_SL g5667 ( 
.A(n_3137),
.B(n_3266),
.Y(n_5667)
);

OAI22xp5_ASAP7_75t_SL g5668 ( 
.A1(n_3577),
.A2(n_3653),
.B1(n_3629),
.B2(n_3670),
.Y(n_5668)
);

INVx1_ASAP7_75t_SL g5669 ( 
.A(n_3303),
.Y(n_5669)
);

AOI221xp5_ASAP7_75t_L g5670 ( 
.A1(n_3587),
.A2(n_3690),
.B1(n_3578),
.B2(n_4057),
.C(n_4200),
.Y(n_5670)
);

INVx2_ASAP7_75t_SL g5671 ( 
.A(n_3137),
.Y(n_5671)
);

INVx1_ASAP7_75t_SL g5672 ( 
.A(n_3680),
.Y(n_5672)
);

INVx3_ASAP7_75t_L g5673 ( 
.A(n_3137),
.Y(n_5673)
);

AND3x1_ASAP7_75t_SL g5674 ( 
.A(n_3546),
.B(n_4333),
.C(n_3371),
.Y(n_5674)
);

NOR2xp33_ASAP7_75t_L g5675 ( 
.A(n_3638),
.B(n_3704),
.Y(n_5675)
);

INVx4_ASAP7_75t_L g5676 ( 
.A(n_3523),
.Y(n_5676)
);

AO22x1_ASAP7_75t_L g5677 ( 
.A1(n_3577),
.A2(n_3607),
.B1(n_3632),
.B2(n_3671),
.Y(n_5677)
);

AOI22xp5_ASAP7_75t_L g5678 ( 
.A1(n_4107),
.A2(n_4372),
.B1(n_4187),
.B2(n_3532),
.Y(n_5678)
);

INVxp67_ASAP7_75t_SL g5679 ( 
.A(n_3584),
.Y(n_5679)
);

INVx3_ASAP7_75t_L g5680 ( 
.A(n_3137),
.Y(n_5680)
);

AOI22xp5_ASAP7_75t_L g5681 ( 
.A1(n_3655),
.A2(n_3671),
.B1(n_3590),
.B2(n_3591),
.Y(n_5681)
);

CKINVDCx5p33_ASAP7_75t_R g5682 ( 
.A(n_4318),
.Y(n_5682)
);

AND3x1_ASAP7_75t_SL g5683 ( 
.A(n_4333),
.B(n_3371),
.C(n_3686),
.Y(n_5683)
);

CKINVDCx5p33_ASAP7_75t_R g5684 ( 
.A(n_4448),
.Y(n_5684)
);

INVx3_ASAP7_75t_L g5685 ( 
.A(n_3266),
.Y(n_5685)
);

INVx4_ASAP7_75t_L g5686 ( 
.A(n_3523),
.Y(n_5686)
);

BUFx12f_ASAP7_75t_L g5687 ( 
.A(n_3689),
.Y(n_5687)
);

AOI22xp33_ASAP7_75t_L g5688 ( 
.A1(n_3685),
.A2(n_3619),
.B1(n_3636),
.B2(n_3654),
.Y(n_5688)
);

OR2x6_ASAP7_75t_L g5689 ( 
.A(n_3584),
.B(n_3592),
.Y(n_5689)
);

BUFx2_ASAP7_75t_L g5690 ( 
.A(n_3618),
.Y(n_5690)
);

AOI22xp33_ASAP7_75t_L g5691 ( 
.A1(n_3685),
.A2(n_3636),
.B1(n_3654),
.B2(n_3662),
.Y(n_5691)
);

INVx2_ASAP7_75t_SL g5692 ( 
.A(n_3266),
.Y(n_5692)
);

BUFx4f_ASAP7_75t_L g5693 ( 
.A(n_3266),
.Y(n_5693)
);

AND3x1_ASAP7_75t_SL g5694 ( 
.A(n_3686),
.B(n_3688),
.C(n_4448),
.Y(n_5694)
);

NOR2xp33_ASAP7_75t_L g5695 ( 
.A(n_3638),
.B(n_3704),
.Y(n_5695)
);

BUFx2_ASAP7_75t_L g5696 ( 
.A(n_3618),
.Y(n_5696)
);

INVx3_ASAP7_75t_SL g5697 ( 
.A(n_4095),
.Y(n_5697)
);

A2O1A1Ixp33_ASAP7_75t_L g5698 ( 
.A1(n_3645),
.A2(n_3637),
.B(n_3643),
.C(n_3669),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_4448),
.Y(n_5699)
);

INVx4_ASAP7_75t_L g5700 ( 
.A(n_3523),
.Y(n_5700)
);

BUFx2_ASAP7_75t_L g5701 ( 
.A(n_3633),
.Y(n_5701)
);

BUFx6f_ASAP7_75t_L g5702 ( 
.A(n_3266),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_3646),
.B(n_3552),
.Y(n_5703)
);

INVx3_ASAP7_75t_L g5704 ( 
.A(n_3355),
.Y(n_5704)
);

BUFx3_ASAP7_75t_L g5705 ( 
.A(n_3632),
.Y(n_5705)
);

HB1xp67_ASAP7_75t_L g5706 ( 
.A(n_3355),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_L g5707 ( 
.A(n_3569),
.B(n_3571),
.Y(n_5707)
);

NAND2xp5_ASAP7_75t_L g5708 ( 
.A(n_3569),
.B(n_3571),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_3545),
.B(n_3551),
.Y(n_5709)
);

NAND2xp5_ASAP7_75t_L g5710 ( 
.A(n_3355),
.B(n_3429),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_SL g5711 ( 
.A(n_3355),
.B(n_3429),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_3613),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_3642),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_L g5714 ( 
.A(n_3355),
.B(n_3429),
.Y(n_5714)
);

INVx5_ASAP7_75t_L g5715 ( 
.A(n_3523),
.Y(n_5715)
);

BUFx10_ASAP7_75t_L g5716 ( 
.A(n_3237),
.Y(n_5716)
);

BUFx3_ASAP7_75t_L g5717 ( 
.A(n_3632),
.Y(n_5717)
);

INVxp67_ASAP7_75t_SL g5718 ( 
.A(n_3592),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_L g5719 ( 
.A(n_3355),
.B(n_3429),
.Y(n_5719)
);

AND2x6_ASAP7_75t_L g5720 ( 
.A(n_3237),
.B(n_3349),
.Y(n_5720)
);

O2A1O1Ixp33_ASAP7_75t_L g5721 ( 
.A1(n_3603),
.A2(n_3633),
.B(n_3644),
.C(n_3694),
.Y(n_5721)
);

NOR2xp33_ASAP7_75t_L g5722 ( 
.A(n_3704),
.B(n_3560),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_3659),
.Y(n_5723)
);

BUFx6f_ASAP7_75t_L g5724 ( 
.A(n_3429),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_3575),
.Y(n_5725)
);

INVx5_ASAP7_75t_L g5726 ( 
.A(n_3733),
.Y(n_5726)
);

A2O1A1Ixp33_ASAP7_75t_L g5727 ( 
.A1(n_4749),
.A2(n_3678),
.B(n_3627),
.C(n_3681),
.Y(n_5727)
);

INVxp67_ASAP7_75t_SL g5728 ( 
.A(n_5229),
.Y(n_5728)
);

BUFx6f_ASAP7_75t_L g5729 ( 
.A(n_4620),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_4488),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_SL g5731 ( 
.A(n_4514),
.B(n_3429),
.Y(n_5731)
);

INVx3_ASAP7_75t_L g5732 ( 
.A(n_5542),
.Y(n_5732)
);

OAI22xp5_ASAP7_75t_L g5733 ( 
.A1(n_4702),
.A2(n_3513),
.B1(n_3585),
.B2(n_3599),
.Y(n_5733)
);

OAI21xp5_ASAP7_75t_L g5734 ( 
.A1(n_4764),
.A2(n_3360),
.B(n_3426),
.Y(n_5734)
);

AND2x2_ASAP7_75t_SL g5735 ( 
.A(n_5061),
.B(n_3360),
.Y(n_5735)
);

AOI21xp5_ASAP7_75t_L g5736 ( 
.A1(n_5514),
.A2(n_3360),
.B(n_3426),
.Y(n_5736)
);

A2O1A1Ixp33_ASAP7_75t_L g5737 ( 
.A1(n_4749),
.A2(n_3580),
.B(n_3626),
.C(n_3676),
.Y(n_5737)
);

AOI21x1_ASAP7_75t_L g5738 ( 
.A1(n_4862),
.A2(n_3557),
.B(n_3508),
.Y(n_5738)
);

NOR2x1_ASAP7_75t_L g5739 ( 
.A(n_5186),
.B(n_3680),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5322),
.Y(n_5740)
);

BUFx2_ASAP7_75t_L g5741 ( 
.A(n_5460),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_5322),
.Y(n_5742)
);

NOR2xp33_ASAP7_75t_L g5743 ( 
.A(n_4828),
.B(n_3688),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_4504),
.B(n_3500),
.Y(n_5744)
);

O2A1O1Ixp33_ASAP7_75t_L g5745 ( 
.A1(n_4764),
.A2(n_3694),
.B(n_3644),
.C(n_3612),
.Y(n_5745)
);

AND2x4_ASAP7_75t_L g5746 ( 
.A(n_5175),
.B(n_3733),
.Y(n_5746)
);

OR2x2_ASAP7_75t_L g5747 ( 
.A(n_4757),
.B(n_3533),
.Y(n_5747)
);

BUFx3_ASAP7_75t_L g5748 ( 
.A(n_5460),
.Y(n_5748)
);

INVx1_ASAP7_75t_SL g5749 ( 
.A(n_4682),
.Y(n_5749)
);

AOI21xp5_ASAP7_75t_L g5750 ( 
.A1(n_5514),
.A2(n_3426),
.B(n_3360),
.Y(n_5750)
);

A2O1A1Ixp33_ASAP7_75t_L g5751 ( 
.A1(n_4933),
.A2(n_3676),
.B(n_3624),
.C(n_3582),
.Y(n_5751)
);

OR2x2_ASAP7_75t_L g5752 ( 
.A(n_4757),
.B(n_3680),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_4488),
.Y(n_5753)
);

AOI22xp33_ASAP7_75t_L g5754 ( 
.A1(n_4933),
.A2(n_3619),
.B1(n_3662),
.B2(n_3506),
.Y(n_5754)
);

OAI21xp33_ASAP7_75t_L g5755 ( 
.A1(n_4514),
.A2(n_3650),
.B(n_3660),
.Y(n_5755)
);

NAND2xp5_ASAP7_75t_L g5756 ( 
.A(n_4504),
.B(n_3500),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_4488),
.Y(n_5757)
);

AOI22xp33_ASAP7_75t_L g5758 ( 
.A1(n_4943),
.A2(n_3674),
.B1(n_3675),
.B2(n_3635),
.Y(n_5758)
);

BUFx6f_ASAP7_75t_L g5759 ( 
.A(n_4620),
.Y(n_5759)
);

INVx2_ASAP7_75t_L g5760 ( 
.A(n_4488),
.Y(n_5760)
);

INVx5_ASAP7_75t_L g5761 ( 
.A(n_4752),
.Y(n_5761)
);

OR2x6_ASAP7_75t_L g5762 ( 
.A(n_4480),
.B(n_4515),
.Y(n_5762)
);

OR2x6_ASAP7_75t_L g5763 ( 
.A(n_4480),
.B(n_3237),
.Y(n_5763)
);

INVx2_ASAP7_75t_SL g5764 ( 
.A(n_5460),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_L g5765 ( 
.A(n_4562),
.B(n_3500),
.Y(n_5765)
);

INVx3_ASAP7_75t_L g5766 ( 
.A(n_5542),
.Y(n_5766)
);

BUFx6f_ASAP7_75t_L g5767 ( 
.A(n_4620),
.Y(n_5767)
);

BUFx2_ASAP7_75t_L g5768 ( 
.A(n_5460),
.Y(n_5768)
);

NOR2xp33_ASAP7_75t_L g5769 ( 
.A(n_4828),
.B(n_3691),
.Y(n_5769)
);

NOR2xp33_ASAP7_75t_L g5770 ( 
.A(n_4820),
.B(n_3691),
.Y(n_5770)
);

INVx1_ASAP7_75t_SL g5771 ( 
.A(n_4682),
.Y(n_5771)
);

AOI22xp33_ASAP7_75t_L g5772 ( 
.A1(n_4943),
.A2(n_3674),
.B1(n_3675),
.B2(n_3593),
.Y(n_5772)
);

AND2x4_ASAP7_75t_L g5773 ( 
.A(n_5175),
.B(n_3733),
.Y(n_5773)
);

CKINVDCx5p33_ASAP7_75t_R g5774 ( 
.A(n_4558),
.Y(n_5774)
);

AND2x4_ASAP7_75t_L g5775 ( 
.A(n_5175),
.B(n_3733),
.Y(n_5775)
);

A2O1A1Ixp33_ASAP7_75t_L g5776 ( 
.A1(n_4582),
.A2(n_3595),
.B(n_3562),
.C(n_3594),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5322),
.Y(n_5777)
);

INVxp67_ASAP7_75t_L g5778 ( 
.A(n_5232),
.Y(n_5778)
);

AOI22xp33_ASAP7_75t_SL g5779 ( 
.A1(n_4582),
.A2(n_4625),
.B1(n_4993),
.B2(n_4977),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_4489),
.Y(n_5780)
);

AOI21xp5_ASAP7_75t_L g5781 ( 
.A1(n_5528),
.A2(n_3426),
.B(n_3494),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5322),
.Y(n_5782)
);

INVx2_ASAP7_75t_L g5783 ( 
.A(n_4492),
.Y(n_5783)
);

BUFx2_ASAP7_75t_L g5784 ( 
.A(n_5460),
.Y(n_5784)
);

OAI22xp5_ASAP7_75t_L g5785 ( 
.A1(n_4702),
.A2(n_3616),
.B1(n_3560),
.B2(n_3585),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5327),
.Y(n_5786)
);

NOR2xp33_ASAP7_75t_L g5787 ( 
.A(n_4820),
.B(n_3691),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5327),
.Y(n_5788)
);

A2O1A1Ixp33_ASAP7_75t_L g5789 ( 
.A1(n_4625),
.A2(n_3606),
.B(n_3567),
.C(n_3572),
.Y(n_5789)
);

NAND2xp5_ASAP7_75t_SL g5790 ( 
.A(n_4594),
.B(n_3500),
.Y(n_5790)
);

AOI21xp5_ASAP7_75t_L g5791 ( 
.A1(n_5528),
.A2(n_3510),
.B(n_3550),
.Y(n_5791)
);

AOI21xp5_ASAP7_75t_L g5792 ( 
.A1(n_4544),
.A2(n_3539),
.B(n_3733),
.Y(n_5792)
);

NAND2xp5_ASAP7_75t_L g5793 ( 
.A(n_4562),
.B(n_3500),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_4492),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_4494),
.Y(n_5795)
);

NOR2xp33_ASAP7_75t_L g5796 ( 
.A(n_4479),
.B(n_3560),
.Y(n_5796)
);

OAI22xp5_ASAP7_75t_SL g5797 ( 
.A1(n_5129),
.A2(n_4993),
.B1(n_4977),
.B2(n_4589),
.Y(n_5797)
);

INVx2_ASAP7_75t_L g5798 ( 
.A(n_4494),
.Y(n_5798)
);

BUFx3_ASAP7_75t_L g5799 ( 
.A(n_4616),
.Y(n_5799)
);

NOR2x1_ASAP7_75t_SL g5800 ( 
.A(n_4968),
.B(n_3733),
.Y(n_5800)
);

INVxp67_ASAP7_75t_SL g5801 ( 
.A(n_5229),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5327),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5327),
.Y(n_5803)
);

AOI21xp5_ASAP7_75t_L g5804 ( 
.A1(n_4544),
.A2(n_3500),
.B(n_3547),
.Y(n_5804)
);

INVx2_ASAP7_75t_SL g5805 ( 
.A(n_5175),
.Y(n_5805)
);

INVx3_ASAP7_75t_L g5806 ( 
.A(n_5542),
.Y(n_5806)
);

OAI22xp5_ASAP7_75t_L g5807 ( 
.A1(n_4716),
.A2(n_3585),
.B1(n_3616),
.B2(n_3560),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5338),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5338),
.Y(n_5809)
);

OAI22xp5_ASAP7_75t_L g5810 ( 
.A1(n_4716),
.A2(n_3585),
.B1(n_3599),
.B2(n_3616),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_4564),
.B(n_4584),
.Y(n_5811)
);

OAI22xp5_ASAP7_75t_L g5812 ( 
.A1(n_4740),
.A2(n_4795),
.B1(n_4589),
.B2(n_4630),
.Y(n_5812)
);

BUFx2_ASAP7_75t_L g5813 ( 
.A(n_4610),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_4494),
.Y(n_5814)
);

INVx1_ASAP7_75t_SL g5815 ( 
.A(n_4714),
.Y(n_5815)
);

OR2x6_ASAP7_75t_L g5816 ( 
.A(n_4480),
.B(n_4515),
.Y(n_5816)
);

HB1xp67_ASAP7_75t_L g5817 ( 
.A(n_4531),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_4497),
.Y(n_5818)
);

NAND2xp5_ASAP7_75t_L g5819 ( 
.A(n_4564),
.B(n_3547),
.Y(n_5819)
);

INVx2_ASAP7_75t_L g5820 ( 
.A(n_4497),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5338),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5338),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5339),
.Y(n_5823)
);

AOI22xp33_ASAP7_75t_L g5824 ( 
.A1(n_4903),
.A2(n_3593),
.B1(n_3519),
.B2(n_3689),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_4497),
.Y(n_5825)
);

BUFx3_ASAP7_75t_L g5826 ( 
.A(n_4616),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_L g5827 ( 
.A(n_4584),
.B(n_3547),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5339),
.Y(n_5828)
);

NOR2xp33_ASAP7_75t_L g5829 ( 
.A(n_4479),
.B(n_3599),
.Y(n_5829)
);

NAND2xp5_ASAP7_75t_L g5830 ( 
.A(n_4617),
.B(n_4785),
.Y(n_5830)
);

O2A1O1Ixp5_ASAP7_75t_L g5831 ( 
.A1(n_4477),
.A2(n_3220),
.B(n_3354),
.C(n_3424),
.Y(n_5831)
);

NOR2xp33_ASAP7_75t_L g5832 ( 
.A(n_4801),
.B(n_3599),
.Y(n_5832)
);

INVxp67_ASAP7_75t_L g5833 ( 
.A(n_5232),
.Y(n_5833)
);

NAND2xp5_ASAP7_75t_L g5834 ( 
.A(n_4617),
.B(n_3220),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_4785),
.B(n_3220),
.Y(n_5835)
);

BUFx3_ASAP7_75t_L g5836 ( 
.A(n_4616),
.Y(n_5836)
);

AND2x2_ASAP7_75t_SL g5837 ( 
.A(n_5061),
.B(n_3237),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5339),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5339),
.Y(n_5839)
);

INVx3_ASAP7_75t_L g5840 ( 
.A(n_5542),
.Y(n_5840)
);

BUFx2_ASAP7_75t_SL g5841 ( 
.A(n_5180),
.Y(n_5841)
);

NAND2xp5_ASAP7_75t_L g5842 ( 
.A(n_4802),
.B(n_3220),
.Y(n_5842)
);

A2O1A1Ixp33_ASAP7_75t_L g5843 ( 
.A1(n_4594),
.A2(n_3696),
.B(n_3692),
.C(n_3701),
.Y(n_5843)
);

AND2x2_ASAP7_75t_L g5844 ( 
.A(n_4680),
.B(n_3616),
.Y(n_5844)
);

AOI22xp5_ASAP7_75t_L g5845 ( 
.A1(n_4885),
.A2(n_3593),
.B1(n_3519),
.B2(n_3702),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5344),
.Y(n_5846)
);

BUFx2_ASAP7_75t_L g5847 ( 
.A(n_4610),
.Y(n_5847)
);

AOI22xp33_ASAP7_75t_L g5848 ( 
.A1(n_4903),
.A2(n_3519),
.B1(n_3689),
.B2(n_3615),
.Y(n_5848)
);

NAND2xp5_ASAP7_75t_L g5849 ( 
.A(n_4802),
.B(n_3354),
.Y(n_5849)
);

OAI22xp5_ASAP7_75t_L g5850 ( 
.A1(n_4740),
.A2(n_3677),
.B1(n_3650),
.B2(n_3706),
.Y(n_5850)
);

BUFx12f_ASAP7_75t_L g5851 ( 
.A(n_4609),
.Y(n_5851)
);

HB1xp67_ASAP7_75t_L g5852 ( 
.A(n_4531),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5344),
.Y(n_5853)
);

OAI22xp5_ASAP7_75t_L g5854 ( 
.A1(n_4795),
.A2(n_3677),
.B1(n_3706),
.B2(n_3700),
.Y(n_5854)
);

AOI21xp5_ASAP7_75t_L g5855 ( 
.A1(n_4719),
.A2(n_3601),
.B(n_3354),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_SL g5856 ( 
.A(n_4630),
.B(n_3424),
.Y(n_5856)
);

BUFx2_ASAP7_75t_L g5857 ( 
.A(n_4610),
.Y(n_5857)
);

O2A1O1Ixp33_ASAP7_75t_L g5858 ( 
.A1(n_4761),
.A2(n_4632),
.B(n_4597),
.C(n_4539),
.Y(n_5858)
);

BUFx12f_ASAP7_75t_L g5859 ( 
.A(n_4609),
.Y(n_5859)
);

A2O1A1Ixp33_ASAP7_75t_L g5860 ( 
.A1(n_4493),
.A2(n_3600),
.B(n_3695),
.C(n_3679),
.Y(n_5860)
);

NAND2xp5_ASAP7_75t_SL g5861 ( 
.A(n_4655),
.B(n_3424),
.Y(n_5861)
);

AOI221xp5_ASAP7_75t_L g5862 ( 
.A1(n_4542),
.A2(n_3709),
.B1(n_3683),
.B2(n_3693),
.C(n_3684),
.Y(n_5862)
);

NOR2xp33_ASAP7_75t_L g5863 ( 
.A(n_4801),
.B(n_3700),
.Y(n_5863)
);

NAND2xp5_ASAP7_75t_L g5864 ( 
.A(n_4835),
.B(n_3354),
.Y(n_5864)
);

BUFx12f_ASAP7_75t_L g5865 ( 
.A(n_4641),
.Y(n_5865)
);

CKINVDCx8_ASAP7_75t_R g5866 ( 
.A(n_5333),
.Y(n_5866)
);

NAND2xp5_ASAP7_75t_L g5867 ( 
.A(n_4835),
.B(n_3424),
.Y(n_5867)
);

NAND2xp5_ASAP7_75t_L g5868 ( 
.A(n_4907),
.B(n_3538),
.Y(n_5868)
);

INVx2_ASAP7_75t_SL g5869 ( 
.A(n_5180),
.Y(n_5869)
);

A2O1A1Ixp33_ASAP7_75t_L g5870 ( 
.A1(n_4493),
.A2(n_3600),
.B(n_3667),
.C(n_3666),
.Y(n_5870)
);

O2A1O1Ixp5_ASAP7_75t_L g5871 ( 
.A1(n_4477),
.A2(n_3625),
.B(n_3609),
.C(n_3687),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_L g5872 ( 
.A(n_4907),
.B(n_3538),
.Y(n_5872)
);

NOR2xp33_ASAP7_75t_L g5873 ( 
.A(n_4858),
.B(n_3557),
.Y(n_5873)
);

OAI22xp5_ASAP7_75t_L g5874 ( 
.A1(n_4696),
.A2(n_3677),
.B1(n_3706),
.B2(n_3639),
.Y(n_5874)
);

AOI21xp5_ASAP7_75t_L g5875 ( 
.A1(n_4719),
.A2(n_3486),
.B(n_3385),
.Y(n_5875)
);

BUFx12f_ASAP7_75t_L g5876 ( 
.A(n_4641),
.Y(n_5876)
);

AOI21xp5_ASAP7_75t_L g5877 ( 
.A1(n_4855),
.A2(n_3486),
.B(n_3385),
.Y(n_5877)
);

INVx2_ASAP7_75t_SL g5878 ( 
.A(n_5180),
.Y(n_5878)
);

AND2x4_ASAP7_75t_L g5879 ( 
.A(n_5180),
.B(n_3349),
.Y(n_5879)
);

AOI21xp5_ASAP7_75t_L g5880 ( 
.A1(n_4855),
.A2(n_3292),
.B(n_3385),
.Y(n_5880)
);

NOR2xp33_ASAP7_75t_L g5881 ( 
.A(n_4858),
.B(n_4867),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5344),
.Y(n_5882)
);

NOR2xp33_ASAP7_75t_L g5883 ( 
.A(n_4867),
.B(n_3703),
.Y(n_5883)
);

O2A1O1Ixp33_ASAP7_75t_L g5884 ( 
.A1(n_4761),
.A2(n_3699),
.B(n_3631),
.C(n_3549),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5344),
.Y(n_5885)
);

OAI22xp5_ASAP7_75t_L g5886 ( 
.A1(n_4696),
.A2(n_3677),
.B1(n_3706),
.B2(n_3292),
.Y(n_5886)
);

INVx2_ASAP7_75t_SL g5887 ( 
.A(n_5180),
.Y(n_5887)
);

NAND2xp5_ASAP7_75t_SL g5888 ( 
.A(n_4655),
.B(n_4781),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_SL g5889 ( 
.A(n_4655),
.B(n_3687),
.Y(n_5889)
);

NOR2xp33_ASAP7_75t_L g5890 ( 
.A(n_4999),
.B(n_3703),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5355),
.Y(n_5891)
);

NOR2x1_ASAP7_75t_SL g5892 ( 
.A(n_4968),
.B(n_3684),
.Y(n_5892)
);

INVx4_ASAP7_75t_SL g5893 ( 
.A(n_5207),
.Y(n_5893)
);

O2A1O1Ixp33_ASAP7_75t_L g5894 ( 
.A1(n_4597),
.A2(n_4632),
.B(n_4677),
.C(n_4539),
.Y(n_5894)
);

A2O1A1Ixp33_ASAP7_75t_SL g5895 ( 
.A1(n_5384),
.A2(n_3621),
.B(n_3610),
.C(n_3581),
.Y(n_5895)
);

AND2x2_ASAP7_75t_L g5896 ( 
.A(n_4680),
.B(n_3292),
.Y(n_5896)
);

AOI22xp33_ASAP7_75t_L g5897 ( 
.A1(n_4723),
.A2(n_3689),
.B1(n_3615),
.B2(n_3665),
.Y(n_5897)
);

OAI21xp5_ASAP7_75t_L g5898 ( 
.A1(n_4677),
.A2(n_3698),
.B(n_3697),
.Y(n_5898)
);

NAND2xp5_ASAP7_75t_L g5899 ( 
.A(n_4931),
.B(n_3622),
.Y(n_5899)
);

AOI22xp33_ASAP7_75t_L g5900 ( 
.A1(n_4723),
.A2(n_4542),
.B1(n_4914),
.B2(n_4755),
.Y(n_5900)
);

O2A1O1Ixp33_ASAP7_75t_L g5901 ( 
.A1(n_4726),
.A2(n_4746),
.B(n_4777),
.C(n_4948),
.Y(n_5901)
);

A2O1A1Ixp33_ASAP7_75t_L g5902 ( 
.A1(n_4554),
.A2(n_3672),
.B(n_3349),
.C(n_3693),
.Y(n_5902)
);

BUFx2_ASAP7_75t_L g5903 ( 
.A(n_4642),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_4931),
.B(n_3611),
.Y(n_5904)
);

INVx1_ASAP7_75t_SL g5905 ( 
.A(n_4714),
.Y(n_5905)
);

NAND2xp5_ASAP7_75t_L g5906 ( 
.A(n_4984),
.B(n_3611),
.Y(n_5906)
);

AOI21xp5_ASAP7_75t_L g5907 ( 
.A1(n_4963),
.A2(n_5090),
.B(n_4990),
.Y(n_5907)
);

NOR2xp33_ASAP7_75t_L g5908 ( 
.A(n_4999),
.B(n_3656),
.Y(n_5908)
);

BUFx2_ASAP7_75t_L g5909 ( 
.A(n_4642),
.Y(n_5909)
);

BUFx2_ASAP7_75t_L g5910 ( 
.A(n_4642),
.Y(n_5910)
);

NAND2xp5_ASAP7_75t_SL g5911 ( 
.A(n_4781),
.B(n_3349),
.Y(n_5911)
);

OAI22xp33_ASAP7_75t_L g5912 ( 
.A1(n_4941),
.A2(n_3537),
.B1(n_3707),
.B2(n_3665),
.Y(n_5912)
);

A2O1A1Ixp33_ASAP7_75t_L g5913 ( 
.A1(n_4554),
.A2(n_3707),
.B(n_3658),
.C(n_3661),
.Y(n_5913)
);

AOI221x1_ASAP7_75t_L g5914 ( 
.A1(n_4726),
.A2(n_3605),
.B1(n_3661),
.B2(n_3652),
.C(n_3651),
.Y(n_5914)
);

BUFx3_ASAP7_75t_L g5915 ( 
.A(n_4616),
.Y(n_5915)
);

BUFx12f_ASAP7_75t_L g5916 ( 
.A(n_4667),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5355),
.Y(n_5917)
);

INVx1_ASAP7_75t_SL g5918 ( 
.A(n_4613),
.Y(n_5918)
);

INVxp67_ASAP7_75t_SL g5919 ( 
.A(n_5044),
.Y(n_5919)
);

NAND2xp5_ASAP7_75t_SL g5920 ( 
.A(n_4797),
.B(n_3537),
.Y(n_5920)
);

AOI22xp33_ASAP7_75t_SL g5921 ( 
.A1(n_5213),
.A2(n_3663),
.B1(n_3604),
.B2(n_3605),
.Y(n_5921)
);

NOR2xp33_ASAP7_75t_R g5922 ( 
.A(n_4751),
.B(n_3623),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5355),
.Y(n_5923)
);

HAxp5_ASAP7_75t_L g5924 ( 
.A(n_5129),
.B(n_3488),
.CON(n_5924),
.SN(n_5924)
);

NAND2xp5_ASAP7_75t_SL g5925 ( 
.A(n_4797),
.B(n_3537),
.Y(n_5925)
);

BUFx8_ASAP7_75t_SL g5926 ( 
.A(n_4558),
.Y(n_5926)
);

NAND2xp5_ASAP7_75t_SL g5927 ( 
.A(n_4746),
.B(n_3604),
.Y(n_5927)
);

CKINVDCx20_ASAP7_75t_R g5928 ( 
.A(n_4637),
.Y(n_5928)
);

NOR2xp33_ASAP7_75t_L g5929 ( 
.A(n_4948),
.B(n_3663),
.Y(n_5929)
);

A2O1A1Ixp33_ASAP7_75t_L g5930 ( 
.A1(n_4635),
.A2(n_3597),
.B(n_3651),
.C(n_3576),
.Y(n_5930)
);

HB1xp67_ASAP7_75t_L g5931 ( 
.A(n_4568),
.Y(n_5931)
);

INVx1_ASAP7_75t_SL g5932 ( 
.A(n_4613),
.Y(n_5932)
);

OR2x6_ASAP7_75t_L g5933 ( 
.A(n_4480),
.B(n_3597),
.Y(n_5933)
);

OAI21xp5_ASAP7_75t_L g5934 ( 
.A1(n_4777),
.A2(n_3541),
.B(n_3570),
.Y(n_5934)
);

INVx2_ASAP7_75t_SL g5935 ( 
.A(n_5180),
.Y(n_5935)
);

AOI21xp5_ASAP7_75t_L g5936 ( 
.A1(n_4963),
.A2(n_3576),
.B(n_3579),
.Y(n_5936)
);

O2A1O1Ixp33_ASAP7_75t_L g5937 ( 
.A1(n_4481),
.A2(n_3579),
.B(n_3652),
.C(n_3589),
.Y(n_5937)
);

AND2x2_ASAP7_75t_SL g5938 ( 
.A(n_5061),
.B(n_3622),
.Y(n_5938)
);

INVx1_ASAP7_75t_SL g5939 ( 
.A(n_4659),
.Y(n_5939)
);

AOI21xp5_ASAP7_75t_L g5940 ( 
.A1(n_4990),
.A2(n_3589),
.B(n_3596),
.Y(n_5940)
);

A2O1A1Ixp33_ASAP7_75t_SL g5941 ( 
.A1(n_5384),
.A2(n_3583),
.B(n_3608),
.C(n_3596),
.Y(n_5941)
);

AOI222xp33_ASAP7_75t_L g5942 ( 
.A1(n_4914),
.A2(n_3630),
.B1(n_3640),
.B2(n_3649),
.C1(n_4755),
.C2(n_4519),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5355),
.Y(n_5943)
);

AOI22xp33_ASAP7_75t_L g5944 ( 
.A1(n_4921),
.A2(n_3630),
.B1(n_3640),
.B2(n_3649),
.Y(n_5944)
);

A2O1A1Ixp33_ASAP7_75t_L g5945 ( 
.A1(n_4635),
.A2(n_4647),
.B(n_5419),
.C(n_5025),
.Y(n_5945)
);

A2O1A1Ixp33_ASAP7_75t_L g5946 ( 
.A1(n_4647),
.A2(n_5419),
.B(n_5025),
.C(n_5091),
.Y(n_5946)
);

CKINVDCx11_ASAP7_75t_R g5947 ( 
.A(n_4637),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5358),
.Y(n_5948)
);

INVxp67_ASAP7_75t_SL g5949 ( 
.A(n_5044),
.Y(n_5949)
);

AOI22xp5_ASAP7_75t_L g5950 ( 
.A1(n_4885),
.A2(n_4946),
.B1(n_4902),
.B2(n_4941),
.Y(n_5950)
);

AOI221xp5_ASAP7_75t_L g5951 ( 
.A1(n_5213),
.A2(n_5316),
.B1(n_4651),
.B2(n_4634),
.C(n_4672),
.Y(n_5951)
);

O2A1O1Ixp33_ASAP7_75t_L g5952 ( 
.A1(n_4481),
.A2(n_4519),
.B(n_4566),
.C(n_4533),
.Y(n_5952)
);

AOI21xp5_ASAP7_75t_L g5953 ( 
.A1(n_5090),
.A2(n_5376),
.B(n_5131),
.Y(n_5953)
);

NAND2xp5_ASAP7_75t_SL g5954 ( 
.A(n_4527),
.B(n_4538),
.Y(n_5954)
);

AND2x6_ASAP7_75t_L g5955 ( 
.A(n_5555),
.B(n_5558),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5442),
.Y(n_5956)
);

INVx2_ASAP7_75t_SL g5957 ( 
.A(n_5180),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5358),
.Y(n_5958)
);

OAI21xp33_ASAP7_75t_SL g5959 ( 
.A1(n_4533),
.A2(n_4596),
.B(n_4566),
.Y(n_5959)
);

A2O1A1Ixp33_ASAP7_75t_L g5960 ( 
.A1(n_5080),
.A2(n_5096),
.B(n_5091),
.C(n_5163),
.Y(n_5960)
);

CKINVDCx5p33_ASAP7_75t_R g5961 ( 
.A(n_4685),
.Y(n_5961)
);

O2A1O1Ixp33_ASAP7_75t_L g5962 ( 
.A1(n_4596),
.A2(n_4623),
.B(n_5151),
.C(n_5121),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5358),
.Y(n_5963)
);

AOI21xp5_ASAP7_75t_L g5964 ( 
.A1(n_5131),
.A2(n_5433),
.B(n_5376),
.Y(n_5964)
);

AOI21xp5_ASAP7_75t_L g5965 ( 
.A1(n_5433),
.A2(n_5445),
.B(n_5519),
.Y(n_5965)
);

INVx2_ASAP7_75t_L g5966 ( 
.A(n_5442),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5358),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5363),
.Y(n_5968)
);

AOI21xp5_ASAP7_75t_L g5969 ( 
.A1(n_5445),
.A2(n_5525),
.B(n_5519),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5363),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5363),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5442),
.Y(n_5972)
);

AOI21xp5_ASAP7_75t_L g5973 ( 
.A1(n_5525),
.A2(n_5536),
.B(n_5520),
.Y(n_5973)
);

O2A1O1Ixp33_ASAP7_75t_L g5974 ( 
.A1(n_4623),
.A2(n_5151),
.B(n_5121),
.C(n_5080),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_4685),
.Y(n_5975)
);

BUFx3_ASAP7_75t_L g5976 ( 
.A(n_4616),
.Y(n_5976)
);

NOR2xp33_ASAP7_75t_SL g5977 ( 
.A(n_5397),
.B(n_5474),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_5442),
.Y(n_5978)
);

INVxp67_ASAP7_75t_SL g5979 ( 
.A(n_4949),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5363),
.Y(n_5980)
);

NAND2xp5_ASAP7_75t_SL g5981 ( 
.A(n_4527),
.B(n_4538),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5377),
.Y(n_5982)
);

AOI22xp5_ASAP7_75t_L g5983 ( 
.A1(n_4902),
.A2(n_4946),
.B1(n_5010),
.B2(n_4942),
.Y(n_5983)
);

OAI22xp5_ASAP7_75t_L g5984 ( 
.A1(n_4541),
.A2(n_4549),
.B1(n_4555),
.B2(n_4548),
.Y(n_5984)
);

AOI21xp33_ASAP7_75t_L g5985 ( 
.A1(n_4690),
.A2(n_4721),
.B(n_5217),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5377),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5377),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5377),
.Y(n_5988)
);

AND2x4_ASAP7_75t_L g5989 ( 
.A(n_5241),
.B(n_5333),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_4984),
.B(n_5074),
.Y(n_5990)
);

OR2x6_ASAP7_75t_L g5991 ( 
.A(n_4480),
.B(n_4515),
.Y(n_5991)
);

INVx2_ASAP7_75t_L g5992 ( 
.A(n_5461),
.Y(n_5992)
);

INVxp67_ASAP7_75t_L g5993 ( 
.A(n_5238),
.Y(n_5993)
);

CKINVDCx20_ASAP7_75t_R g5994 ( 
.A(n_4684),
.Y(n_5994)
);

AOI22xp33_ASAP7_75t_SL g5995 ( 
.A1(n_5328),
.A2(n_5163),
.B1(n_4563),
.B2(n_4548),
.Y(n_5995)
);

INVx2_ASAP7_75t_L g5996 ( 
.A(n_5461),
.Y(n_5996)
);

AOI22xp5_ASAP7_75t_L g5997 ( 
.A1(n_4942),
.A2(n_5105),
.B1(n_5010),
.B2(n_4577),
.Y(n_5997)
);

INVx6_ASAP7_75t_L g5998 ( 
.A(n_5333),
.Y(n_5998)
);

AOI22xp33_ASAP7_75t_L g5999 ( 
.A1(n_4921),
.A2(n_4672),
.B1(n_5106),
.B2(n_5096),
.Y(n_5999)
);

AOI22xp33_ASAP7_75t_L g6000 ( 
.A1(n_5106),
.A2(n_4967),
.B1(n_4937),
.B2(n_4651),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5382),
.Y(n_6001)
);

AND2x4_ASAP7_75t_L g6002 ( 
.A(n_5241),
.B(n_5333),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5382),
.Y(n_6003)
);

INVx2_ASAP7_75t_L g6004 ( 
.A(n_5461),
.Y(n_6004)
);

HB1xp67_ASAP7_75t_L g6005 ( 
.A(n_4568),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5641),
.Y(n_6006)
);

INVx6_ASAP7_75t_L g6007 ( 
.A(n_5333),
.Y(n_6007)
);

NAND2xp5_ASAP7_75t_L g6008 ( 
.A(n_5074),
.B(n_5092),
.Y(n_6008)
);

BUFx2_ASAP7_75t_L g6009 ( 
.A(n_4502),
.Y(n_6009)
);

AOI21xp33_ASAP7_75t_L g6010 ( 
.A1(n_4690),
.A2(n_4721),
.B(n_5217),
.Y(n_6010)
);

AOI21xp5_ASAP7_75t_L g6011 ( 
.A1(n_5536),
.A2(n_5520),
.B(n_5346),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_4703),
.B(n_4733),
.Y(n_6012)
);

NOR2xp33_ASAP7_75t_L g6013 ( 
.A(n_4843),
.B(n_4845),
.Y(n_6013)
);

NAND2xp5_ASAP7_75t_L g6014 ( 
.A(n_5092),
.B(n_5100),
.Y(n_6014)
);

NOR2xp33_ASAP7_75t_L g6015 ( 
.A(n_4843),
.B(n_4845),
.Y(n_6015)
);

OAI22xp5_ASAP7_75t_L g6016 ( 
.A1(n_4541),
.A2(n_4555),
.B1(n_4560),
.B2(n_4549),
.Y(n_6016)
);

BUFx3_ASAP7_75t_L g6017 ( 
.A(n_4799),
.Y(n_6017)
);

NAND2xp5_ASAP7_75t_L g6018 ( 
.A(n_5100),
.B(n_4648),
.Y(n_6018)
);

NAND2x1p5_ASAP7_75t_L g6019 ( 
.A(n_4524),
.B(n_4511),
.Y(n_6019)
);

CKINVDCx8_ASAP7_75t_R g6020 ( 
.A(n_5333),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5461),
.Y(n_6021)
);

O2A1O1Ixp33_ASAP7_75t_L g6022 ( 
.A1(n_5117),
.A2(n_5057),
.B(n_4563),
.C(n_4565),
.Y(n_6022)
);

AOI22xp33_ASAP7_75t_L g6023 ( 
.A1(n_4937),
.A2(n_4967),
.B1(n_4634),
.B2(n_4986),
.Y(n_6023)
);

OAI22xp5_ASAP7_75t_L g6024 ( 
.A1(n_4560),
.A2(n_4569),
.B1(n_4574),
.B2(n_4565),
.Y(n_6024)
);

O2A1O1Ixp33_ASAP7_75t_L g6025 ( 
.A1(n_5117),
.A2(n_5057),
.B(n_4574),
.C(n_4585),
.Y(n_6025)
);

AOI21xp5_ASAP7_75t_L g6026 ( 
.A1(n_5337),
.A2(n_5347),
.B(n_5346),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5382),
.Y(n_6027)
);

NOR2xp33_ASAP7_75t_L g6028 ( 
.A(n_4847),
.B(n_4851),
.Y(n_6028)
);

A2O1A1Ixp33_ASAP7_75t_SL g6029 ( 
.A1(n_5387),
.A2(n_5218),
.B(n_5059),
.C(n_5119),
.Y(n_6029)
);

INVx6_ASAP7_75t_L g6030 ( 
.A(n_5333),
.Y(n_6030)
);

NAND2xp5_ASAP7_75t_L g6031 ( 
.A(n_4648),
.B(n_4687),
.Y(n_6031)
);

INVx6_ASAP7_75t_L g6032 ( 
.A(n_5241),
.Y(n_6032)
);

INVx6_ASAP7_75t_SL g6033 ( 
.A(n_4698),
.Y(n_6033)
);

OAI21x1_ASAP7_75t_SL g6034 ( 
.A1(n_4569),
.A2(n_4591),
.B(n_4585),
.Y(n_6034)
);

AND2x2_ASAP7_75t_L g6035 ( 
.A(n_4703),
.B(n_4733),
.Y(n_6035)
);

AOI21xp5_ASAP7_75t_L g6036 ( 
.A1(n_5337),
.A2(n_5424),
.B(n_5347),
.Y(n_6036)
);

OR2x2_ASAP7_75t_L g6037 ( 
.A(n_4670),
.B(n_4681),
.Y(n_6037)
);

AND2x4_ASAP7_75t_L g6038 ( 
.A(n_5241),
.B(n_5356),
.Y(n_6038)
);

HB1xp67_ASAP7_75t_L g6039 ( 
.A(n_4580),
.Y(n_6039)
);

HB1xp67_ASAP7_75t_L g6040 ( 
.A(n_4580),
.Y(n_6040)
);

INVx3_ASAP7_75t_L g6041 ( 
.A(n_5641),
.Y(n_6041)
);

AOI221xp5_ASAP7_75t_L g6042 ( 
.A1(n_5316),
.A2(n_5370),
.B1(n_5491),
.B2(n_5492),
.C(n_5185),
.Y(n_6042)
);

AO21x2_ASAP7_75t_L g6043 ( 
.A1(n_4717),
.A2(n_4789),
.B(n_4775),
.Y(n_6043)
);

AND2x2_ASAP7_75t_L g6044 ( 
.A(n_5412),
.B(n_5415),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5382),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_SL g6046 ( 
.A(n_4591),
.B(n_4593),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5391),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5391),
.Y(n_6048)
);

NOR2xp33_ASAP7_75t_L g6049 ( 
.A(n_4847),
.B(n_4851),
.Y(n_6049)
);

NAND2xp5_ASAP7_75t_L g6050 ( 
.A(n_4687),
.B(n_4693),
.Y(n_6050)
);

NOR2xp33_ASAP7_75t_L g6051 ( 
.A(n_4853),
.B(n_4856),
.Y(n_6051)
);

AOI21xp5_ASAP7_75t_L g6052 ( 
.A1(n_5424),
.A2(n_5540),
.B(n_5427),
.Y(n_6052)
);

AOI22xp33_ASAP7_75t_SL g6053 ( 
.A1(n_5328),
.A2(n_4600),
.B1(n_4602),
.B2(n_4593),
.Y(n_6053)
);

O2A1O1Ixp33_ASAP7_75t_SL g6054 ( 
.A1(n_4600),
.A2(n_4602),
.B(n_4611),
.C(n_4603),
.Y(n_6054)
);

AND2x4_ASAP7_75t_L g6055 ( 
.A(n_5241),
.B(n_5356),
.Y(n_6055)
);

NAND2xp5_ASAP7_75t_L g6056 ( 
.A(n_4693),
.B(n_4709),
.Y(n_6056)
);

BUFx6f_ASAP7_75t_SL g6057 ( 
.A(n_5397),
.Y(n_6057)
);

INVx4_ASAP7_75t_L g6058 ( 
.A(n_4511),
.Y(n_6058)
);

CKINVDCx20_ASAP7_75t_R g6059 ( 
.A(n_4684),
.Y(n_6059)
);

AOI21xp5_ASAP7_75t_L g6060 ( 
.A1(n_5427),
.A2(n_5552),
.B(n_5540),
.Y(n_6060)
);

AOI21xp5_ASAP7_75t_L g6061 ( 
.A1(n_5552),
.A2(n_5571),
.B(n_5566),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_SL g6062 ( 
.A(n_4603),
.B(n_4611),
.Y(n_6062)
);

INVx1_ASAP7_75t_SL g6063 ( 
.A(n_4659),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5391),
.Y(n_6064)
);

A2O1A1Ixp33_ASAP7_75t_L g6065 ( 
.A1(n_5218),
.A2(n_5541),
.B(n_4966),
.C(n_4636),
.Y(n_6065)
);

BUFx4f_ASAP7_75t_L g6066 ( 
.A(n_4524),
.Y(n_6066)
);

AOI21xp5_ASAP7_75t_L g6067 ( 
.A1(n_5566),
.A2(n_5571),
.B(n_4929),
.Y(n_6067)
);

BUFx2_ASAP7_75t_SL g6068 ( 
.A(n_5587),
.Y(n_6068)
);

AOI22xp5_ASAP7_75t_L g6069 ( 
.A1(n_5105),
.A2(n_4577),
.B1(n_5047),
.B2(n_4986),
.Y(n_6069)
);

HB1xp67_ASAP7_75t_L g6070 ( 
.A(n_4709),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_SL g6071 ( 
.A(n_4612),
.B(n_4619),
.Y(n_6071)
);

AND2x4_ASAP7_75t_L g6072 ( 
.A(n_5356),
.B(n_5398),
.Y(n_6072)
);

AOI21xp5_ASAP7_75t_L g6073 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6073)
);

NAND2x1p5_ASAP7_75t_L g6074 ( 
.A(n_4524),
.B(n_4511),
.Y(n_6074)
);

INVx2_ASAP7_75t_SL g6075 ( 
.A(n_5597),
.Y(n_6075)
);

NAND2xp5_ASAP7_75t_L g6076 ( 
.A(n_4873),
.B(n_4874),
.Y(n_6076)
);

O2A1O1Ixp33_ASAP7_75t_L g6077 ( 
.A1(n_4612),
.A2(n_4619),
.B(n_5492),
.C(n_5491),
.Y(n_6077)
);

OAI22xp5_ASAP7_75t_L g6078 ( 
.A1(n_4853),
.A2(n_4865),
.B1(n_4883),
.B2(n_4856),
.Y(n_6078)
);

NAND2xp5_ASAP7_75t_L g6079 ( 
.A(n_4873),
.B(n_4874),
.Y(n_6079)
);

AOI22xp33_ASAP7_75t_L g6080 ( 
.A1(n_5047),
.A2(n_5069),
.B1(n_5541),
.B2(n_5185),
.Y(n_6080)
);

AND2x4_ASAP7_75t_L g6081 ( 
.A(n_5356),
.B(n_5398),
.Y(n_6081)
);

BUFx12f_ASAP7_75t_L g6082 ( 
.A(n_4667),
.Y(n_6082)
);

AND2x4_ASAP7_75t_L g6083 ( 
.A(n_5398),
.B(n_5478),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5391),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_SL g6085 ( 
.A(n_5059),
.B(n_5115),
.Y(n_6085)
);

AOI222xp33_ASAP7_75t_L g6086 ( 
.A1(n_5046),
.A2(n_5069),
.B1(n_4883),
.B2(n_4884),
.C1(n_4893),
.C2(n_4888),
.Y(n_6086)
);

AOI22xp5_ASAP7_75t_L g6087 ( 
.A1(n_4567),
.A2(n_4573),
.B1(n_5046),
.B2(n_5360),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5249),
.Y(n_6088)
);

AOI21xp5_ASAP7_75t_L g6089 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5249),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5249),
.Y(n_6091)
);

A2O1A1Ixp33_ASAP7_75t_L g6092 ( 
.A1(n_4966),
.A2(n_4636),
.B(n_5343),
.C(n_5633),
.Y(n_6092)
);

AND2x2_ASAP7_75t_L g6093 ( 
.A(n_5412),
.B(n_5415),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_4887),
.B(n_4889),
.Y(n_6094)
);

BUFx2_ASAP7_75t_L g6095 ( 
.A(n_4502),
.Y(n_6095)
);

AOI221xp5_ASAP7_75t_L g6096 ( 
.A1(n_5370),
.A2(n_5332),
.B1(n_5329),
.B2(n_5260),
.C(n_4980),
.Y(n_6096)
);

CKINVDCx8_ASAP7_75t_R g6097 ( 
.A(n_5666),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5259),
.Y(n_6098)
);

AOI22xp5_ASAP7_75t_L g6099 ( 
.A1(n_4567),
.A2(n_4573),
.B1(n_5360),
.B2(n_5071),
.Y(n_6099)
);

NAND2xp5_ASAP7_75t_SL g6100 ( 
.A(n_5115),
.B(n_5119),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_4887),
.B(n_4889),
.Y(n_6101)
);

AND2x2_ASAP7_75t_L g6102 ( 
.A(n_5412),
.B(n_5415),
.Y(n_6102)
);

O2A1O1Ixp33_ASAP7_75t_L g6103 ( 
.A1(n_5329),
.A2(n_4865),
.B(n_4888),
.C(n_4884),
.Y(n_6103)
);

NAND2xp5_ASAP7_75t_SL g6104 ( 
.A(n_5120),
.B(n_5122),
.Y(n_6104)
);

INVx5_ASAP7_75t_L g6105 ( 
.A(n_4752),
.Y(n_6105)
);

NOR3xp33_ASAP7_75t_L g6106 ( 
.A(n_5084),
.B(n_4908),
.C(n_4980),
.Y(n_6106)
);

AOI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_SL g6108 ( 
.A(n_5120),
.B(n_5122),
.Y(n_6108)
);

BUFx12f_ASAP7_75t_L g6109 ( 
.A(n_4710),
.Y(n_6109)
);

INVx1_ASAP7_75t_SL g6110 ( 
.A(n_4974),
.Y(n_6110)
);

OAI22xp5_ASAP7_75t_L g6111 ( 
.A1(n_4893),
.A2(n_4896),
.B1(n_4895),
.B2(n_5144),
.Y(n_6111)
);

AOI22xp33_ASAP7_75t_L g6112 ( 
.A1(n_5127),
.A2(n_5137),
.B1(n_5071),
.B2(n_4841),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5259),
.Y(n_6113)
);

NAND2xp5_ASAP7_75t_L g6114 ( 
.A(n_4892),
.B(n_4951),
.Y(n_6114)
);

AND2x4_ASAP7_75t_L g6115 ( 
.A(n_5398),
.B(n_5478),
.Y(n_6115)
);

NAND2xp5_ASAP7_75t_SL g6116 ( 
.A(n_5127),
.B(n_5137),
.Y(n_6116)
);

AND2x4_ASAP7_75t_L g6117 ( 
.A(n_5398),
.B(n_5478),
.Y(n_6117)
);

AND2x4_ASAP7_75t_L g6118 ( 
.A(n_5398),
.B(n_5478),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5259),
.Y(n_6119)
);

O2A1O1Ixp33_ASAP7_75t_L g6120 ( 
.A1(n_4895),
.A2(n_4896),
.B(n_4908),
.C(n_5236),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_4892),
.B(n_4951),
.Y(n_6121)
);

NOR2xp33_ASAP7_75t_SL g6122 ( 
.A(n_5397),
.B(n_5474),
.Y(n_6122)
);

HAxp5_ASAP7_75t_L g6123 ( 
.A(n_4721),
.B(n_5189),
.CON(n_6123),
.SN(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5275),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_4953),
.B(n_4979),
.Y(n_6125)
);

NAND2xp5_ASAP7_75t_SL g6126 ( 
.A(n_4547),
.B(n_5061),
.Y(n_6126)
);

NAND3xp33_ASAP7_75t_L g6127 ( 
.A(n_5293),
.B(n_5343),
.C(n_4919),
.Y(n_6127)
);

INVx6_ASAP7_75t_L g6128 ( 
.A(n_4713),
.Y(n_6128)
);

O2A1O1Ixp5_ASAP7_75t_L g6129 ( 
.A1(n_5136),
.A2(n_5236),
.B(n_5250),
.C(n_5166),
.Y(n_6129)
);

INVxp67_ASAP7_75t_L g6130 ( 
.A(n_5238),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5275),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5275),
.Y(n_6132)
);

AOI22xp5_ASAP7_75t_L g6133 ( 
.A1(n_4841),
.A2(n_5170),
.B1(n_4520),
.B2(n_5268),
.Y(n_6133)
);

CKINVDCx11_ASAP7_75t_R g6134 ( 
.A(n_4759),
.Y(n_6134)
);

INVx1_ASAP7_75t_L g6135 ( 
.A(n_5278),
.Y(n_6135)
);

AOI22xp5_ASAP7_75t_L g6136 ( 
.A1(n_5170),
.A2(n_4520),
.B1(n_5268),
.B2(n_5136),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5278),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5278),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_SL g6139 ( 
.A(n_4547),
.B(n_5144),
.Y(n_6139)
);

AND2x2_ASAP7_75t_L g6140 ( 
.A(n_5468),
.B(n_5330),
.Y(n_6140)
);

NOR2xp33_ASAP7_75t_L g6141 ( 
.A(n_5231),
.B(n_5240),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5287),
.Y(n_6142)
);

O2A1O1Ixp33_ASAP7_75t_L g6143 ( 
.A1(n_5098),
.A2(n_5332),
.B(n_5084),
.C(n_5250),
.Y(n_6143)
);

BUFx2_ASAP7_75t_L g6144 ( 
.A(n_4502),
.Y(n_6144)
);

AND2x4_ASAP7_75t_L g6145 ( 
.A(n_5478),
.B(n_5483),
.Y(n_6145)
);

O2A1O1Ixp33_ASAP7_75t_L g6146 ( 
.A1(n_5098),
.A2(n_5582),
.B(n_4919),
.C(n_4920),
.Y(n_6146)
);

INVx4_ASAP7_75t_L g6147 ( 
.A(n_4511),
.Y(n_6147)
);

O2A1O1Ixp33_ASAP7_75t_L g6148 ( 
.A1(n_5582),
.A2(n_4920),
.B(n_4922),
.C(n_4913),
.Y(n_6148)
);

OAI22xp5_ASAP7_75t_L g6149 ( 
.A1(n_5189),
.A2(n_5199),
.B1(n_5210),
.B2(n_4501),
.Y(n_6149)
);

NAND2xp5_ASAP7_75t_SL g6150 ( 
.A(n_4957),
.B(n_4952),
.Y(n_6150)
);

INVx2_ASAP7_75t_SL g6151 ( 
.A(n_5597),
.Y(n_6151)
);

OAI321xp33_ASAP7_75t_L g6152 ( 
.A1(n_5293),
.A2(n_4789),
.A3(n_4717),
.B1(n_4821),
.B2(n_4775),
.C(n_5260),
.Y(n_6152)
);

A2O1A1Ixp33_ASAP7_75t_SL g6153 ( 
.A1(n_5387),
.A2(n_5619),
.B(n_5655),
.C(n_5480),
.Y(n_6153)
);

AOI22xp33_ASAP7_75t_SL g6154 ( 
.A1(n_5301),
.A2(n_5303),
.B1(n_5464),
.B2(n_4803),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_5468),
.B(n_5330),
.Y(n_6155)
);

NAND2xp5_ASAP7_75t_L g6156 ( 
.A(n_4953),
.B(n_4979),
.Y(n_6156)
);

OR2x2_ASAP7_75t_L g6157 ( 
.A(n_4670),
.B(n_4681),
.Y(n_6157)
);

OAI22xp5_ASAP7_75t_L g6158 ( 
.A1(n_5199),
.A2(n_5210),
.B1(n_4501),
.B2(n_4922),
.Y(n_6158)
);

O2A1O1Ixp33_ASAP7_75t_L g6159 ( 
.A1(n_4913),
.A2(n_4928),
.B(n_4944),
.C(n_4926),
.Y(n_6159)
);

NAND2xp5_ASAP7_75t_SL g6160 ( 
.A(n_4957),
.B(n_4952),
.Y(n_6160)
);

O2A1O1Ixp33_ASAP7_75t_L g6161 ( 
.A1(n_4926),
.A2(n_4944),
.B(n_4928),
.C(n_5231),
.Y(n_6161)
);

AOI22xp33_ASAP7_75t_L g6162 ( 
.A1(n_5116),
.A2(n_5132),
.B1(n_5182),
.B2(n_5164),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_SL g6163 ( 
.A(n_5221),
.B(n_4973),
.Y(n_6163)
);

BUFx2_ASAP7_75t_L g6164 ( 
.A(n_4509),
.Y(n_6164)
);

AOI22xp5_ASAP7_75t_L g6165 ( 
.A1(n_5464),
.A2(n_5235),
.B1(n_5184),
.B2(n_5156),
.Y(n_6165)
);

OAI21x1_ASAP7_75t_L g6166 ( 
.A1(n_4862),
.A2(n_5437),
.B(n_5302),
.Y(n_6166)
);

NAND2xp5_ASAP7_75t_L g6167 ( 
.A(n_4991),
.B(n_4996),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5287),
.Y(n_6168)
);

OAI22xp5_ASAP7_75t_L g6169 ( 
.A1(n_4501),
.A2(n_5156),
.B1(n_5336),
.B2(n_5613),
.Y(n_6169)
);

INVx5_ASAP7_75t_L g6170 ( 
.A(n_4752),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_5287),
.Y(n_6171)
);

INVx2_ASAP7_75t_SL g6172 ( 
.A(n_5597),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5288),
.Y(n_6173)
);

AOI21xp5_ASAP7_75t_L g6174 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6174)
);

A2O1A1Ixp33_ASAP7_75t_L g6175 ( 
.A1(n_5633),
.A2(n_5642),
.B(n_5247),
.C(n_5155),
.Y(n_6175)
);

AOI21xp5_ASAP7_75t_L g6176 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5288),
.Y(n_6177)
);

NAND2xp5_ASAP7_75t_SL g6178 ( 
.A(n_5221),
.B(n_4973),
.Y(n_6178)
);

INVx8_ASAP7_75t_L g6179 ( 
.A(n_5207),
.Y(n_6179)
);

NAND2xp5_ASAP7_75t_L g6180 ( 
.A(n_4991),
.B(n_4996),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_SL g6181 ( 
.A(n_4524),
.B(n_5619),
.Y(n_6181)
);

NAND2xp5_ASAP7_75t_L g6182 ( 
.A(n_5012),
.B(n_5027),
.Y(n_6182)
);

AO21x2_ASAP7_75t_L g6183 ( 
.A1(n_4821),
.A2(n_5141),
.B(n_5135),
.Y(n_6183)
);

INVx2_ASAP7_75t_SL g6184 ( 
.A(n_5597),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_5012),
.B(n_5027),
.Y(n_6185)
);

AOI21xp5_ASAP7_75t_L g6186 ( 
.A1(n_4792),
.A2(n_4939),
.B(n_4929),
.Y(n_6186)
);

AOI21xp5_ASAP7_75t_L g6187 ( 
.A1(n_4792),
.A2(n_5009),
.B(n_4939),
.Y(n_6187)
);

INVx2_ASAP7_75t_SL g6188 ( 
.A(n_5597),
.Y(n_6188)
);

AND2x2_ASAP7_75t_L g6189 ( 
.A(n_5468),
.B(n_5330),
.Y(n_6189)
);

AND2x4_ASAP7_75t_L g6190 ( 
.A(n_5478),
.B(n_5483),
.Y(n_6190)
);

INVx5_ASAP7_75t_L g6191 ( 
.A(n_4752),
.Y(n_6191)
);

OAI22xp5_ASAP7_75t_L g6192 ( 
.A1(n_5336),
.A2(n_5613),
.B1(n_5240),
.B2(n_5590),
.Y(n_6192)
);

AND2x4_ASAP7_75t_L g6193 ( 
.A(n_5483),
.B(n_5527),
.Y(n_6193)
);

O2A1O1Ixp5_ASAP7_75t_SL g6194 ( 
.A1(n_5171),
.A2(n_5508),
.B(n_5309),
.C(n_5160),
.Y(n_6194)
);

AND2x4_ASAP7_75t_L g6195 ( 
.A(n_5483),
.B(n_5527),
.Y(n_6195)
);

BUFx2_ASAP7_75t_L g6196 ( 
.A(n_4509),
.Y(n_6196)
);

NOR2xp33_ASAP7_75t_L g6197 ( 
.A(n_5642),
.B(n_5589),
.Y(n_6197)
);

NAND2xp5_ASAP7_75t_L g6198 ( 
.A(n_5030),
.B(n_5041),
.Y(n_6198)
);

NAND2xp5_ASAP7_75t_L g6199 ( 
.A(n_5030),
.B(n_5041),
.Y(n_6199)
);

O2A1O1Ixp33_ASAP7_75t_L g6200 ( 
.A1(n_5497),
.A2(n_4643),
.B(n_5261),
.C(n_5166),
.Y(n_6200)
);

AND2x2_ASAP7_75t_L g6201 ( 
.A(n_5361),
.B(n_4670),
.Y(n_6201)
);

INVxp67_ASAP7_75t_L g6202 ( 
.A(n_5072),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_5361),
.B(n_4681),
.Y(n_6203)
);

AOI222xp33_ASAP7_75t_L g6204 ( 
.A1(n_4812),
.A2(n_4819),
.B1(n_5341),
.B2(n_5351),
.C1(n_5342),
.C2(n_5590),
.Y(n_6204)
);

INVxp67_ASAP7_75t_L g6205 ( 
.A(n_5072),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5288),
.Y(n_6206)
);

OAI22xp5_ASAP7_75t_L g6207 ( 
.A1(n_5301),
.A2(n_5303),
.B1(n_4643),
.B2(n_5477),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_5078),
.B(n_4482),
.Y(n_6208)
);

INVxp67_ASAP7_75t_SL g6209 ( 
.A(n_4949),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5289),
.Y(n_6210)
);

AOI21xp5_ASAP7_75t_L g6211 ( 
.A1(n_5009),
.A2(n_5181),
.B(n_5034),
.Y(n_6211)
);

A2O1A1Ixp33_ASAP7_75t_L g6212 ( 
.A1(n_5247),
.A2(n_5155),
.B(n_5235),
.C(n_5184),
.Y(n_6212)
);

INVx2_ASAP7_75t_SL g6213 ( 
.A(n_5597),
.Y(n_6213)
);

INVx2_ASAP7_75t_SL g6214 ( 
.A(n_5597),
.Y(n_6214)
);

INVx5_ASAP7_75t_SL g6215 ( 
.A(n_5397),
.Y(n_6215)
);

AND2x4_ASAP7_75t_L g6216 ( 
.A(n_5483),
.B(n_5527),
.Y(n_6216)
);

AOI22xp33_ASAP7_75t_L g6217 ( 
.A1(n_5116),
.A2(n_5132),
.B1(n_5182),
.B2(n_5164),
.Y(n_6217)
);

NAND2xp5_ASAP7_75t_L g6218 ( 
.A(n_5078),
.B(n_4482),
.Y(n_6218)
);

INVx3_ASAP7_75t_L g6219 ( 
.A(n_4640),
.Y(n_6219)
);

HB1xp67_ASAP7_75t_L g6220 ( 
.A(n_4509),
.Y(n_6220)
);

OR2x6_ASAP7_75t_L g6221 ( 
.A(n_4515),
.B(n_4698),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_5289),
.Y(n_6222)
);

INVx4_ASAP7_75t_L g6223 ( 
.A(n_4511),
.Y(n_6223)
);

NOR2xp67_ASAP7_75t_SL g6224 ( 
.A(n_5587),
.B(n_5666),
.Y(n_6224)
);

BUFx8_ASAP7_75t_L g6225 ( 
.A(n_4772),
.Y(n_6225)
);

AND2x4_ASAP7_75t_L g6226 ( 
.A(n_5483),
.B(n_5527),
.Y(n_6226)
);

INVx5_ASAP7_75t_L g6227 ( 
.A(n_4752),
.Y(n_6227)
);

CKINVDCx8_ASAP7_75t_R g6228 ( 
.A(n_5666),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_5289),
.Y(n_6229)
);

OR2x6_ASAP7_75t_L g6230 ( 
.A(n_4515),
.B(n_4698),
.Y(n_6230)
);

INVx3_ASAP7_75t_L g6231 ( 
.A(n_4640),
.Y(n_6231)
);

AOI21xp5_ASAP7_75t_L g6232 ( 
.A1(n_5009),
.A2(n_5181),
.B(n_5034),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_5297),
.Y(n_6233)
);

AOI22xp5_ASAP7_75t_L g6234 ( 
.A1(n_4812),
.A2(n_4819),
.B1(n_5083),
.B2(n_5257),
.Y(n_6234)
);

CKINVDCx5p33_ASAP7_75t_R g6235 ( 
.A(n_4906),
.Y(n_6235)
);

NAND2xp5_ASAP7_75t_L g6236 ( 
.A(n_4482),
.B(n_4483),
.Y(n_6236)
);

AOI21xp5_ASAP7_75t_L g6237 ( 
.A1(n_5009),
.A2(n_5181),
.B(n_5034),
.Y(n_6237)
);

INVx3_ASAP7_75t_L g6238 ( 
.A(n_4644),
.Y(n_6238)
);

NAND2xp5_ASAP7_75t_L g6239 ( 
.A(n_4483),
.B(n_4484),
.Y(n_6239)
);

AOI21xp5_ASAP7_75t_L g6240 ( 
.A1(n_5009),
.A2(n_5181),
.B(n_5034),
.Y(n_6240)
);

AOI22xp33_ASAP7_75t_L g6241 ( 
.A1(n_5271),
.A2(n_5295),
.B1(n_5257),
.B2(n_5499),
.Y(n_6241)
);

BUFx2_ASAP7_75t_L g6242 ( 
.A(n_4523),
.Y(n_6242)
);

BUFx3_ASAP7_75t_L g6243 ( 
.A(n_4799),
.Y(n_6243)
);

O2A1O1Ixp33_ASAP7_75t_L g6244 ( 
.A1(n_5497),
.A2(n_5261),
.B(n_5147),
.C(n_5309),
.Y(n_6244)
);

NOR2xp33_ASAP7_75t_L g6245 ( 
.A(n_5589),
.B(n_5438),
.Y(n_6245)
);

NAND2xp5_ASAP7_75t_L g6246 ( 
.A(n_4483),
.B(n_4484),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_L g6247 ( 
.A(n_4484),
.B(n_4487),
.Y(n_6247)
);

NOR2xp33_ASAP7_75t_SL g6248 ( 
.A(n_5474),
.B(n_4526),
.Y(n_6248)
);

AOI21xp5_ASAP7_75t_L g6249 ( 
.A1(n_5009),
.A2(n_5181),
.B(n_5034),
.Y(n_6249)
);

NOR2xp33_ASAP7_75t_L g6250 ( 
.A(n_5438),
.B(n_5447),
.Y(n_6250)
);

BUFx3_ASAP7_75t_L g6251 ( 
.A(n_4799),
.Y(n_6251)
);

NAND2x1_ASAP7_75t_SL g6252 ( 
.A(n_4882),
.B(n_5043),
.Y(n_6252)
);

INVx2_ASAP7_75t_SL g6253 ( 
.A(n_5597),
.Y(n_6253)
);

BUFx2_ASAP7_75t_L g6254 ( 
.A(n_4523),
.Y(n_6254)
);

NOR2xp33_ASAP7_75t_L g6255 ( 
.A(n_5447),
.B(n_5451),
.Y(n_6255)
);

AND2x4_ASAP7_75t_L g6256 ( 
.A(n_5527),
.B(n_4758),
.Y(n_6256)
);

AOI22xp33_ASAP7_75t_SL g6257 ( 
.A1(n_4803),
.A2(n_5609),
.B1(n_4813),
.B2(n_4817),
.Y(n_6257)
);

INVx1_ASAP7_75t_SL g6258 ( 
.A(n_4974),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_4487),
.B(n_4490),
.Y(n_6259)
);

A2O1A1Ixp33_ASAP7_75t_L g6260 ( 
.A1(n_5609),
.A2(n_4803),
.B(n_5480),
.C(n_4813),
.Y(n_6260)
);

INVx1_ASAP7_75t_L g6261 ( 
.A(n_5297),
.Y(n_6261)
);

CKINVDCx6p67_ASAP7_75t_R g6262 ( 
.A(n_4521),
.Y(n_6262)
);

INVx4_ASAP7_75t_L g6263 ( 
.A(n_4526),
.Y(n_6263)
);

INVx3_ASAP7_75t_L g6264 ( 
.A(n_4644),
.Y(n_6264)
);

NOR2xp33_ASAP7_75t_L g6265 ( 
.A(n_5451),
.B(n_5458),
.Y(n_6265)
);

OAI22xp5_ASAP7_75t_L g6266 ( 
.A1(n_5477),
.A2(n_5481),
.B1(n_5149),
.B2(n_5467),
.Y(n_6266)
);

BUFx8_ASAP7_75t_L g6267 ( 
.A(n_4772),
.Y(n_6267)
);

BUFx3_ASAP7_75t_L g6268 ( 
.A(n_4799),
.Y(n_6268)
);

HB1xp67_ASAP7_75t_L g6269 ( 
.A(n_4523),
.Y(n_6269)
);

OR2x6_ASAP7_75t_L g6270 ( 
.A(n_4698),
.B(n_4752),
.Y(n_6270)
);

O2A1O1Ixp33_ASAP7_75t_L g6271 ( 
.A1(n_5147),
.A2(n_5262),
.B(n_4947),
.C(n_5187),
.Y(n_6271)
);

INVx5_ASAP7_75t_L g6272 ( 
.A(n_4752),
.Y(n_6272)
);

AND2x4_ASAP7_75t_L g6273 ( 
.A(n_5527),
.B(n_4758),
.Y(n_6273)
);

A2O1A1Ixp33_ASAP7_75t_L g6274 ( 
.A1(n_4803),
.A2(n_4817),
.B(n_4827),
.C(n_4787),
.Y(n_6274)
);

CKINVDCx5p33_ASAP7_75t_R g6275 ( 
.A(n_4906),
.Y(n_6275)
);

O2A1O1Ixp33_ASAP7_75t_L g6276 ( 
.A1(n_5262),
.A2(n_4947),
.B(n_5187),
.C(n_5186),
.Y(n_6276)
);

AOI22xp33_ASAP7_75t_L g6277 ( 
.A1(n_5271),
.A2(n_5295),
.B1(n_5499),
.B2(n_5312),
.Y(n_6277)
);

O2A1O1Ixp33_ASAP7_75t_L g6278 ( 
.A1(n_5188),
.A2(n_5197),
.B(n_5206),
.C(n_5204),
.Y(n_6278)
);

NOR2xp33_ASAP7_75t_L g6279 ( 
.A(n_5458),
.B(n_4498),
.Y(n_6279)
);

AND2x4_ASAP7_75t_L g6280 ( 
.A(n_4758),
.B(n_4644),
.Y(n_6280)
);

OAI21xp5_ASAP7_75t_L g6281 ( 
.A1(n_4959),
.A2(n_5352),
.B(n_5203),
.Y(n_6281)
);

INVx3_ASAP7_75t_L g6282 ( 
.A(n_4644),
.Y(n_6282)
);

INVx3_ASAP7_75t_SL g6283 ( 
.A(n_5009),
.Y(n_6283)
);

AOI21xp5_ASAP7_75t_L g6284 ( 
.A1(n_5034),
.A2(n_5194),
.B(n_5181),
.Y(n_6284)
);

BUFx3_ASAP7_75t_L g6285 ( 
.A(n_4799),
.Y(n_6285)
);

O2A1O1Ixp33_ASAP7_75t_L g6286 ( 
.A1(n_5188),
.A2(n_5197),
.B(n_5206),
.C(n_5204),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_5361),
.B(n_5507),
.Y(n_6287)
);

NAND2xp5_ASAP7_75t_L g6288 ( 
.A(n_4487),
.B(n_4490),
.Y(n_6288)
);

OR2x6_ASAP7_75t_SL g6289 ( 
.A(n_4981),
.B(n_5310),
.Y(n_6289)
);

HB1xp67_ASAP7_75t_L g6290 ( 
.A(n_4536),
.Y(n_6290)
);

INVx3_ASAP7_75t_L g6291 ( 
.A(n_4644),
.Y(n_6291)
);

NAND2xp5_ASAP7_75t_SL g6292 ( 
.A(n_5721),
.B(n_4513),
.Y(n_6292)
);

NAND2xp5_ASAP7_75t_L g6293 ( 
.A(n_4490),
.B(n_4525),
.Y(n_6293)
);

NOR2xp67_ASAP7_75t_L g6294 ( 
.A(n_4510),
.B(n_4767),
.Y(n_6294)
);

AOI21x1_ASAP7_75t_L g6295 ( 
.A1(n_4862),
.A2(n_5171),
.B(n_4864),
.Y(n_6295)
);

AOI22xp33_ASAP7_75t_L g6296 ( 
.A1(n_5311),
.A2(n_5313),
.B1(n_5321),
.B2(n_5312),
.Y(n_6296)
);

AND2x2_ASAP7_75t_L g6297 ( 
.A(n_5507),
.B(n_5511),
.Y(n_6297)
);

AOI21x1_ASAP7_75t_L g6298 ( 
.A1(n_4852),
.A2(n_4976),
.B(n_4864),
.Y(n_6298)
);

AND2x2_ASAP7_75t_L g6299 ( 
.A(n_5507),
.B(n_5511),
.Y(n_6299)
);

CKINVDCx5p33_ASAP7_75t_R g6300 ( 
.A(n_4978),
.Y(n_6300)
);

AOI221xp5_ASAP7_75t_L g6301 ( 
.A1(n_4812),
.A2(n_4819),
.B1(n_4498),
.B2(n_4499),
.C(n_4981),
.Y(n_6301)
);

AOI22xp33_ASAP7_75t_L g6302 ( 
.A1(n_5311),
.A2(n_5313),
.B1(n_5323),
.B2(n_5321),
.Y(n_6302)
);

AND2x4_ASAP7_75t_L g6303 ( 
.A(n_4758),
.B(n_4644),
.Y(n_6303)
);

AOI21xp5_ASAP7_75t_L g6304 ( 
.A1(n_5034),
.A2(n_5194),
.B(n_5181),
.Y(n_6304)
);

AOI22xp5_ASAP7_75t_L g6305 ( 
.A1(n_5083),
.A2(n_5446),
.B1(n_5467),
.B2(n_5453),
.Y(n_6305)
);

AOI21xp5_ASAP7_75t_L g6306 ( 
.A1(n_5194),
.A2(n_5335),
.B(n_5200),
.Y(n_6306)
);

INVx3_ASAP7_75t_L g6307 ( 
.A(n_4645),
.Y(n_6307)
);

INVx5_ASAP7_75t_L g6308 ( 
.A(n_4698),
.Y(n_6308)
);

NAND2xp5_ASAP7_75t_L g6309 ( 
.A(n_4525),
.B(n_4529),
.Y(n_6309)
);

INVx2_ASAP7_75t_SL g6310 ( 
.A(n_5597),
.Y(n_6310)
);

INVxp67_ASAP7_75t_SL g6311 ( 
.A(n_5146),
.Y(n_6311)
);

OR2x2_ASAP7_75t_L g6312 ( 
.A(n_5201),
.B(n_5239),
.Y(n_6312)
);

AND2x4_ASAP7_75t_L g6313 ( 
.A(n_4758),
.B(n_4645),
.Y(n_6313)
);

BUFx2_ASAP7_75t_L g6314 ( 
.A(n_4536),
.Y(n_6314)
);

NOR2xp33_ASAP7_75t_L g6315 ( 
.A(n_4499),
.B(n_5215),
.Y(n_6315)
);

AOI21xp5_ASAP7_75t_L g6316 ( 
.A1(n_5194),
.A2(n_5335),
.B(n_5200),
.Y(n_6316)
);

NAND2xp5_ASAP7_75t_L g6317 ( 
.A(n_4525),
.B(n_4529),
.Y(n_6317)
);

CKINVDCx11_ASAP7_75t_R g6318 ( 
.A(n_4759),
.Y(n_6318)
);

INVx5_ASAP7_75t_L g6319 ( 
.A(n_4698),
.Y(n_6319)
);

INVxp67_ASAP7_75t_SL g6320 ( 
.A(n_5146),
.Y(n_6320)
);

AND2x2_ASAP7_75t_L g6321 ( 
.A(n_5511),
.B(n_5531),
.Y(n_6321)
);

O2A1O1Ixp33_ASAP7_75t_SL g6322 ( 
.A1(n_5000),
.A2(n_4891),
.B(n_4916),
.C(n_4859),
.Y(n_6322)
);

INVx4_ASAP7_75t_L g6323 ( 
.A(n_4526),
.Y(n_6323)
);

BUFx2_ASAP7_75t_L g6324 ( 
.A(n_4536),
.Y(n_6324)
);

INVx1_ASAP7_75t_SL g6325 ( 
.A(n_4983),
.Y(n_6325)
);

INVx3_ASAP7_75t_L g6326 ( 
.A(n_4645),
.Y(n_6326)
);

OR2x6_ASAP7_75t_SL g6327 ( 
.A(n_5310),
.B(n_4787),
.Y(n_6327)
);

INVx3_ASAP7_75t_L g6328 ( 
.A(n_4645),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_L g6329 ( 
.A(n_4529),
.B(n_4530),
.Y(n_6329)
);

NOR2xp33_ASAP7_75t_L g6330 ( 
.A(n_5215),
.B(n_5455),
.Y(n_6330)
);

O2A1O1Ixp33_ASAP7_75t_L g6331 ( 
.A1(n_5352),
.A2(n_5000),
.B(n_4767),
.C(n_4768),
.Y(n_6331)
);

OR2x6_ASAP7_75t_L g6332 ( 
.A(n_4698),
.B(n_4760),
.Y(n_6332)
);

BUFx2_ASAP7_75t_L g6333 ( 
.A(n_4543),
.Y(n_6333)
);

AOI21xp5_ASAP7_75t_L g6334 ( 
.A1(n_5194),
.A2(n_5335),
.B(n_5200),
.Y(n_6334)
);

OR2x6_ASAP7_75t_L g6335 ( 
.A(n_4760),
.B(n_4605),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_4530),
.B(n_4535),
.Y(n_6336)
);

INVx4_ASAP7_75t_L g6337 ( 
.A(n_4526),
.Y(n_6337)
);

INVx2_ASAP7_75t_SL g6338 ( 
.A(n_4875),
.Y(n_6338)
);

BUFx2_ASAP7_75t_L g6339 ( 
.A(n_4543),
.Y(n_6339)
);

INVx4_ASAP7_75t_L g6340 ( 
.A(n_4526),
.Y(n_6340)
);

AOI21xp5_ASAP7_75t_L g6341 ( 
.A1(n_5194),
.A2(n_5335),
.B(n_5200),
.Y(n_6341)
);

OAI22xp5_ASAP7_75t_L g6342 ( 
.A1(n_5481),
.A2(n_5149),
.B1(n_5446),
.B2(n_5489),
.Y(n_6342)
);

OAI22xp5_ASAP7_75t_L g6343 ( 
.A1(n_5489),
.A2(n_5296),
.B1(n_5392),
.B2(n_5524),
.Y(n_6343)
);

INVx2_ASAP7_75t_L g6344 ( 
.A(n_5212),
.Y(n_6344)
);

BUFx2_ASAP7_75t_L g6345 ( 
.A(n_4543),
.Y(n_6345)
);

BUFx4f_ASAP7_75t_SL g6346 ( 
.A(n_4780),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_5212),
.Y(n_6347)
);

AOI22xp5_ASAP7_75t_L g6348 ( 
.A1(n_5443),
.A2(n_5453),
.B1(n_5500),
.B2(n_5473),
.Y(n_6348)
);

BUFx12f_ASAP7_75t_L g6349 ( 
.A(n_4710),
.Y(n_6349)
);

AOI22xp33_ASAP7_75t_SL g6350 ( 
.A1(n_4803),
.A2(n_4830),
.B1(n_4832),
.B2(n_4827),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_5531),
.B(n_5556),
.Y(n_6351)
);

AND2x4_ASAP7_75t_L g6352 ( 
.A(n_4663),
.B(n_4671),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_5212),
.Y(n_6353)
);

O2A1O1Ixp33_ASAP7_75t_L g6354 ( 
.A1(n_4510),
.A2(n_4768),
.B(n_4771),
.C(n_4650),
.Y(n_6354)
);

NOR2xp33_ASAP7_75t_L g6355 ( 
.A(n_5455),
.B(n_5602),
.Y(n_6355)
);

HB1xp67_ASAP7_75t_L g6356 ( 
.A(n_4546),
.Y(n_6356)
);

OAI22xp5_ASAP7_75t_L g6357 ( 
.A1(n_5296),
.A2(n_5392),
.B1(n_5524),
.B2(n_5341),
.Y(n_6357)
);

AND2x4_ASAP7_75t_L g6358 ( 
.A(n_4663),
.B(n_4671),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_4530),
.B(n_4535),
.Y(n_6359)
);

OAI22xp5_ASAP7_75t_L g6360 ( 
.A1(n_5342),
.A2(n_5351),
.B1(n_5348),
.B2(n_4959),
.Y(n_6360)
);

OR2x6_ASAP7_75t_L g6361 ( 
.A(n_4760),
.B(n_4605),
.Y(n_6361)
);

NAND2xp5_ASAP7_75t_L g6362 ( 
.A(n_4535),
.B(n_4553),
.Y(n_6362)
);

AOI21xp5_ASAP7_75t_L g6363 ( 
.A1(n_5194),
.A2(n_5335),
.B(n_5200),
.Y(n_6363)
);

BUFx12f_ASAP7_75t_L g6364 ( 
.A(n_4731),
.Y(n_6364)
);

AOI21x1_ASAP7_75t_L g6365 ( 
.A1(n_4852),
.A2(n_5040),
.B(n_4976),
.Y(n_6365)
);

A2O1A1Ixp33_ASAP7_75t_L g6366 ( 
.A1(n_4830),
.A2(n_4833),
.B(n_4837),
.C(n_4832),
.Y(n_6366)
);

BUFx2_ASAP7_75t_L g6367 ( 
.A(n_4546),
.Y(n_6367)
);

AO22x1_ASAP7_75t_L g6368 ( 
.A1(n_5697),
.A2(n_5279),
.B1(n_5366),
.B2(n_5207),
.Y(n_6368)
);

AND2x2_ASAP7_75t_L g6369 ( 
.A(n_5531),
.B(n_5556),
.Y(n_6369)
);

NOR2xp33_ASAP7_75t_L g6370 ( 
.A(n_5602),
.B(n_5348),
.Y(n_6370)
);

INVx4_ASAP7_75t_L g6371 ( 
.A(n_4570),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_4553),
.B(n_4572),
.Y(n_6372)
);

CKINVDCx5p33_ASAP7_75t_R g6373 ( 
.A(n_4978),
.Y(n_6373)
);

AOI22xp33_ASAP7_75t_L g6374 ( 
.A1(n_5323),
.A2(n_5325),
.B1(n_5324),
.B2(n_5310),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_5212),
.Y(n_6375)
);

INVx2_ASAP7_75t_L g6376 ( 
.A(n_5216),
.Y(n_6376)
);

NAND2xp5_ASAP7_75t_L g6377 ( 
.A(n_4553),
.B(n_4572),
.Y(n_6377)
);

OAI22xp5_ASAP7_75t_L g6378 ( 
.A1(n_4959),
.A2(n_5599),
.B1(n_4778),
.B2(n_4784),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_4546),
.Y(n_6379)
);

O2A1O1Ixp33_ASAP7_75t_L g6380 ( 
.A1(n_4771),
.A2(n_4650),
.B(n_5573),
.C(n_5618),
.Y(n_6380)
);

INVx2_ASAP7_75t_L g6381 ( 
.A(n_5216),
.Y(n_6381)
);

OR2x2_ASAP7_75t_L g6382 ( 
.A(n_5201),
.B(n_5239),
.Y(n_6382)
);

A2O1A1Ixp33_ASAP7_75t_L g6383 ( 
.A1(n_4833),
.A2(n_4837),
.B(n_5599),
.C(n_5618),
.Y(n_6383)
);

CKINVDCx16_ASAP7_75t_R g6384 ( 
.A(n_4521),
.Y(n_6384)
);

NAND2x1p5_ASAP7_75t_L g6385 ( 
.A(n_4570),
.B(n_4628),
.Y(n_6385)
);

OAI22xp5_ASAP7_75t_L g6386 ( 
.A1(n_4778),
.A2(n_4784),
.B1(n_4669),
.B2(n_5559),
.Y(n_6386)
);

A2O1A1Ixp33_ASAP7_75t_L g6387 ( 
.A1(n_5017),
.A2(n_5066),
.B(n_4570),
.C(n_4656),
.Y(n_6387)
);

AO22x1_ASAP7_75t_L g6388 ( 
.A1(n_5697),
.A2(n_5279),
.B1(n_5366),
.B2(n_5207),
.Y(n_6388)
);

INVx5_ASAP7_75t_L g6389 ( 
.A(n_4605),
.Y(n_6389)
);

AOI22xp33_ASAP7_75t_L g6390 ( 
.A1(n_5324),
.A2(n_5325),
.B1(n_4809),
.B2(n_5646),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_4572),
.B(n_4576),
.Y(n_6391)
);

O2A1O1Ixp33_ASAP7_75t_L g6392 ( 
.A1(n_5573),
.A2(n_5501),
.B(n_5504),
.C(n_5498),
.Y(n_6392)
);

OR2x6_ASAP7_75t_L g6393 ( 
.A(n_4760),
.B(n_4605),
.Y(n_6393)
);

AOI21xp5_ASAP7_75t_L g6394 ( 
.A1(n_5200),
.A2(n_5475),
.B(n_5335),
.Y(n_6394)
);

NOR2xp33_ASAP7_75t_L g6395 ( 
.A(n_5459),
.B(n_5485),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_5216),
.Y(n_6396)
);

BUFx2_ASAP7_75t_L g6397 ( 
.A(n_4586),
.Y(n_6397)
);

CKINVDCx5p33_ASAP7_75t_R g6398 ( 
.A(n_5032),
.Y(n_6398)
);

NAND2xp5_ASAP7_75t_L g6399 ( 
.A(n_4576),
.B(n_4578),
.Y(n_6399)
);

AOI21xp5_ASAP7_75t_L g6400 ( 
.A1(n_5200),
.A2(n_5475),
.B(n_5335),
.Y(n_6400)
);

O2A1O1Ixp33_ASAP7_75t_L g6401 ( 
.A1(n_5498),
.A2(n_5504),
.B(n_5515),
.C(n_5501),
.Y(n_6401)
);

BUFx8_ASAP7_75t_SL g6402 ( 
.A(n_4731),
.Y(n_6402)
);

AOI21xp5_ASAP7_75t_L g6403 ( 
.A1(n_5475),
.A2(n_5509),
.B(n_5515),
.Y(n_6403)
);

A2O1A1Ixp33_ASAP7_75t_SL g6404 ( 
.A1(n_5655),
.A2(n_5637),
.B(n_5663),
.C(n_5658),
.Y(n_6404)
);

INVx4_ASAP7_75t_L g6405 ( 
.A(n_4570),
.Y(n_6405)
);

OAI22xp5_ASAP7_75t_L g6406 ( 
.A1(n_4669),
.A2(n_5559),
.B1(n_5043),
.B2(n_4882),
.Y(n_6406)
);

OR2x2_ASAP7_75t_L g6407 ( 
.A(n_4766),
.B(n_4897),
.Y(n_6407)
);

AOI222xp33_ASAP7_75t_L g6408 ( 
.A1(n_5157),
.A2(n_5522),
.B1(n_5443),
.B2(n_5500),
.C1(n_5473),
.C2(n_5577),
.Y(n_6408)
);

OAI21xp33_ASAP7_75t_L g6409 ( 
.A1(n_5516),
.A2(n_5546),
.B(n_5530),
.Y(n_6409)
);

NOR2xp33_ASAP7_75t_L g6410 ( 
.A(n_5459),
.B(n_5485),
.Y(n_6410)
);

INVx4_ASAP7_75t_L g6411 ( 
.A(n_4570),
.Y(n_6411)
);

OAI22xp5_ASAP7_75t_L g6412 ( 
.A1(n_4669),
.A2(n_5043),
.B1(n_4882),
.B2(n_5017),
.Y(n_6412)
);

OR2x2_ASAP7_75t_L g6413 ( 
.A(n_4766),
.B(n_4897),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_L g6414 ( 
.A(n_4576),
.B(n_4578),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_4578),
.B(n_4588),
.Y(n_6415)
);

INVx5_ASAP7_75t_L g6416 ( 
.A(n_4605),
.Y(n_6416)
);

HB1xp67_ASAP7_75t_L g6417 ( 
.A(n_4586),
.Y(n_6417)
);

NAND2xp5_ASAP7_75t_L g6418 ( 
.A(n_4588),
.B(n_4595),
.Y(n_6418)
);

NOR2xp67_ASAP7_75t_L g6419 ( 
.A(n_5508),
.B(n_5726),
.Y(n_6419)
);

BUFx2_ASAP7_75t_L g6420 ( 
.A(n_4586),
.Y(n_6420)
);

BUFx2_ASAP7_75t_L g6421 ( 
.A(n_4601),
.Y(n_6421)
);

AOI22xp5_ASAP7_75t_L g6422 ( 
.A1(n_5522),
.A2(n_5157),
.B1(n_4809),
.B2(n_5626),
.Y(n_6422)
);

OAI22xp5_ASAP7_75t_L g6423 ( 
.A1(n_4669),
.A2(n_5043),
.B1(n_4882),
.B2(n_5066),
.Y(n_6423)
);

HB1xp67_ASAP7_75t_L g6424 ( 
.A(n_4601),
.Y(n_6424)
);

BUFx2_ASAP7_75t_L g6425 ( 
.A(n_4601),
.Y(n_6425)
);

AOI22xp5_ASAP7_75t_L g6426 ( 
.A1(n_5157),
.A2(n_4809),
.B1(n_5626),
.B2(n_5474),
.Y(n_6426)
);

NOR2xp33_ASAP7_75t_L g6427 ( 
.A(n_5631),
.B(n_5304),
.Y(n_6427)
);

AOI21xp5_ASAP7_75t_L g6428 ( 
.A1(n_5475),
.A2(n_5509),
.B(n_5516),
.Y(n_6428)
);

BUFx2_ASAP7_75t_L g6429 ( 
.A(n_4607),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_5556),
.B(n_4552),
.Y(n_6430)
);

BUFx4f_ASAP7_75t_L g6431 ( 
.A(n_5207),
.Y(n_6431)
);

HB1xp67_ASAP7_75t_L g6432 ( 
.A(n_4607),
.Y(n_6432)
);

NOR2xp67_ASAP7_75t_L g6433 ( 
.A(n_5726),
.B(n_5666),
.Y(n_6433)
);

NOR2xp33_ASAP7_75t_SL g6434 ( 
.A(n_4628),
.B(n_4656),
.Y(n_6434)
);

INVx5_ASAP7_75t_L g6435 ( 
.A(n_4605),
.Y(n_6435)
);

INVx5_ASAP7_75t_L g6436 ( 
.A(n_4605),
.Y(n_6436)
);

AOI21xp33_ASAP7_75t_L g6437 ( 
.A1(n_4809),
.A2(n_5141),
.B(n_5135),
.Y(n_6437)
);

NAND2xp5_ASAP7_75t_SL g6438 ( 
.A(n_5721),
.B(n_4513),
.Y(n_6438)
);

O2A1O1Ixp33_ASAP7_75t_L g6439 ( 
.A1(n_5530),
.A2(n_5549),
.B(n_5565),
.C(n_5546),
.Y(n_6439)
);

BUFx2_ASAP7_75t_L g6440 ( 
.A(n_4607),
.Y(n_6440)
);

NAND2xp5_ASAP7_75t_L g6441 ( 
.A(n_4588),
.B(n_4595),
.Y(n_6441)
);

O2A1O1Ixp5_ASAP7_75t_L g6442 ( 
.A1(n_5620),
.A2(n_5565),
.B(n_5569),
.C(n_5549),
.Y(n_6442)
);

AOI221xp5_ASAP7_75t_L g6443 ( 
.A1(n_5246),
.A2(n_5254),
.B1(n_5484),
.B2(n_5423),
.C(n_5135),
.Y(n_6443)
);

AND2x2_ASAP7_75t_SL g6444 ( 
.A(n_4628),
.B(n_4656),
.Y(n_6444)
);

AND2x2_ASAP7_75t_L g6445 ( 
.A(n_4552),
.B(n_4652),
.Y(n_6445)
);

CKINVDCx14_ASAP7_75t_R g6446 ( 
.A(n_4751),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_4595),
.B(n_4615),
.Y(n_6447)
);

NAND2xp5_ASAP7_75t_L g6448 ( 
.A(n_4615),
.B(n_4631),
.Y(n_6448)
);

AOI22xp5_ASAP7_75t_L g6449 ( 
.A1(n_4809),
.A2(n_5577),
.B1(n_5537),
.B2(n_5535),
.Y(n_6449)
);

OAI22xp5_ASAP7_75t_L g6450 ( 
.A1(n_5475),
.A2(n_5423),
.B1(n_5484),
.B2(n_5494),
.Y(n_6450)
);

NAND2xp5_ASAP7_75t_L g6451 ( 
.A(n_4615),
.B(n_4631),
.Y(n_6451)
);

NOR2xp33_ASAP7_75t_L g6452 ( 
.A(n_5631),
.B(n_5304),
.Y(n_6452)
);

CKINVDCx5p33_ASAP7_75t_R g6453 ( 
.A(n_5032),
.Y(n_6453)
);

AOI21xp5_ASAP7_75t_L g6454 ( 
.A1(n_5475),
.A2(n_5569),
.B(n_5203),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_4552),
.B(n_4652),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_SL g6456 ( 
.A(n_4649),
.B(n_4692),
.Y(n_6456)
);

NAND2xp5_ASAP7_75t_SL g6457 ( 
.A(n_4649),
.B(n_4692),
.Y(n_6457)
);

A2O1A1Ixp33_ASAP7_75t_L g6458 ( 
.A1(n_4628),
.A2(n_4656),
.B(n_4938),
.C(n_4915),
.Y(n_6458)
);

NOR2xp67_ASAP7_75t_SL g6459 ( 
.A(n_5587),
.B(n_5666),
.Y(n_6459)
);

NAND2xp5_ASAP7_75t_L g6460 ( 
.A(n_4631),
.B(n_4638),
.Y(n_6460)
);

NAND2xp5_ASAP7_75t_L g6461 ( 
.A(n_4638),
.B(n_4654),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_L g6462 ( 
.A(n_4638),
.B(n_4654),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_4654),
.B(n_4662),
.Y(n_6463)
);

OAI22xp5_ASAP7_75t_L g6464 ( 
.A1(n_5475),
.A2(n_5423),
.B1(n_5484),
.B2(n_5494),
.Y(n_6464)
);

AOI21xp5_ASAP7_75t_L g6465 ( 
.A1(n_5203),
.A2(n_5437),
.B(n_5302),
.Y(n_6465)
);

AOI222xp33_ASAP7_75t_L g6466 ( 
.A1(n_5668),
.A2(n_5506),
.B1(n_5646),
.B2(n_5628),
.C1(n_5624),
.C2(n_5254),
.Y(n_6466)
);

OAI21x1_ASAP7_75t_L g6467 ( 
.A1(n_5302),
.A2(n_5465),
.B(n_5437),
.Y(n_6467)
);

OR2x6_ASAP7_75t_L g6468 ( 
.A(n_4760),
.B(n_5677),
.Y(n_6468)
);

AOI22xp5_ASAP7_75t_L g6469 ( 
.A1(n_5535),
.A2(n_5610),
.B1(n_5537),
.B2(n_5670),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_4662),
.B(n_4673),
.Y(n_6470)
);

AOI22xp33_ASAP7_75t_SL g6471 ( 
.A1(n_4756),
.A2(n_5246),
.B1(n_5141),
.B2(n_5153),
.Y(n_6471)
);

A2O1A1Ixp33_ASAP7_75t_L g6472 ( 
.A1(n_4628),
.A2(n_4656),
.B(n_4938),
.C(n_4915),
.Y(n_6472)
);

INVx1_ASAP7_75t_SL g6473 ( 
.A(n_4983),
.Y(n_6473)
);

OR2x2_ASAP7_75t_L g6474 ( 
.A(n_4897),
.B(n_4909),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_SL g6475 ( 
.A(n_4756),
.B(n_4915),
.Y(n_6475)
);

CKINVDCx5p33_ASAP7_75t_R g6476 ( 
.A(n_5284),
.Y(n_6476)
);

INVx2_ASAP7_75t_SL g6477 ( 
.A(n_4875),
.Y(n_6477)
);

OAI22xp5_ASAP7_75t_L g6478 ( 
.A1(n_5494),
.A2(n_5547),
.B1(n_5523),
.B2(n_5465),
.Y(n_6478)
);

AND2x4_ASAP7_75t_L g6479 ( 
.A(n_4674),
.B(n_5317),
.Y(n_6479)
);

OAI21xp5_ASAP7_75t_L g6480 ( 
.A1(n_4825),
.A2(n_4701),
.B(n_5040),
.Y(n_6480)
);

INVx5_ASAP7_75t_L g6481 ( 
.A(n_4760),
.Y(n_6481)
);

AOI22xp33_ASAP7_75t_L g6482 ( 
.A1(n_5697),
.A2(n_5153),
.B1(n_5150),
.B2(n_5669),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_SL g6483 ( 
.A(n_4915),
.B(n_4938),
.Y(n_6483)
);

A2O1A1Ixp33_ASAP7_75t_L g6484 ( 
.A1(n_4915),
.A2(n_4938),
.B(n_5214),
.C(n_5198),
.Y(n_6484)
);

INVx8_ASAP7_75t_L g6485 ( 
.A(n_5207),
.Y(n_6485)
);

A2O1A1Ixp33_ASAP7_75t_L g6486 ( 
.A1(n_4938),
.A2(n_5198),
.B(n_5253),
.C(n_5214),
.Y(n_6486)
);

O2A1O1Ixp33_ASAP7_75t_L g6487 ( 
.A1(n_5620),
.A2(n_4701),
.B(n_5263),
.C(n_5563),
.Y(n_6487)
);

AOI21xp5_ASAP7_75t_L g6488 ( 
.A1(n_5465),
.A2(n_5523),
.B(n_4760),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_4652),
.B(n_4870),
.Y(n_6489)
);

A2O1A1Ixp33_ASAP7_75t_L g6490 ( 
.A1(n_5198),
.A2(n_5253),
.B(n_5282),
.C(n_5214),
.Y(n_6490)
);

NOR2xp33_ASAP7_75t_L g6491 ( 
.A(n_5305),
.B(n_5637),
.Y(n_6491)
);

INVx2_ASAP7_75t_SL g6492 ( 
.A(n_4875),
.Y(n_6492)
);

CKINVDCx11_ASAP7_75t_R g6493 ( 
.A(n_4780),
.Y(n_6493)
);

AOI22xp5_ASAP7_75t_L g6494 ( 
.A1(n_5610),
.A2(n_5670),
.B1(n_4606),
.B2(n_4590),
.Y(n_6494)
);

NAND2xp5_ASAP7_75t_L g6495 ( 
.A(n_4662),
.B(n_4673),
.Y(n_6495)
);

NAND2xp5_ASAP7_75t_L g6496 ( 
.A(n_4673),
.B(n_4675),
.Y(n_6496)
);

O2A1O1Ixp33_ASAP7_75t_L g6497 ( 
.A1(n_5263),
.A2(n_5564),
.B(n_5567),
.C(n_5563),
.Y(n_6497)
);

AOI21xp5_ASAP7_75t_L g6498 ( 
.A1(n_5523),
.A2(n_5564),
.B(n_5563),
.Y(n_6498)
);

NAND2xp5_ASAP7_75t_L g6499 ( 
.A(n_4675),
.B(n_4679),
.Y(n_6499)
);

OR2x2_ASAP7_75t_L g6500 ( 
.A(n_4909),
.B(n_5004),
.Y(n_6500)
);

AOI21xp5_ASAP7_75t_L g6501 ( 
.A1(n_5564),
.A2(n_5568),
.B(n_5567),
.Y(n_6501)
);

AOI21xp5_ASAP7_75t_L g6502 ( 
.A1(n_5567),
.A2(n_5570),
.B(n_5568),
.Y(n_6502)
);

O2A1O1Ixp33_ASAP7_75t_L g6503 ( 
.A1(n_5568),
.A2(n_5572),
.B(n_5570),
.C(n_5153),
.Y(n_6503)
);

INVxp67_ASAP7_75t_L g6504 ( 
.A(n_4872),
.Y(n_6504)
);

AOI22xp33_ASAP7_75t_L g6505 ( 
.A1(n_5697),
.A2(n_5150),
.B1(n_5669),
.B2(n_5668),
.Y(n_6505)
);

AOI21xp5_ASAP7_75t_L g6506 ( 
.A1(n_5570),
.A2(n_5572),
.B(n_5644),
.Y(n_6506)
);

NAND2x1p5_ASAP7_75t_L g6507 ( 
.A(n_5198),
.B(n_5214),
.Y(n_6507)
);

O2A1O1Ixp33_ASAP7_75t_L g6508 ( 
.A1(n_5572),
.A2(n_5150),
.B(n_5698),
.C(n_4825),
.Y(n_6508)
);

AOI22xp5_ASAP7_75t_L g6509 ( 
.A1(n_4590),
.A2(n_4606),
.B1(n_5506),
.B2(n_5640),
.Y(n_6509)
);

NOR2xp33_ASAP7_75t_L g6510 ( 
.A(n_5305),
.B(n_5466),
.Y(n_6510)
);

AOI21xp5_ASAP7_75t_L g6511 ( 
.A1(n_5644),
.A2(n_4661),
.B(n_5580),
.Y(n_6511)
);

AOI21xp5_ASAP7_75t_L g6512 ( 
.A1(n_4661),
.A2(n_5584),
.B(n_5580),
.Y(n_6512)
);

NOR2xp33_ASAP7_75t_L g6513 ( 
.A(n_5466),
.B(n_5690),
.Y(n_6513)
);

NAND2xp5_ASAP7_75t_SL g6514 ( 
.A(n_5198),
.B(n_5214),
.Y(n_6514)
);

NOR2xp33_ASAP7_75t_L g6515 ( 
.A(n_5690),
.B(n_5696),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_L g6516 ( 
.A(n_4675),
.B(n_4679),
.Y(n_6516)
);

AOI21xp5_ASAP7_75t_L g6517 ( 
.A1(n_4661),
.A2(n_5591),
.B(n_5584),
.Y(n_6517)
);

AND2x4_ASAP7_75t_L g6518 ( 
.A(n_5317),
.B(n_5554),
.Y(n_6518)
);

NAND2xp5_ASAP7_75t_L g6519 ( 
.A(n_4679),
.B(n_4683),
.Y(n_6519)
);

O2A1O1Ixp33_ASAP7_75t_L g6520 ( 
.A1(n_5698),
.A2(n_4646),
.B(n_5493),
.C(n_5591),
.Y(n_6520)
);

NAND2xp5_ASAP7_75t_L g6521 ( 
.A(n_4683),
.B(n_4697),
.Y(n_6521)
);

OAI22xp5_ASAP7_75t_L g6522 ( 
.A1(n_5547),
.A2(n_5434),
.B1(n_5538),
.B2(n_4891),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_SL g6523 ( 
.A(n_5253),
.B(n_5282),
.Y(n_6523)
);

INVxp67_ASAP7_75t_SL g6524 ( 
.A(n_5160),
.Y(n_6524)
);

OR2x2_ASAP7_75t_L g6525 ( 
.A(n_4909),
.B(n_5004),
.Y(n_6525)
);

NOR2xp33_ASAP7_75t_L g6526 ( 
.A(n_5690),
.B(n_5696),
.Y(n_6526)
);

AOI21xp5_ASAP7_75t_L g6527 ( 
.A1(n_5592),
.A2(n_5654),
.B(n_5648),
.Y(n_6527)
);

NOR2xp33_ASAP7_75t_L g6528 ( 
.A(n_5696),
.B(n_5701),
.Y(n_6528)
);

INVx1_ASAP7_75t_SL g6529 ( 
.A(n_5125),
.Y(n_6529)
);

INVx3_ASAP7_75t_L g6530 ( 
.A(n_4491),
.Y(n_6530)
);

HB1xp67_ASAP7_75t_L g6531 ( 
.A(n_5306),
.Y(n_6531)
);

AOI22xp5_ASAP7_75t_L g6532 ( 
.A1(n_5640),
.A2(n_5635),
.B1(n_5678),
.B2(n_5681),
.Y(n_6532)
);

INVx5_ASAP7_75t_L g6533 ( 
.A(n_4664),
.Y(n_6533)
);

NOR2xp33_ASAP7_75t_L g6534 ( 
.A(n_5701),
.B(n_5561),
.Y(n_6534)
);

HB1xp67_ASAP7_75t_L g6535 ( 
.A(n_5306),
.Y(n_6535)
);

AOI21xp5_ASAP7_75t_L g6536 ( 
.A1(n_5592),
.A2(n_5654),
.B(n_5648),
.Y(n_6536)
);

NAND2xp5_ASAP7_75t_L g6537 ( 
.A(n_4683),
.B(n_4697),
.Y(n_6537)
);

NAND2xp5_ASAP7_75t_L g6538 ( 
.A(n_4697),
.B(n_4699),
.Y(n_6538)
);

BUFx2_ASAP7_75t_L g6539 ( 
.A(n_4686),
.Y(n_6539)
);

INVx1_ASAP7_75t_SL g6540 ( 
.A(n_5125),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_L g6541 ( 
.A(n_4699),
.B(n_4706),
.Y(n_6541)
);

O2A1O1Ixp5_ASAP7_75t_L g6542 ( 
.A1(n_5677),
.A2(n_5625),
.B(n_5650),
.C(n_5657),
.Y(n_6542)
);

OR2x6_ASAP7_75t_L g6543 ( 
.A(n_5677),
.B(n_4734),
.Y(n_6543)
);

AOI21xp5_ASAP7_75t_L g6544 ( 
.A1(n_5636),
.A2(n_5638),
.B(n_4916),
.Y(n_6544)
);

AND2x2_ASAP7_75t_SL g6545 ( 
.A(n_5253),
.B(n_5282),
.Y(n_6545)
);

BUFx2_ASAP7_75t_L g6546 ( 
.A(n_4686),
.Y(n_6546)
);

AND2x2_ASAP7_75t_L g6547 ( 
.A(n_4870),
.B(n_4936),
.Y(n_6547)
);

OAI22xp5_ASAP7_75t_L g6548 ( 
.A1(n_5547),
.A2(n_5434),
.B1(n_5538),
.B2(n_4930),
.Y(n_6548)
);

INVx3_ASAP7_75t_L g6549 ( 
.A(n_4491),
.Y(n_6549)
);

NOR3xp33_ASAP7_75t_L g6550 ( 
.A(n_5345),
.B(n_5353),
.C(n_5493),
.Y(n_6550)
);

HB1xp67_ASAP7_75t_L g6551 ( 
.A(n_5314),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_4699),
.B(n_4706),
.Y(n_6552)
);

A2O1A1Ixp33_ASAP7_75t_SL g6553 ( 
.A1(n_5658),
.A2(n_5664),
.B(n_5663),
.C(n_5722),
.Y(n_6553)
);

BUFx2_ASAP7_75t_L g6554 ( 
.A(n_4836),
.Y(n_6554)
);

AO32x1_ASAP7_75t_L g6555 ( 
.A1(n_4850),
.A2(n_5013),
.A3(n_5023),
.B1(n_4955),
.B2(n_4912),
.Y(n_6555)
);

HB1xp67_ASAP7_75t_L g6556 ( 
.A(n_5314),
.Y(n_6556)
);

A2O1A1Ixp33_ASAP7_75t_SL g6557 ( 
.A1(n_5664),
.A2(n_5722),
.B(n_5576),
.C(n_5611),
.Y(n_6557)
);

BUFx2_ASAP7_75t_L g6558 ( 
.A(n_4836),
.Y(n_6558)
);

INVx1_ASAP7_75t_SL g6559 ( 
.A(n_5434),
.Y(n_6559)
);

O2A1O1Ixp33_ASAP7_75t_L g6560 ( 
.A1(n_4646),
.A2(n_5371),
.B(n_5383),
.C(n_5331),
.Y(n_6560)
);

NOR2xp33_ASAP7_75t_L g6561 ( 
.A(n_5701),
.B(n_5561),
.Y(n_6561)
);

INVx2_ASAP7_75t_SL g6562 ( 
.A(n_4875),
.Y(n_6562)
);

NOR2x1_ASAP7_75t_L g6563 ( 
.A(n_4706),
.B(n_4707),
.Y(n_6563)
);

INVxp67_ASAP7_75t_L g6564 ( 
.A(n_4872),
.Y(n_6564)
);

OAI22xp5_ASAP7_75t_L g6565 ( 
.A1(n_5538),
.A2(n_4930),
.B1(n_4859),
.B2(n_5253),
.Y(n_6565)
);

OAI21x1_ASAP7_75t_L g6566 ( 
.A1(n_5290),
.A2(n_5298),
.B(n_5294),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_4707),
.B(n_4712),
.Y(n_6567)
);

BUFx12f_ASAP7_75t_L g6568 ( 
.A(n_4736),
.Y(n_6568)
);

AOI21xp5_ASAP7_75t_L g6569 ( 
.A1(n_5636),
.A2(n_5638),
.B(n_5226),
.Y(n_6569)
);

AOI22xp33_ASAP7_75t_L g6570 ( 
.A1(n_5647),
.A2(n_5628),
.B1(n_5624),
.B2(n_5688),
.Y(n_6570)
);

INVx3_ASAP7_75t_SL g6571 ( 
.A(n_5666),
.Y(n_6571)
);

CKINVDCx5p33_ASAP7_75t_R g6572 ( 
.A(n_5284),
.Y(n_6572)
);

BUFx2_ASAP7_75t_L g6573 ( 
.A(n_5502),
.Y(n_6573)
);

CKINVDCx5p33_ASAP7_75t_R g6574 ( 
.A(n_5319),
.Y(n_6574)
);

INVx3_ASAP7_75t_L g6575 ( 
.A(n_4491),
.Y(n_6575)
);

OAI22xp5_ASAP7_75t_L g6576 ( 
.A1(n_5538),
.A2(n_5394),
.B1(n_5282),
.B2(n_4750),
.Y(n_6576)
);

INVx3_ASAP7_75t_L g6577 ( 
.A(n_4491),
.Y(n_6577)
);

INVx3_ASAP7_75t_L g6578 ( 
.A(n_4491),
.Y(n_6578)
);

BUFx4f_ASAP7_75t_L g6579 ( 
.A(n_5207),
.Y(n_6579)
);

AOI22xp5_ASAP7_75t_L g6580 ( 
.A1(n_5635),
.A2(n_5678),
.B1(n_5681),
.B2(n_5683),
.Y(n_6580)
);

OAI22xp5_ASAP7_75t_L g6581 ( 
.A1(n_5538),
.A2(n_5394),
.B1(n_5282),
.B2(n_4678),
.Y(n_6581)
);

A2O1A1Ixp33_ASAP7_75t_L g6582 ( 
.A1(n_5394),
.A2(n_5353),
.B(n_5533),
.C(n_4639),
.Y(n_6582)
);

OR2x6_ASAP7_75t_L g6583 ( 
.A(n_4734),
.B(n_4754),
.Y(n_6583)
);

CKINVDCx5p33_ASAP7_75t_R g6584 ( 
.A(n_5319),
.Y(n_6584)
);

HB1xp67_ASAP7_75t_L g6585 ( 
.A(n_5331),
.Y(n_6585)
);

AOI22xp33_ASAP7_75t_L g6586 ( 
.A1(n_5647),
.A2(n_5691),
.B1(n_5688),
.B2(n_4579),
.Y(n_6586)
);

NAND2xp5_ASAP7_75t_SL g6587 ( 
.A(n_5394),
.B(n_4810),
.Y(n_6587)
);

BUFx4f_ASAP7_75t_L g6588 ( 
.A(n_5207),
.Y(n_6588)
);

NAND2xp5_ASAP7_75t_SL g6589 ( 
.A(n_5394),
.B(n_4810),
.Y(n_6589)
);

NAND2xp5_ASAP7_75t_SL g6590 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6590)
);

A2O1A1Ixp33_ASAP7_75t_L g6591 ( 
.A1(n_5533),
.A2(n_4639),
.B(n_4627),
.C(n_4734),
.Y(n_6591)
);

HB1xp67_ASAP7_75t_L g6592 ( 
.A(n_5371),
.Y(n_6592)
);

AOI21xp33_ASAP7_75t_L g6593 ( 
.A1(n_5267),
.A2(n_5430),
.B(n_5413),
.Y(n_6593)
);

AOI21xp5_ASAP7_75t_L g6594 ( 
.A1(n_5226),
.A2(n_5657),
.B(n_5650),
.Y(n_6594)
);

NAND2xp5_ASAP7_75t_L g6595 ( 
.A(n_4707),
.B(n_4712),
.Y(n_6595)
);

BUFx12f_ASAP7_75t_L g6596 ( 
.A(n_4736),
.Y(n_6596)
);

INVxp67_ASAP7_75t_L g6597 ( 
.A(n_5018),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_5004),
.B(n_5020),
.Y(n_6598)
);

INVx1_ASAP7_75t_SL g6599 ( 
.A(n_5020),
.Y(n_6599)
);

INVx1_ASAP7_75t_SL g6600 ( 
.A(n_5020),
.Y(n_6600)
);

CKINVDCx20_ASAP7_75t_R g6601 ( 
.A(n_4806),
.Y(n_6601)
);

CKINVDCx20_ASAP7_75t_R g6602 ( 
.A(n_4806),
.Y(n_6602)
);

A2O1A1Ixp33_ASAP7_75t_L g6603 ( 
.A1(n_4627),
.A2(n_4754),
.B(n_4765),
.C(n_4734),
.Y(n_6603)
);

AOI21xp5_ASAP7_75t_L g6604 ( 
.A1(n_5625),
.A2(n_5667),
.B(n_5660),
.Y(n_6604)
);

BUFx12f_ASAP7_75t_L g6605 ( 
.A(n_4762),
.Y(n_6605)
);

AOI21xp5_ASAP7_75t_L g6606 ( 
.A1(n_5660),
.A2(n_5711),
.B(n_5667),
.Y(n_6606)
);

NAND2x1p5_ASAP7_75t_L g6607 ( 
.A(n_5666),
.B(n_5715),
.Y(n_6607)
);

NOR2xp33_ASAP7_75t_L g6608 ( 
.A(n_5101),
.B(n_5408),
.Y(n_6608)
);

NOR2xp33_ASAP7_75t_L g6609 ( 
.A(n_5101),
.B(n_5408),
.Y(n_6609)
);

INVx2_ASAP7_75t_SL g6610 ( 
.A(n_4875),
.Y(n_6610)
);

AOI33xp33_ASAP7_75t_L g6611 ( 
.A1(n_5362),
.A2(n_5380),
.A3(n_5411),
.B1(n_5425),
.B2(n_5421),
.B3(n_5408),
.Y(n_6611)
);

O2A1O1Ixp33_ASAP7_75t_SL g6612 ( 
.A1(n_5444),
.A2(n_5118),
.B(n_5237),
.C(n_5077),
.Y(n_6612)
);

NAND2x1p5_ASAP7_75t_L g6613 ( 
.A(n_5666),
.B(n_5715),
.Y(n_6613)
);

NOR2xp33_ASAP7_75t_SL g6614 ( 
.A(n_5281),
.B(n_4571),
.Y(n_6614)
);

AOI21xp5_ASAP7_75t_L g6615 ( 
.A1(n_5711),
.A2(n_5693),
.B(n_5596),
.Y(n_6615)
);

OAI22xp5_ASAP7_75t_L g6616 ( 
.A1(n_4653),
.A2(n_4718),
.B1(n_4657),
.B2(n_4676),
.Y(n_6616)
);

NAND2xp5_ASAP7_75t_L g6617 ( 
.A(n_4712),
.B(n_4729),
.Y(n_6617)
);

AOI22xp5_ASAP7_75t_L g6618 ( 
.A1(n_5683),
.A2(n_5639),
.B1(n_5366),
.B2(n_5279),
.Y(n_6618)
);

BUFx2_ASAP7_75t_L g6619 ( 
.A(n_5502),
.Y(n_6619)
);

AOI21xp5_ASAP7_75t_L g6620 ( 
.A1(n_5596),
.A2(n_5693),
.B(n_5158),
.Y(n_6620)
);

A2O1A1Ixp33_ASAP7_75t_SL g6621 ( 
.A1(n_5576),
.A2(n_5583),
.B(n_5614),
.C(n_5611),
.Y(n_6621)
);

AND2x6_ASAP7_75t_SL g6622 ( 
.A(n_4910),
.B(n_5079),
.Y(n_6622)
);

BUFx2_ASAP7_75t_SL g6623 ( 
.A(n_5666),
.Y(n_6623)
);

OAI22xp5_ASAP7_75t_L g6624 ( 
.A1(n_4653),
.A2(n_4750),
.B1(n_4657),
.B2(n_4676),
.Y(n_6624)
);

NAND2xp5_ASAP7_75t_L g6625 ( 
.A(n_4729),
.B(n_4737),
.Y(n_6625)
);

OR2x6_ASAP7_75t_L g6626 ( 
.A(n_4754),
.B(n_4765),
.Y(n_6626)
);

AOI21xp5_ASAP7_75t_L g6627 ( 
.A1(n_5596),
.A2(n_5693),
.B(n_5158),
.Y(n_6627)
);

NOR2xp33_ASAP7_75t_L g6628 ( 
.A(n_5101),
.B(n_5411),
.Y(n_6628)
);

NOR2xp33_ASAP7_75t_L g6629 ( 
.A(n_5411),
.B(n_5421),
.Y(n_6629)
);

INVx4_ASAP7_75t_L g6630 ( 
.A(n_5715),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_4729),
.B(n_4737),
.Y(n_6631)
);

AOI21xp5_ASAP7_75t_L g6632 ( 
.A1(n_5596),
.A2(n_5693),
.B(n_5404),
.Y(n_6632)
);

INVx2_ASAP7_75t_SL g6633 ( 
.A(n_4875),
.Y(n_6633)
);

CKINVDCx8_ASAP7_75t_R g6634 ( 
.A(n_5715),
.Y(n_6634)
);

BUFx2_ASAP7_75t_L g6635 ( 
.A(n_5562),
.Y(n_6635)
);

BUFx2_ASAP7_75t_L g6636 ( 
.A(n_5562),
.Y(n_6636)
);

INVx2_ASAP7_75t_SL g6637 ( 
.A(n_4875),
.Y(n_6637)
);

OAI21xp33_ASAP7_75t_SL g6638 ( 
.A1(n_5183),
.A2(n_5426),
.B(n_5381),
.Y(n_6638)
);

NOR2xp33_ASAP7_75t_L g6639 ( 
.A(n_5421),
.B(n_5425),
.Y(n_6639)
);

INVx8_ASAP7_75t_L g6640 ( 
.A(n_5279),
.Y(n_6640)
);

NOR2xp33_ASAP7_75t_L g6641 ( 
.A(n_5425),
.B(n_5435),
.Y(n_6641)
);

OAI22xp5_ASAP7_75t_L g6642 ( 
.A1(n_4694),
.A2(n_4724),
.B1(n_4745),
.B2(n_4695),
.Y(n_6642)
);

OAI22xp5_ASAP7_75t_L g6643 ( 
.A1(n_4695),
.A2(n_4747),
.B1(n_4715),
.B2(n_4678),
.Y(n_6643)
);

NAND2xp5_ASAP7_75t_SL g6644 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6644)
);

BUFx2_ASAP7_75t_L g6645 ( 
.A(n_5562),
.Y(n_6645)
);

NOR2xp33_ASAP7_75t_L g6646 ( 
.A(n_5435),
.B(n_5448),
.Y(n_6646)
);

A2O1A1Ixp33_ASAP7_75t_L g6647 ( 
.A1(n_4754),
.A2(n_4765),
.B(n_5718),
.C(n_5022),
.Y(n_6647)
);

OR2x2_ASAP7_75t_L g6648 ( 
.A(n_4665),
.B(n_4688),
.Y(n_6648)
);

BUFx2_ASAP7_75t_L g6649 ( 
.A(n_5578),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_4737),
.B(n_4742),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_5216),
.Y(n_6651)
);

BUFx2_ASAP7_75t_L g6652 ( 
.A(n_5578),
.Y(n_6652)
);

INVx6_ASAP7_75t_L g6653 ( 
.A(n_4713),
.Y(n_6653)
);

AOI21xp5_ASAP7_75t_L g6654 ( 
.A1(n_5596),
.A2(n_5693),
.B(n_5404),
.Y(n_6654)
);

NAND2xp5_ASAP7_75t_L g6655 ( 
.A(n_4742),
.B(n_4743),
.Y(n_6655)
);

INVx2_ASAP7_75t_SL g6656 ( 
.A(n_4875),
.Y(n_6656)
);

INVx2_ASAP7_75t_SL g6657 ( 
.A(n_4875),
.Y(n_6657)
);

A2O1A1Ixp33_ASAP7_75t_L g6658 ( 
.A1(n_4765),
.A2(n_5718),
.B(n_5022),
.C(n_5026),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_5222),
.Y(n_6659)
);

O2A1O1Ixp33_ASAP7_75t_L g6660 ( 
.A1(n_5383),
.A2(n_5409),
.B(n_5410),
.C(n_5385),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_5222),
.Y(n_6661)
);

HB1xp67_ASAP7_75t_L g6662 ( 
.A(n_5385),
.Y(n_6662)
);

AOI21xp5_ASAP7_75t_L g6663 ( 
.A1(n_5401),
.A2(n_5404),
.B(n_5726),
.Y(n_6663)
);

INVx1_ASAP7_75t_SL g6664 ( 
.A(n_4633),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_5222),
.Y(n_6665)
);

O2A1O1Ixp33_ASAP7_75t_L g6666 ( 
.A1(n_5409),
.A2(n_5410),
.B(n_5450),
.C(n_5439),
.Y(n_6666)
);

AOI22xp5_ASAP7_75t_L g6667 ( 
.A1(n_5639),
.A2(n_5366),
.B1(n_5279),
.B2(n_5674),
.Y(n_6667)
);

BUFx2_ASAP7_75t_L g6668 ( 
.A(n_5578),
.Y(n_6668)
);

OR2x2_ASAP7_75t_L g6669 ( 
.A(n_4665),
.B(n_4688),
.Y(n_6669)
);

BUFx2_ASAP7_75t_L g6670 ( 
.A(n_5598),
.Y(n_6670)
);

HB1xp67_ASAP7_75t_L g6671 ( 
.A(n_5439),
.Y(n_6671)
);

INVx4_ASAP7_75t_L g6672 ( 
.A(n_5715),
.Y(n_6672)
);

NAND2xp5_ASAP7_75t_L g6673 ( 
.A(n_4742),
.B(n_4743),
.Y(n_6673)
);

O2A1O1Ixp33_ASAP7_75t_L g6674 ( 
.A1(n_5450),
.A2(n_5479),
.B(n_5413),
.C(n_5414),
.Y(n_6674)
);

NOR2x1_ASAP7_75t_L g6675 ( 
.A(n_4743),
.B(n_4744),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_SL g6676 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_5222),
.Y(n_6677)
);

INVx2_ASAP7_75t_SL g6678 ( 
.A(n_5051),
.Y(n_6678)
);

INVxp67_ASAP7_75t_L g6679 ( 
.A(n_5018),
.Y(n_6679)
);

AOI21xp5_ASAP7_75t_L g6680 ( 
.A1(n_5401),
.A2(n_5726),
.B(n_5715),
.Y(n_6680)
);

INVx1_ASAP7_75t_SL g6681 ( 
.A(n_4633),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_5251),
.Y(n_6682)
);

OAI22xp5_ASAP7_75t_L g6683 ( 
.A1(n_4718),
.A2(n_4745),
.B1(n_4730),
.B2(n_4694),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_5251),
.Y(n_6684)
);

INVxp67_ASAP7_75t_SL g6685 ( 
.A(n_5193),
.Y(n_6685)
);

CKINVDCx20_ASAP7_75t_R g6686 ( 
.A(n_5077),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_4744),
.B(n_4753),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_5251),
.Y(n_6688)
);

AOI21xp5_ASAP7_75t_L g6689 ( 
.A1(n_5401),
.A2(n_5726),
.B(n_5715),
.Y(n_6689)
);

NAND2xp5_ASAP7_75t_L g6690 ( 
.A(n_4744),
.B(n_4753),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_5286),
.Y(n_6691)
);

A2O1A1Ixp33_ASAP7_75t_L g6692 ( 
.A1(n_5026),
.A2(n_4500),
.B(n_4545),
.C(n_4512),
.Y(n_6692)
);

INVx3_ASAP7_75t_L g6693 ( 
.A(n_4495),
.Y(n_6693)
);

O2A1O1Ixp5_ASAP7_75t_L g6694 ( 
.A1(n_5607),
.A2(n_5653),
.B(n_5403),
.C(n_5430),
.Y(n_6694)
);

CKINVDCx20_ASAP7_75t_R g6695 ( 
.A(n_5118),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_5286),
.Y(n_6696)
);

NAND2xp5_ASAP7_75t_L g6697 ( 
.A(n_4753),
.B(n_4770),
.Y(n_6697)
);

A2O1A1Ixp33_ASAP7_75t_L g6698 ( 
.A1(n_4500),
.A2(n_4512),
.B(n_4545),
.C(n_4506),
.Y(n_6698)
);

INVxp67_ASAP7_75t_L g6699 ( 
.A(n_5479),
.Y(n_6699)
);

OR2x2_ASAP7_75t_L g6700 ( 
.A(n_4691),
.B(n_4700),
.Y(n_6700)
);

AOI21xp5_ASAP7_75t_L g6701 ( 
.A1(n_5726),
.A2(n_5715),
.B(n_5354),
.Y(n_6701)
);

O2A1O1Ixp33_ASAP7_75t_L g6702 ( 
.A1(n_5403),
.A2(n_5420),
.B(n_5414),
.C(n_5601),
.Y(n_6702)
);

NAND2xp5_ASAP7_75t_L g6703 ( 
.A(n_4770),
.B(n_4773),
.Y(n_6703)
);

INVx3_ASAP7_75t_L g6704 ( 
.A(n_4495),
.Y(n_6704)
);

NAND2xp5_ASAP7_75t_SL g6705 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6705)
);

INVx3_ASAP7_75t_L g6706 ( 
.A(n_4495),
.Y(n_6706)
);

AOI21xp5_ASAP7_75t_L g6707 ( 
.A1(n_5726),
.A2(n_5715),
.B(n_5354),
.Y(n_6707)
);

AND3x1_ASAP7_75t_SL g6708 ( 
.A(n_5510),
.B(n_5665),
.C(n_4910),
.Y(n_6708)
);

INVx2_ASAP7_75t_SL g6709 ( 
.A(n_5051),
.Y(n_6709)
);

AOI22xp5_ASAP7_75t_L g6710 ( 
.A1(n_5279),
.A2(n_5366),
.B1(n_5674),
.B2(n_5558),
.Y(n_6710)
);

INVx2_ASAP7_75t_SL g6711 ( 
.A(n_5051),
.Y(n_6711)
);

O2A1O1Ixp33_ASAP7_75t_L g6712 ( 
.A1(n_5420),
.A2(n_5601),
.B(n_5647),
.C(n_4886),
.Y(n_6712)
);

AOI21xp5_ASAP7_75t_L g6713 ( 
.A1(n_5726),
.A2(n_5354),
.B(n_5320),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_5286),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_5286),
.Y(n_6715)
);

NAND2xp5_ASAP7_75t_L g6716 ( 
.A(n_4770),
.B(n_4773),
.Y(n_6716)
);

AOI22xp33_ASAP7_75t_L g6717 ( 
.A1(n_5691),
.A2(n_4579),
.B1(n_4587),
.B2(n_4571),
.Y(n_6717)
);

OAI22xp5_ASAP7_75t_L g6718 ( 
.A1(n_4732),
.A2(n_4735),
.B1(n_4700),
.B2(n_4708),
.Y(n_6718)
);

AOI22xp33_ASAP7_75t_L g6719 ( 
.A1(n_4571),
.A2(n_4587),
.B1(n_4598),
.B2(n_4579),
.Y(n_6719)
);

NAND2x1p5_ASAP7_75t_L g6720 ( 
.A(n_5726),
.B(n_4571),
.Y(n_6720)
);

OA22x2_ASAP7_75t_L g6721 ( 
.A1(n_4486),
.A2(n_4522),
.B1(n_4528),
.B2(n_4505),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_5318),
.Y(n_6722)
);

INVx2_ASAP7_75t_L g6723 ( 
.A(n_5318),
.Y(n_6723)
);

AOI21xp5_ASAP7_75t_L g6724 ( 
.A1(n_5320),
.A2(n_5405),
.B(n_5354),
.Y(n_6724)
);

A2O1A1Ixp33_ASAP7_75t_L g6725 ( 
.A1(n_4500),
.A2(n_4512),
.B(n_4545),
.C(n_4506),
.Y(n_6725)
);

AOI21xp5_ASAP7_75t_L g6726 ( 
.A1(n_5320),
.A2(n_5405),
.B(n_5354),
.Y(n_6726)
);

NAND2xp5_ASAP7_75t_L g6727 ( 
.A(n_4773),
.B(n_4776),
.Y(n_6727)
);

AOI222xp33_ASAP7_75t_L g6728 ( 
.A1(n_5607),
.A2(n_4537),
.B1(n_5575),
.B2(n_5134),
.C1(n_5133),
.C2(n_5707),
.Y(n_6728)
);

BUFx2_ASAP7_75t_L g6729 ( 
.A(n_5598),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_5318),
.Y(n_6730)
);

AOI22xp5_ASAP7_75t_L g6731 ( 
.A1(n_5366),
.A2(n_5558),
.B1(n_5585),
.B2(n_5555),
.Y(n_6731)
);

AOI21xp33_ASAP7_75t_L g6732 ( 
.A1(n_5267),
.A2(n_5579),
.B(n_5219),
.Y(n_6732)
);

AOI22x1_ASAP7_75t_L g6733 ( 
.A1(n_4537),
.A2(n_5496),
.B1(n_5539),
.B2(n_5486),
.Y(n_6733)
);

AOI21xp5_ASAP7_75t_L g6734 ( 
.A1(n_5320),
.A2(n_5417),
.B(n_5405),
.Y(n_6734)
);

A2O1A1Ixp33_ASAP7_75t_L g6735 ( 
.A1(n_4500),
.A2(n_4512),
.B(n_4545),
.C(n_4506),
.Y(n_6735)
);

A2O1A1Ixp33_ASAP7_75t_L g6736 ( 
.A1(n_4506),
.A2(n_4551),
.B(n_4575),
.C(n_4550),
.Y(n_6736)
);

NOR2xp67_ASAP7_75t_L g6737 ( 
.A(n_5267),
.B(n_5193),
.Y(n_6737)
);

AOI21xp5_ASAP7_75t_L g6738 ( 
.A1(n_5320),
.A2(n_5417),
.B(n_5405),
.Y(n_6738)
);

HB1xp67_ASAP7_75t_L g6739 ( 
.A(n_4850),
.Y(n_6739)
);

NAND2xp5_ASAP7_75t_L g6740 ( 
.A(n_4776),
.B(n_4782),
.Y(n_6740)
);

CKINVDCx5p33_ASAP7_75t_R g6741 ( 
.A(n_5389),
.Y(n_6741)
);

CKINVDCx5p33_ASAP7_75t_R g6742 ( 
.A(n_5389),
.Y(n_6742)
);

OAI22xp5_ASAP7_75t_L g6743 ( 
.A1(n_4730),
.A2(n_4732),
.B1(n_4708),
.B2(n_4715),
.Y(n_6743)
);

AOI22xp5_ASAP7_75t_L g6744 ( 
.A1(n_5366),
.A2(n_5558),
.B1(n_5585),
.B2(n_5555),
.Y(n_6744)
);

AOI22xp5_ASAP7_75t_L g6745 ( 
.A1(n_5366),
.A2(n_5585),
.B1(n_5616),
.B2(n_5555),
.Y(n_6745)
);

INVx2_ASAP7_75t_L g6746 ( 
.A(n_5396),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_4534),
.Y(n_6747)
);

NOR2xp33_ASAP7_75t_L g6748 ( 
.A(n_5435),
.B(n_5448),
.Y(n_6748)
);

INVxp67_ASAP7_75t_SL g6749 ( 
.A(n_5219),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_5396),
.Y(n_6750)
);

NAND2xp5_ASAP7_75t_L g6751 ( 
.A(n_4776),
.B(n_4782),
.Y(n_6751)
);

HB1xp67_ASAP7_75t_L g6752 ( 
.A(n_4850),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_4534),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_4534),
.Y(n_6754)
);

OAI22xp5_ASAP7_75t_L g6755 ( 
.A1(n_4738),
.A2(n_4724),
.B1(n_4725),
.B2(n_4691),
.Y(n_6755)
);

NAND2xp5_ASAP7_75t_SL g6756 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6756)
);

O2A1O1Ixp33_ASAP7_75t_L g6757 ( 
.A1(n_4728),
.A2(n_5006),
.B(n_5428),
.C(n_4886),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_SL g6758 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6758)
);

AOI22xp33_ASAP7_75t_L g6759 ( 
.A1(n_4571),
.A2(n_4587),
.B1(n_4598),
.B2(n_4579),
.Y(n_6759)
);

AOI22xp33_ASAP7_75t_L g6760 ( 
.A1(n_4579),
.A2(n_4598),
.B1(n_4626),
.B2(n_4587),
.Y(n_6760)
);

NOR2xp33_ASAP7_75t_R g6761 ( 
.A(n_5237),
.B(n_5274),
.Y(n_6761)
);

INVx4_ASAP7_75t_L g6762 ( 
.A(n_4772),
.Y(n_6762)
);

NOR2xp33_ASAP7_75t_L g6763 ( 
.A(n_5448),
.B(n_5449),
.Y(n_6763)
);

OAI22xp5_ASAP7_75t_SL g6764 ( 
.A1(n_5444),
.A2(n_5274),
.B1(n_5575),
.B2(n_5687),
.Y(n_6764)
);

A2O1A1Ixp33_ASAP7_75t_L g6765 ( 
.A1(n_4551),
.A2(n_4575),
.B(n_4583),
.C(n_4550),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_5396),
.Y(n_6766)
);

BUFx6f_ASAP7_75t_SL g6767 ( 
.A(n_4587),
.Y(n_6767)
);

AOI21xp5_ASAP7_75t_L g6768 ( 
.A1(n_5405),
.A2(n_5417),
.B(n_5581),
.Y(n_6768)
);

INVx2_ASAP7_75t_L g6769 ( 
.A(n_5396),
.Y(n_6769)
);

NOR2x1_ASAP7_75t_L g6770 ( 
.A(n_4782),
.B(n_4783),
.Y(n_6770)
);

AOI21xp5_ASAP7_75t_L g6771 ( 
.A1(n_5417),
.A2(n_5586),
.B(n_5581),
.Y(n_6771)
);

OAI22xp5_ASAP7_75t_L g6772 ( 
.A1(n_4735),
.A2(n_4738),
.B1(n_4747),
.B2(n_4725),
.Y(n_6772)
);

INVxp67_ASAP7_75t_L g6773 ( 
.A(n_5340),
.Y(n_6773)
);

INVx2_ASAP7_75t_SL g6774 ( 
.A(n_5051),
.Y(n_6774)
);

OR2x6_ASAP7_75t_L g6775 ( 
.A(n_4587),
.B(n_4598),
.Y(n_6775)
);

NAND2xp5_ASAP7_75t_L g6776 ( 
.A(n_4783),
.B(n_4786),
.Y(n_6776)
);

NOR2x1_ASAP7_75t_L g6777 ( 
.A(n_4783),
.B(n_4786),
.Y(n_6777)
);

BUFx12f_ASAP7_75t_L g6778 ( 
.A(n_4762),
.Y(n_6778)
);

NAND2xp5_ASAP7_75t_SL g6779 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6779)
);

BUFx2_ASAP7_75t_L g6780 ( 
.A(n_5598),
.Y(n_6780)
);

AOI21x1_ASAP7_75t_L g6781 ( 
.A1(n_5223),
.A2(n_5227),
.B(n_5579),
.Y(n_6781)
);

BUFx2_ASAP7_75t_L g6782 ( 
.A(n_5645),
.Y(n_6782)
);

OAI22xp5_ASAP7_75t_L g6783 ( 
.A1(n_4748),
.A2(n_4626),
.B1(n_4668),
.B2(n_4598),
.Y(n_6783)
);

NAND2xp5_ASAP7_75t_L g6784 ( 
.A(n_4786),
.B(n_4794),
.Y(n_6784)
);

CKINVDCx14_ASAP7_75t_R g6785 ( 
.A(n_5463),
.Y(n_6785)
);

AOI22xp33_ASAP7_75t_L g6786 ( 
.A1(n_4598),
.A2(n_4668),
.B1(n_4849),
.B2(n_4626),
.Y(n_6786)
);

NAND2xp5_ASAP7_75t_SL g6787 ( 
.A(n_5512),
.B(n_5513),
.Y(n_6787)
);

O2A1O1Ixp33_ASAP7_75t_L g6788 ( 
.A1(n_4728),
.A2(n_5006),
.B(n_5428),
.C(n_4886),
.Y(n_6788)
);

O2A1O1Ixp5_ASAP7_75t_SL g6789 ( 
.A1(n_5223),
.A2(n_5227),
.B(n_5192),
.C(n_5202),
.Y(n_6789)
);

INVx3_ASAP7_75t_L g6790 ( 
.A(n_4495),
.Y(n_6790)
);

OR2x2_ASAP7_75t_L g6791 ( 
.A(n_4748),
.B(n_4763),
.Y(n_6791)
);

NAND2xp5_ASAP7_75t_L g6792 ( 
.A(n_4794),
.B(n_4796),
.Y(n_6792)
);

AOI21xp5_ASAP7_75t_L g6793 ( 
.A1(n_5417),
.A2(n_5586),
.B(n_5581),
.Y(n_6793)
);

CKINVDCx6p67_ASAP7_75t_R g6794 ( 
.A(n_4521),
.Y(n_6794)
);

OAI22xp5_ASAP7_75t_L g6795 ( 
.A1(n_4626),
.A2(n_4668),
.B1(n_4860),
.B2(n_4849),
.Y(n_6795)
);

NOR2xp33_ASAP7_75t_L g6796 ( 
.A(n_5449),
.B(n_5452),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_L g6797 ( 
.A(n_4794),
.B(n_4796),
.Y(n_6797)
);

INVxp67_ASAP7_75t_L g6798 ( 
.A(n_5340),
.Y(n_6798)
);

NAND2xp5_ASAP7_75t_L g6799 ( 
.A(n_4796),
.B(n_4798),
.Y(n_6799)
);

HB1xp67_ASAP7_75t_L g6800 ( 
.A(n_4912),
.Y(n_6800)
);

CKINVDCx20_ASAP7_75t_R g6801 ( 
.A(n_4846),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_SL g6802 ( 
.A(n_5643),
.B(n_5617),
.Y(n_6802)
);

NOR2xp33_ASAP7_75t_R g6803 ( 
.A(n_5463),
.B(n_5471),
.Y(n_6803)
);

BUFx3_ASAP7_75t_L g6804 ( 
.A(n_4478),
.Y(n_6804)
);

CKINVDCx5p33_ASAP7_75t_R g6805 ( 
.A(n_5436),
.Y(n_6805)
);

AOI21xp5_ASAP7_75t_L g6806 ( 
.A1(n_5586),
.A2(n_5656),
.B(n_5651),
.Y(n_6806)
);

BUFx3_ASAP7_75t_L g6807 ( 
.A(n_4478),
.Y(n_6807)
);

INVxp67_ASAP7_75t_L g6808 ( 
.A(n_5340),
.Y(n_6808)
);

HB1xp67_ASAP7_75t_L g6809 ( 
.A(n_4912),
.Y(n_6809)
);

AOI22xp5_ASAP7_75t_L g6810 ( 
.A1(n_5585),
.A2(n_5616),
.B1(n_5607),
.B2(n_4521),
.Y(n_6810)
);

NAND2xp5_ASAP7_75t_L g6811 ( 
.A(n_4798),
.B(n_4800),
.Y(n_6811)
);

BUFx8_ASAP7_75t_L g6812 ( 
.A(n_4772),
.Y(n_6812)
);

AOI21xp5_ASAP7_75t_L g6813 ( 
.A1(n_5651),
.A2(n_5656),
.B(n_5381),
.Y(n_6813)
);

AOI21xp5_ASAP7_75t_L g6814 ( 
.A1(n_5651),
.A2(n_5656),
.B(n_5381),
.Y(n_6814)
);

NOR2xp33_ASAP7_75t_L g6815 ( 
.A(n_5449),
.B(n_5452),
.Y(n_6815)
);

INVx4_ASAP7_75t_L g6816 ( 
.A(n_4772),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_4798),
.B(n_4800),
.Y(n_6817)
);

AOI22xp5_ASAP7_75t_L g6818 ( 
.A1(n_5616),
.A2(n_4559),
.B1(n_5191),
.B2(n_4608),
.Y(n_6818)
);

O2A1O1Ixp33_ASAP7_75t_L g6819 ( 
.A1(n_4728),
.A2(n_5006),
.B(n_5428),
.C(n_4886),
.Y(n_6819)
);

OAI22xp5_ASAP7_75t_L g6820 ( 
.A1(n_4626),
.A2(n_4668),
.B1(n_4860),
.B2(n_4849),
.Y(n_6820)
);

AOI21xp5_ASAP7_75t_L g6821 ( 
.A1(n_5183),
.A2(n_5469),
.B(n_5426),
.Y(n_6821)
);

OAI22xp33_ASAP7_75t_L g6822 ( 
.A1(n_4668),
.A2(n_4860),
.B1(n_4868),
.B2(n_4849),
.Y(n_6822)
);

NAND2xp5_ASAP7_75t_L g6823 ( 
.A(n_4800),
.B(n_4804),
.Y(n_6823)
);

BUFx3_ASAP7_75t_L g6824 ( 
.A(n_4478),
.Y(n_6824)
);

INVxp67_ASAP7_75t_SL g6825 ( 
.A(n_5290),
.Y(n_6825)
);

NAND2xp5_ASAP7_75t_SL g6826 ( 
.A(n_5643),
.B(n_5617),
.Y(n_6826)
);

BUFx3_ASAP7_75t_L g6827 ( 
.A(n_4478),
.Y(n_6827)
);

NAND2xp5_ASAP7_75t_L g6828 ( 
.A(n_4804),
.B(n_4808),
.Y(n_6828)
);

A2O1A1Ixp33_ASAP7_75t_L g6829 ( 
.A1(n_4550),
.A2(n_4575),
.B(n_4583),
.C(n_4551),
.Y(n_6829)
);

CKINVDCx20_ASAP7_75t_R g6830 ( 
.A(n_4846),
.Y(n_6830)
);

AOI21xp5_ASAP7_75t_L g6831 ( 
.A1(n_5183),
.A2(n_5469),
.B(n_5426),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_4804),
.B(n_4808),
.Y(n_6832)
);

NOR2xp33_ASAP7_75t_L g6833 ( 
.A(n_5452),
.B(n_5457),
.Y(n_6833)
);

AOI21xp33_ASAP7_75t_L g6834 ( 
.A1(n_5579),
.A2(n_5400),
.B(n_5593),
.Y(n_6834)
);

NAND2xp5_ASAP7_75t_L g6835 ( 
.A(n_4808),
.B(n_4815),
.Y(n_6835)
);

HB1xp67_ASAP7_75t_L g6836 ( 
.A(n_4955),
.Y(n_6836)
);

BUFx4f_ASAP7_75t_L g6837 ( 
.A(n_4772),
.Y(n_6837)
);

HB1xp67_ASAP7_75t_L g6838 ( 
.A(n_4955),
.Y(n_6838)
);

NOR2xp33_ASAP7_75t_L g6839 ( 
.A(n_5457),
.B(n_5462),
.Y(n_6839)
);

INVx1_ASAP7_75t_SL g6840 ( 
.A(n_4633),
.Y(n_6840)
);

AOI22xp33_ASAP7_75t_L g6841 ( 
.A1(n_4849),
.A2(n_4868),
.B1(n_4899),
.B2(n_4860),
.Y(n_6841)
);

NOR2xp33_ASAP7_75t_L g6842 ( 
.A(n_5457),
.B(n_5462),
.Y(n_6842)
);

AOI21xp5_ASAP7_75t_L g6843 ( 
.A1(n_5469),
.A2(n_5529),
.B(n_4886),
.Y(n_6843)
);

NOR2xp33_ASAP7_75t_L g6844 ( 
.A(n_5462),
.B(n_5470),
.Y(n_6844)
);

AOI21xp5_ASAP7_75t_L g6845 ( 
.A1(n_5529),
.A2(n_5006),
.B(n_4728),
.Y(n_6845)
);

HB1xp67_ASAP7_75t_L g6846 ( 
.A(n_5013),
.Y(n_6846)
);

O2A1O1Ixp33_ASAP7_75t_L g6847 ( 
.A1(n_4728),
.A2(n_5428),
.B(n_5006),
.C(n_5269),
.Y(n_6847)
);

NAND2xp5_ASAP7_75t_SL g6848 ( 
.A(n_5643),
.B(n_5617),
.Y(n_6848)
);

INVx1_ASAP7_75t_SL g6849 ( 
.A(n_5264),
.Y(n_6849)
);

INVx1_ASAP7_75t_SL g6850 ( 
.A(n_5264),
.Y(n_6850)
);

BUFx3_ASAP7_75t_L g6851 ( 
.A(n_4478),
.Y(n_6851)
);

OAI22xp5_ASAP7_75t_L g6852 ( 
.A1(n_4860),
.A2(n_4899),
.B1(n_4901),
.B2(n_4868),
.Y(n_6852)
);

NAND2xp5_ASAP7_75t_L g6853 ( 
.A(n_4815),
.B(n_4823),
.Y(n_6853)
);

NOR2xp33_ASAP7_75t_L g6854 ( 
.A(n_5470),
.B(n_5476),
.Y(n_6854)
);

NAND2x2_ASAP7_75t_L g6855 ( 
.A(n_4722),
.B(n_5627),
.Y(n_6855)
);

HB1xp67_ASAP7_75t_L g6856 ( 
.A(n_5013),
.Y(n_6856)
);

AND2x4_ASAP7_75t_L g6857 ( 
.A(n_4722),
.B(n_4486),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_SL g6858 ( 
.A(n_5617),
.B(n_5623),
.Y(n_6858)
);

AOI21xp5_ASAP7_75t_L g6859 ( 
.A1(n_5529),
.A2(n_5428),
.B(n_5645),
.Y(n_6859)
);

AOI22xp5_ASAP7_75t_L g6860 ( 
.A1(n_5616),
.A2(n_4559),
.B1(n_5233),
.B2(n_5191),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_4815),
.B(n_4823),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_SL g6862 ( 
.A(n_5623),
.B(n_5023),
.Y(n_6862)
);

INVx2_ASAP7_75t_SL g6863 ( 
.A(n_5051),
.Y(n_6863)
);

AOI21xp5_ASAP7_75t_L g6864 ( 
.A1(n_5645),
.A2(n_5161),
.B(n_5154),
.Y(n_6864)
);

AOI22xp33_ASAP7_75t_L g6865 ( 
.A1(n_4868),
.A2(n_4901),
.B1(n_4964),
.B2(n_4899),
.Y(n_6865)
);

AOI22xp5_ASAP7_75t_L g6866 ( 
.A1(n_4559),
.A2(n_4608),
.B1(n_5233),
.B2(n_5191),
.Y(n_6866)
);

NOR2xp33_ASAP7_75t_L g6867 ( 
.A(n_5470),
.B(n_5476),
.Y(n_6867)
);

BUFx3_ASAP7_75t_L g6868 ( 
.A(n_4478),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_4823),
.B(n_4826),
.Y(n_6869)
);

BUFx2_ASAP7_75t_L g6870 ( 
.A(n_4689),
.Y(n_6870)
);

NAND2xp33_ASAP7_75t_L g6871 ( 
.A(n_4772),
.B(n_4814),
.Y(n_6871)
);

AOI21x1_ASAP7_75t_L g6872 ( 
.A1(n_5290),
.A2(n_5298),
.B(n_5294),
.Y(n_6872)
);

NAND2xp5_ASAP7_75t_L g6873 ( 
.A(n_4826),
.B(n_4834),
.Y(n_6873)
);

NOR3xp33_ASAP7_75t_L g6874 ( 
.A(n_5345),
.B(n_5269),
.C(n_5270),
.Y(n_6874)
);

BUFx3_ASAP7_75t_L g6875 ( 
.A(n_4478),
.Y(n_6875)
);

BUFx12f_ASAP7_75t_L g6876 ( 
.A(n_4866),
.Y(n_6876)
);

AOI21xp5_ASAP7_75t_L g6877 ( 
.A1(n_5154),
.A2(n_5161),
.B(n_5290),
.Y(n_6877)
);

AOI22xp5_ASAP7_75t_L g6878 ( 
.A1(n_4559),
.A2(n_4608),
.B1(n_5191),
.B2(n_5233),
.Y(n_6878)
);

NAND2xp5_ASAP7_75t_L g6879 ( 
.A(n_4826),
.B(n_4834),
.Y(n_6879)
);

CKINVDCx20_ASAP7_75t_R g6880 ( 
.A(n_4866),
.Y(n_6880)
);

CKINVDCx16_ASAP7_75t_R g6881 ( 
.A(n_4608),
.Y(n_6881)
);

INVxp67_ASAP7_75t_SL g6882 ( 
.A(n_5294),
.Y(n_6882)
);

CKINVDCx5p33_ASAP7_75t_R g6883 ( 
.A(n_5436),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_4834),
.B(n_4838),
.Y(n_6884)
);

AOI22xp33_ASAP7_75t_L g6885 ( 
.A1(n_4868),
.A2(n_4901),
.B1(n_4964),
.B2(n_4899),
.Y(n_6885)
);

CKINVDCx5p33_ASAP7_75t_R g6886 ( 
.A(n_4880),
.Y(n_6886)
);

OAI22xp5_ASAP7_75t_L g6887 ( 
.A1(n_4899),
.A2(n_4964),
.B1(n_4965),
.B2(n_4901),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_SL g6888 ( 
.A(n_5623),
.B(n_5023),
.Y(n_6888)
);

O2A1O1Ixp33_ASAP7_75t_L g6889 ( 
.A1(n_5270),
.A2(n_5280),
.B(n_5283),
.C(n_5277),
.Y(n_6889)
);

BUFx2_ASAP7_75t_L g6890 ( 
.A(n_4689),
.Y(n_6890)
);

INVx2_ASAP7_75t_SL g6891 ( 
.A(n_5051),
.Y(n_6891)
);

NAND2xp5_ASAP7_75t_L g6892 ( 
.A(n_4838),
.B(n_4839),
.Y(n_6892)
);

INVx6_ASAP7_75t_SL g6893 ( 
.A(n_5716),
.Y(n_6893)
);

OAI321xp33_ASAP7_75t_L g6894 ( 
.A1(n_4557),
.A2(n_4561),
.A3(n_5600),
.B1(n_5606),
.B2(n_5595),
.C(n_5593),
.Y(n_6894)
);

CKINVDCx16_ASAP7_75t_R g6895 ( 
.A(n_5233),
.Y(n_6895)
);

AOI21xp5_ASAP7_75t_L g6896 ( 
.A1(n_5154),
.A2(n_5161),
.B(n_5294),
.Y(n_6896)
);

NAND2x1p5_ASAP7_75t_L g6897 ( 
.A(n_4964),
.B(n_4965),
.Y(n_6897)
);

INVx4_ASAP7_75t_L g6898 ( 
.A(n_4772),
.Y(n_6898)
);

INVxp67_ASAP7_75t_SL g6899 ( 
.A(n_5298),
.Y(n_6899)
);

BUFx3_ASAP7_75t_L g6900 ( 
.A(n_4478),
.Y(n_6900)
);

CKINVDCx16_ASAP7_75t_R g6901 ( 
.A(n_5349),
.Y(n_6901)
);

INVx4_ASAP7_75t_L g6902 ( 
.A(n_4814),
.Y(n_6902)
);

INVx3_ASAP7_75t_L g6903 ( 
.A(n_4516),
.Y(n_6903)
);

OAI22xp5_ASAP7_75t_L g6904 ( 
.A1(n_4965),
.A2(n_5687),
.B1(n_4814),
.B2(n_4788),
.Y(n_6904)
);

NAND2xp5_ASAP7_75t_SL g6905 ( 
.A(n_5623),
.B(n_5062),
.Y(n_6905)
);

BUFx2_ASAP7_75t_L g6906 ( 
.A(n_4689),
.Y(n_6906)
);

AOI21xp5_ASAP7_75t_L g6907 ( 
.A1(n_5298),
.A2(n_5299),
.B(n_5350),
.Y(n_6907)
);

BUFx2_ASAP7_75t_L g6908 ( 
.A(n_4711),
.Y(n_6908)
);

AOI21xp5_ASAP7_75t_L g6909 ( 
.A1(n_5299),
.A2(n_5373),
.B(n_5350),
.Y(n_6909)
);

NOR2xp33_ASAP7_75t_R g6910 ( 
.A(n_5471),
.B(n_5349),
.Y(n_6910)
);

INVx2_ASAP7_75t_SL g6911 ( 
.A(n_5051),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_SL g6912 ( 
.A(n_5062),
.B(n_5068),
.Y(n_6912)
);

OAI22xp5_ASAP7_75t_L g6913 ( 
.A1(n_4965),
.A2(n_5687),
.B1(n_4814),
.B2(n_4763),
.Y(n_6913)
);

BUFx3_ASAP7_75t_L g6914 ( 
.A(n_4478),
.Y(n_6914)
);

AOI21xp5_ASAP7_75t_L g6915 ( 
.A1(n_5299),
.A2(n_5373),
.B(n_5350),
.Y(n_6915)
);

BUFx2_ASAP7_75t_L g6916 ( 
.A(n_4711),
.Y(n_6916)
);

NAND2xp5_ASAP7_75t_L g6917 ( 
.A(n_4838),
.B(n_4839),
.Y(n_6917)
);

NAND2xp5_ASAP7_75t_SL g6918 ( 
.A(n_5062),
.B(n_5068),
.Y(n_6918)
);

O2A1O1Ixp33_ASAP7_75t_L g6919 ( 
.A1(n_5277),
.A2(n_5283),
.B(n_5285),
.C(n_5280),
.Y(n_6919)
);

A2O1A1Ixp33_ASAP7_75t_SL g6920 ( 
.A1(n_5576),
.A2(n_5583),
.B(n_5614),
.C(n_5611),
.Y(n_6920)
);

OAI21xp33_ASAP7_75t_SL g6921 ( 
.A1(n_5574),
.A2(n_4788),
.B(n_4763),
.Y(n_6921)
);

OR2x2_ASAP7_75t_L g6922 ( 
.A(n_4788),
.B(n_4790),
.Y(n_6922)
);

AOI22xp5_ASAP7_75t_L g6923 ( 
.A1(n_5900),
.A2(n_4965),
.B1(n_4660),
.B2(n_4666),
.Y(n_6923)
);

INVx3_ASAP7_75t_L g6924 ( 
.A(n_5732),
.Y(n_6924)
);

A2O1A1Ixp33_ASAP7_75t_L g6925 ( 
.A1(n_5946),
.A2(n_4551),
.B(n_4575),
.C(n_4550),
.Y(n_6925)
);

BUFx6f_ASAP7_75t_L g6926 ( 
.A(n_6467),
.Y(n_6926)
);

AOI22xp5_ASAP7_75t_L g6927 ( 
.A1(n_5900),
.A2(n_4660),
.B1(n_4666),
.B2(n_4478),
.Y(n_6927)
);

CKINVDCx5p33_ASAP7_75t_R g6928 ( 
.A(n_6134),
.Y(n_6928)
);

INVx2_ASAP7_75t_L g6929 ( 
.A(n_6722),
.Y(n_6929)
);

BUFx8_ASAP7_75t_SL g6930 ( 
.A(n_6402),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_6722),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6651),
.Y(n_6932)
);

AOI22xp5_ASAP7_75t_L g6933 ( 
.A1(n_5983),
.A2(n_4660),
.B1(n_4666),
.B2(n_4478),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6651),
.Y(n_6934)
);

INVx2_ASAP7_75t_SL g6935 ( 
.A(n_6855),
.Y(n_6935)
);

INVx1_ASAP7_75t_L g6936 ( 
.A(n_6659),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6659),
.Y(n_6937)
);

NAND2xp5_ASAP7_75t_L g6938 ( 
.A(n_5979),
.B(n_6209),
.Y(n_6938)
);

NAND2xp5_ASAP7_75t_L g6939 ( 
.A(n_5979),
.B(n_6209),
.Y(n_6939)
);

INVx3_ASAP7_75t_L g6940 ( 
.A(n_5732),
.Y(n_6940)
);

CKINVDCx11_ASAP7_75t_R g6941 ( 
.A(n_6134),
.Y(n_6941)
);

BUFx3_ASAP7_75t_L g6942 ( 
.A(n_6804),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6661),
.Y(n_6943)
);

INVx2_ASAP7_75t_L g6944 ( 
.A(n_6722),
.Y(n_6944)
);

OR2x6_ASAP7_75t_L g6945 ( 
.A(n_6368),
.B(n_5689),
.Y(n_6945)
);

AND2x2_ASAP7_75t_L g6946 ( 
.A(n_6044),
.B(n_5248),
.Y(n_6946)
);

BUFx3_ASAP7_75t_L g6947 ( 
.A(n_6804),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_5728),
.B(n_4839),
.Y(n_6948)
);

BUFx6f_ASAP7_75t_L g6949 ( 
.A(n_6467),
.Y(n_6949)
);

INVx2_ASAP7_75t_L g6950 ( 
.A(n_6722),
.Y(n_6950)
);

CKINVDCx5p33_ASAP7_75t_R g6951 ( 
.A(n_6318),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6723),
.Y(n_6952)
);

INVx3_ASAP7_75t_L g6953 ( 
.A(n_5732),
.Y(n_6953)
);

NAND2x1p5_ASAP7_75t_L g6954 ( 
.A(n_6224),
.B(n_5676),
.Y(n_6954)
);

BUFx6f_ASAP7_75t_L g6955 ( 
.A(n_6467),
.Y(n_6955)
);

CKINVDCx5p33_ASAP7_75t_R g6956 ( 
.A(n_6318),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6661),
.Y(n_6957)
);

AO32x2_ASAP7_75t_L g6958 ( 
.A1(n_6616),
.A2(n_4840),
.A3(n_4818),
.B1(n_4790),
.B2(n_5068),
.Y(n_6958)
);

INVx3_ASAP7_75t_L g6959 ( 
.A(n_5732),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6665),
.Y(n_6960)
);

NAND2xp5_ASAP7_75t_L g6961 ( 
.A(n_5728),
.B(n_4842),
.Y(n_6961)
);

AOI22xp33_ASAP7_75t_L g6962 ( 
.A1(n_5951),
.A2(n_4814),
.B1(n_5349),
.B2(n_5725),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_5801),
.B(n_4842),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6665),
.Y(n_6964)
);

INVx8_ASAP7_75t_L g6965 ( 
.A(n_6179),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6677),
.Y(n_6966)
);

INVx3_ASAP7_75t_L g6967 ( 
.A(n_5732),
.Y(n_6967)
);

AOI22xp5_ASAP7_75t_L g6968 ( 
.A1(n_5983),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_5801),
.B(n_4842),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6677),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6684),
.Y(n_6971)
);

NAND2x1p5_ASAP7_75t_L g6972 ( 
.A(n_6224),
.B(n_5676),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6684),
.Y(n_6973)
);

NAND2xp5_ASAP7_75t_L g6974 ( 
.A(n_6315),
.B(n_4854),
.Y(n_6974)
);

OR2x6_ASAP7_75t_SL g6975 ( 
.A(n_6158),
.B(n_5133),
.Y(n_6975)
);

BUFx6f_ASAP7_75t_L g6976 ( 
.A(n_6283),
.Y(n_6976)
);

HB1xp67_ASAP7_75t_L g6977 ( 
.A(n_5817),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6688),
.Y(n_6978)
);

AND2x2_ASAP7_75t_L g6979 ( 
.A(n_6044),
.B(n_5248),
.Y(n_6979)
);

CKINVDCx5p33_ASAP7_75t_R g6980 ( 
.A(n_5926),
.Y(n_6980)
);

AND2x2_ASAP7_75t_L g6981 ( 
.A(n_6044),
.B(n_5256),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6688),
.Y(n_6982)
);

BUFx3_ASAP7_75t_L g6983 ( 
.A(n_6804),
.Y(n_6983)
);

AOI21xp33_ASAP7_75t_L g6984 ( 
.A1(n_5894),
.A2(n_5177),
.B(n_5167),
.Y(n_6984)
);

NAND2xp5_ASAP7_75t_L g6985 ( 
.A(n_6315),
.B(n_6077),
.Y(n_6985)
);

AND2x2_ASAP7_75t_L g6986 ( 
.A(n_6093),
.B(n_5256),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6691),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_6723),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6691),
.Y(n_6989)
);

INVxp67_ASAP7_75t_L g6990 ( 
.A(n_6563),
.Y(n_6990)
);

AOI21x1_ASAP7_75t_L g6991 ( 
.A1(n_6295),
.A2(n_5299),
.B(n_5345),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6696),
.Y(n_6992)
);

INVx2_ASAP7_75t_L g6993 ( 
.A(n_6723),
.Y(n_6993)
);

BUFx3_ASAP7_75t_L g6994 ( 
.A(n_6804),
.Y(n_6994)
);

AND2x2_ASAP7_75t_L g6995 ( 
.A(n_6093),
.B(n_5256),
.Y(n_6995)
);

AOI21xp5_ASAP7_75t_L g6996 ( 
.A1(n_5907),
.A2(n_5653),
.B(n_4741),
.Y(n_6996)
);

BUFx2_ASAP7_75t_L g6997 ( 
.A(n_6638),
.Y(n_6997)
);

AOI22xp33_ASAP7_75t_L g6998 ( 
.A1(n_5951),
.A2(n_4814),
.B1(n_5349),
.B2(n_5725),
.Y(n_6998)
);

CKINVDCx5p33_ASAP7_75t_R g6999 ( 
.A(n_5926),
.Y(n_6999)
);

AOI22xp33_ASAP7_75t_L g7000 ( 
.A1(n_5999),
.A2(n_4814),
.B1(n_5725),
.B2(n_5134),
.Y(n_7000)
);

CKINVDCx20_ASAP7_75t_R g7001 ( 
.A(n_5928),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6093),
.B(n_4711),
.Y(n_7002)
);

INVx2_ASAP7_75t_L g7003 ( 
.A(n_6723),
.Y(n_7003)
);

INVx3_ASAP7_75t_SL g7004 ( 
.A(n_6571),
.Y(n_7004)
);

BUFx2_ASAP7_75t_SL g7005 ( 
.A(n_6097),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_L g7006 ( 
.A(n_6077),
.B(n_4854),
.Y(n_7006)
);

NAND2xp5_ASAP7_75t_L g7007 ( 
.A(n_6294),
.B(n_4854),
.Y(n_7007)
);

CKINVDCx6p67_ASAP7_75t_R g7008 ( 
.A(n_6571),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_6294),
.B(n_4857),
.Y(n_7009)
);

AOI22xp33_ASAP7_75t_L g7010 ( 
.A1(n_5999),
.A2(n_4814),
.B1(n_5687),
.B2(n_5177),
.Y(n_7010)
);

NAND2xp33_ASAP7_75t_L g7011 ( 
.A(n_5797),
.B(n_5431),
.Y(n_7011)
);

NAND2xp5_ASAP7_75t_SL g7012 ( 
.A(n_5959),
.B(n_4790),
.Y(n_7012)
);

INVx3_ASAP7_75t_L g7013 ( 
.A(n_5766),
.Y(n_7013)
);

AND2x2_ASAP7_75t_L g7014 ( 
.A(n_6102),
.B(n_4739),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6730),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_6696),
.Y(n_7016)
);

HB1xp67_ASAP7_75t_L g7017 ( 
.A(n_5817),
.Y(n_7017)
);

INVx4_ASAP7_75t_L g7018 ( 
.A(n_6571),
.Y(n_7018)
);

CKINVDCx16_ASAP7_75t_R g7019 ( 
.A(n_6289),
.Y(n_7019)
);

AOI21xp5_ASAP7_75t_L g7020 ( 
.A1(n_5907),
.A2(n_4741),
.B(n_4727),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6715),
.Y(n_7021)
);

BUFx12f_ASAP7_75t_L g7022 ( 
.A(n_6622),
.Y(n_7022)
);

CKINVDCx20_ASAP7_75t_R g7023 ( 
.A(n_5928),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6715),
.Y(n_7024)
);

INVx4_ASAP7_75t_L g7025 ( 
.A(n_6571),
.Y(n_7025)
);

NAND2xp5_ASAP7_75t_L g7026 ( 
.A(n_6330),
.B(n_4857),
.Y(n_7026)
);

NAND2x1p5_ASAP7_75t_L g7027 ( 
.A(n_6224),
.B(n_5676),
.Y(n_7027)
);

O2A1O1Ixp5_ASAP7_75t_SL g7028 ( 
.A1(n_6437),
.A2(n_5192),
.B(n_5202),
.C(n_5195),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_5740),
.Y(n_7029)
);

NAND2xp5_ASAP7_75t_L g7030 ( 
.A(n_6330),
.B(n_4857),
.Y(n_7030)
);

NAND2xp5_ASAP7_75t_L g7031 ( 
.A(n_6161),
.B(n_6279),
.Y(n_7031)
);

INVx2_ASAP7_75t_SL g7032 ( 
.A(n_6855),
.Y(n_7032)
);

AOI21xp5_ASAP7_75t_L g7033 ( 
.A1(n_5953),
.A2(n_4741),
.B(n_4727),
.Y(n_7033)
);

HB1xp67_ASAP7_75t_L g7034 ( 
.A(n_5852),
.Y(n_7034)
);

AOI21xp5_ASAP7_75t_L g7035 ( 
.A1(n_5953),
.A2(n_4741),
.B(n_4727),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_5740),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_6161),
.B(n_4869),
.Y(n_7037)
);

BUFx2_ASAP7_75t_L g7038 ( 
.A(n_6638),
.Y(n_7038)
);

AND2x4_ASAP7_75t_L g7039 ( 
.A(n_6280),
.B(n_6303),
.Y(n_7039)
);

BUFx6f_ASAP7_75t_L g7040 ( 
.A(n_6283),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_L g7041 ( 
.A1(n_5950),
.A2(n_5177),
.B1(n_5244),
.B2(n_5167),
.Y(n_7041)
);

AOI22xp5_ASAP7_75t_L g7042 ( 
.A1(n_5997),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7042)
);

AOI22x1_ASAP7_75t_L g7043 ( 
.A1(n_5973),
.A2(n_5486),
.B1(n_5539),
.B2(n_5496),
.Y(n_7043)
);

NAND2x1_ASAP7_75t_SL g7044 ( 
.A(n_6426),
.B(n_4486),
.Y(n_7044)
);

CKINVDCx5p33_ASAP7_75t_R g7045 ( 
.A(n_5947),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_5742),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6279),
.B(n_4869),
.Y(n_7047)
);

AND2x2_ASAP7_75t_L g7048 ( 
.A(n_6102),
.B(n_4739),
.Y(n_7048)
);

INVx3_ASAP7_75t_SL g7049 ( 
.A(n_6262),
.Y(n_7049)
);

NAND2xp5_ASAP7_75t_L g7050 ( 
.A(n_6159),
.B(n_6278),
.Y(n_7050)
);

AOI21xp5_ASAP7_75t_L g7051 ( 
.A1(n_5964),
.A2(n_5965),
.B(n_5969),
.Y(n_7051)
);

OR2x6_ASAP7_75t_L g7052 ( 
.A(n_6368),
.B(n_5689),
.Y(n_7052)
);

BUFx3_ASAP7_75t_L g7053 ( 
.A(n_6807),
.Y(n_7053)
);

CKINVDCx20_ASAP7_75t_R g7054 ( 
.A(n_5994),
.Y(n_7054)
);

NAND2x1p5_ASAP7_75t_L g7055 ( 
.A(n_6459),
.B(n_5676),
.Y(n_7055)
);

AOI22xp5_ASAP7_75t_L g7056 ( 
.A1(n_5997),
.A2(n_5950),
.B1(n_6069),
.B2(n_5812),
.Y(n_7056)
);

AOI21xp5_ASAP7_75t_L g7057 ( 
.A1(n_5964),
.A2(n_4741),
.B(n_4727),
.Y(n_7057)
);

AND2x2_ASAP7_75t_L g7058 ( 
.A(n_6102),
.B(n_4739),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_5742),
.Y(n_7059)
);

INVx1_ASAP7_75t_SL g7060 ( 
.A(n_6539),
.Y(n_7060)
);

BUFx3_ASAP7_75t_L g7061 ( 
.A(n_6807),
.Y(n_7061)
);

INVx3_ASAP7_75t_L g7062 ( 
.A(n_5766),
.Y(n_7062)
);

OAI22xp5_ASAP7_75t_L g7063 ( 
.A1(n_5779),
.A2(n_5390),
.B1(n_4840),
.B2(n_4818),
.Y(n_7063)
);

AOI22xp33_ASAP7_75t_L g7064 ( 
.A1(n_6000),
.A2(n_5177),
.B1(n_5178),
.B2(n_5167),
.Y(n_7064)
);

INVx2_ASAP7_75t_SL g7065 ( 
.A(n_6855),
.Y(n_7065)
);

INVx4_ASAP7_75t_L g7066 ( 
.A(n_6066),
.Y(n_7066)
);

AOI22xp33_ASAP7_75t_L g7067 ( 
.A1(n_6000),
.A2(n_5177),
.B1(n_5178),
.B2(n_5167),
.Y(n_7067)
);

INVx3_ASAP7_75t_L g7068 ( 
.A(n_5766),
.Y(n_7068)
);

NAND2xp5_ASAP7_75t_L g7069 ( 
.A(n_6159),
.B(n_4869),
.Y(n_7069)
);

AOI221xp5_ASAP7_75t_L g7070 ( 
.A1(n_5858),
.A2(n_4878),
.B1(n_4881),
.B2(n_4877),
.C(n_4871),
.Y(n_7070)
);

BUFx6f_ASAP7_75t_L g7071 ( 
.A(n_6283),
.Y(n_7071)
);

NAND2xp5_ASAP7_75t_L g7072 ( 
.A(n_6278),
.B(n_6286),
.Y(n_7072)
);

OA21x2_ASAP7_75t_L g7073 ( 
.A1(n_5965),
.A2(n_5195),
.B(n_5192),
.Y(n_7073)
);

BUFx3_ASAP7_75t_L g7074 ( 
.A(n_6807),
.Y(n_7074)
);

HB1xp67_ASAP7_75t_L g7075 ( 
.A(n_5852),
.Y(n_7075)
);

CKINVDCx6p67_ASAP7_75t_R g7076 ( 
.A(n_6262),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_5777),
.Y(n_7077)
);

HB1xp67_ASAP7_75t_L g7078 ( 
.A(n_5931),
.Y(n_7078)
);

BUFx2_ASAP7_75t_L g7079 ( 
.A(n_6921),
.Y(n_7079)
);

INVx2_ASAP7_75t_SL g7080 ( 
.A(n_6855),
.Y(n_7080)
);

AND2x4_ASAP7_75t_L g7081 ( 
.A(n_6303),
.B(n_6313),
.Y(n_7081)
);

AOI22xp5_ASAP7_75t_L g7082 ( 
.A1(n_6069),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7082)
);

NAND2xp5_ASAP7_75t_L g7083 ( 
.A(n_6286),
.B(n_6355),
.Y(n_7083)
);

INVx1_ASAP7_75t_SL g7084 ( 
.A(n_6539),
.Y(n_7084)
);

BUFx3_ASAP7_75t_L g7085 ( 
.A(n_6807),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_5777),
.Y(n_7086)
);

NOR2x1_ASAP7_75t_SL g7087 ( 
.A(n_6623),
.B(n_4583),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_5782),
.Y(n_7088)
);

A2O1A1Ixp33_ASAP7_75t_L g7089 ( 
.A1(n_5946),
.A2(n_4583),
.B(n_5375),
.C(n_5334),
.Y(n_7089)
);

AOI22xp33_ASAP7_75t_L g7090 ( 
.A1(n_5797),
.A2(n_5177),
.B1(n_5178),
.B2(n_5167),
.Y(n_7090)
);

INVx3_ASAP7_75t_L g7091 ( 
.A(n_5766),
.Y(n_7091)
);

INVx3_ASAP7_75t_L g7092 ( 
.A(n_5766),
.Y(n_7092)
);

BUFx12f_ASAP7_75t_L g7093 ( 
.A(n_6622),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_L g7094 ( 
.A(n_6355),
.B(n_4871),
.Y(n_7094)
);

AO21x1_ASAP7_75t_L g7095 ( 
.A1(n_6158),
.A2(n_4992),
.B(n_4985),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_5782),
.Y(n_7096)
);

HB1xp67_ASAP7_75t_L g7097 ( 
.A(n_5931),
.Y(n_7097)
);

BUFx6f_ASAP7_75t_L g7098 ( 
.A(n_6283),
.Y(n_7098)
);

OAI22xp5_ASAP7_75t_L g7099 ( 
.A1(n_5779),
.A2(n_5390),
.B1(n_4818),
.B2(n_4840),
.Y(n_7099)
);

NOR2xp33_ASAP7_75t_L g7100 ( 
.A(n_5881),
.B(n_5476),
.Y(n_7100)
);

INVx2_ASAP7_75t_L g7101 ( 
.A(n_6746),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6746),
.Y(n_7102)
);

CKINVDCx5p33_ASAP7_75t_R g7103 ( 
.A(n_5947),
.Y(n_7103)
);

OR2x2_ASAP7_75t_L g7104 ( 
.A(n_6407),
.B(n_4985),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_5786),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_6354),
.B(n_4871),
.Y(n_7106)
);

AOI21xp5_ASAP7_75t_L g7107 ( 
.A1(n_5969),
.A2(n_4741),
.B(n_4727),
.Y(n_7107)
);

AOI22xp33_ASAP7_75t_L g7108 ( 
.A1(n_6023),
.A2(n_5178),
.B1(n_5244),
.B2(n_5167),
.Y(n_7108)
);

NOR2x1_ASAP7_75t_SL g7109 ( 
.A(n_6623),
.B(n_4485),
.Y(n_7109)
);

AOI21xp5_ASAP7_75t_L g7110 ( 
.A1(n_5973),
.A2(n_4741),
.B(n_4727),
.Y(n_7110)
);

INVx1_ASAP7_75t_SL g7111 ( 
.A(n_6539),
.Y(n_7111)
);

INVx2_ASAP7_75t_L g7112 ( 
.A(n_6746),
.Y(n_7112)
);

AOI22xp33_ASAP7_75t_L g7113 ( 
.A1(n_6023),
.A2(n_5178),
.B1(n_5244),
.B2(n_5167),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_5786),
.Y(n_7114)
);

BUFx2_ASAP7_75t_L g7115 ( 
.A(n_6921),
.Y(n_7115)
);

NAND2xp5_ASAP7_75t_L g7116 ( 
.A(n_6354),
.B(n_4877),
.Y(n_7116)
);

INVx1_ASAP7_75t_SL g7117 ( 
.A(n_6546),
.Y(n_7117)
);

BUFx6f_ASAP7_75t_L g7118 ( 
.A(n_5762),
.Y(n_7118)
);

INVxp67_ASAP7_75t_SL g7119 ( 
.A(n_6546),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_5788),
.Y(n_7120)
);

OAI221xp5_ASAP7_75t_L g7121 ( 
.A1(n_5858),
.A2(n_4561),
.B1(n_4557),
.B2(n_4705),
.C(n_4704),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_L g7122 ( 
.A(n_5984),
.B(n_6016),
.Y(n_7122)
);

BUFx6f_ASAP7_75t_L g7123 ( 
.A(n_5762),
.Y(n_7123)
);

AOI22xp33_ASAP7_75t_L g7124 ( 
.A1(n_6080),
.A2(n_5178),
.B1(n_5244),
.B2(n_5167),
.Y(n_7124)
);

INVx2_ASAP7_75t_L g7125 ( 
.A(n_6746),
.Y(n_7125)
);

INVx5_ASAP7_75t_L g7126 ( 
.A(n_6468),
.Y(n_7126)
);

INVx1_ASAP7_75t_SL g7127 ( 
.A(n_6546),
.Y(n_7127)
);

AOI21xp5_ASAP7_75t_L g7128 ( 
.A1(n_6073),
.A2(n_4741),
.B(n_4727),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_5788),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_6750),
.Y(n_7130)
);

INVx2_ASAP7_75t_L g7131 ( 
.A(n_6750),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_5984),
.B(n_4877),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_5802),
.Y(n_7133)
);

INVx2_ASAP7_75t_SL g7134 ( 
.A(n_6721),
.Y(n_7134)
);

AOI22xp5_ASAP7_75t_L g7135 ( 
.A1(n_5812),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_5802),
.Y(n_7136)
);

NAND2x1_ASAP7_75t_SL g7137 ( 
.A(n_6426),
.B(n_4486),
.Y(n_7137)
);

BUFx12f_ASAP7_75t_L g7138 ( 
.A(n_5851),
.Y(n_7138)
);

CKINVDCx20_ASAP7_75t_R g7139 ( 
.A(n_5994),
.Y(n_7139)
);

NAND2xp5_ASAP7_75t_L g7140 ( 
.A(n_6016),
.B(n_6024),
.Y(n_7140)
);

INVx3_ASAP7_75t_L g7141 ( 
.A(n_5806),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6750),
.Y(n_7142)
);

A2O1A1Ixp33_ASAP7_75t_L g7143 ( 
.A1(n_6175),
.A2(n_5375),
.B(n_5393),
.C(n_5334),
.Y(n_7143)
);

INVx4_ASAP7_75t_L g7144 ( 
.A(n_6066),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_L g7145 ( 
.A(n_6024),
.B(n_4878),
.Y(n_7145)
);

AO21x2_ASAP7_75t_L g7146 ( 
.A1(n_6437),
.A2(n_5595),
.B(n_5593),
.Y(n_7146)
);

AOI22xp33_ASAP7_75t_L g7147 ( 
.A1(n_6080),
.A2(n_5178),
.B1(n_5252),
.B2(n_5177),
.Y(n_7147)
);

BUFx6f_ASAP7_75t_L g7148 ( 
.A(n_5762),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_L g7149 ( 
.A(n_6276),
.B(n_4878),
.Y(n_7149)
);

INVx3_ASAP7_75t_L g7150 ( 
.A(n_5806),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_5803),
.Y(n_7151)
);

INVx2_ASAP7_75t_L g7152 ( 
.A(n_6750),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_5803),
.Y(n_7153)
);

INVx2_ASAP7_75t_SL g7154 ( 
.A(n_6721),
.Y(n_7154)
);

INVx2_ASAP7_75t_L g7155 ( 
.A(n_6766),
.Y(n_7155)
);

INVx3_ASAP7_75t_L g7156 ( 
.A(n_5806),
.Y(n_7156)
);

NOR2xp67_ASAP7_75t_L g7157 ( 
.A(n_5761),
.B(n_5051),
.Y(n_7157)
);

HB1xp67_ASAP7_75t_L g7158 ( 
.A(n_6005),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6766),
.Y(n_7159)
);

BUFx2_ASAP7_75t_L g7160 ( 
.A(n_5741),
.Y(n_7160)
);

BUFx8_ASAP7_75t_L g7161 ( 
.A(n_6767),
.Y(n_7161)
);

BUFx2_ASAP7_75t_L g7162 ( 
.A(n_5741),
.Y(n_7162)
);

AOI21xp5_ASAP7_75t_L g7163 ( 
.A1(n_6073),
.A2(n_4727),
.B(n_5710),
.Y(n_7163)
);

CKINVDCx8_ASAP7_75t_R g7164 ( 
.A(n_6068),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_5808),
.Y(n_7165)
);

BUFx12f_ASAP7_75t_L g7166 ( 
.A(n_5851),
.Y(n_7166)
);

OAI22xp33_ASAP7_75t_L g7167 ( 
.A1(n_6099),
.A2(n_5281),
.B1(n_5375),
.B2(n_5334),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_5808),
.Y(n_7168)
);

NOR3xp33_ASAP7_75t_L g7169 ( 
.A(n_6042),
.B(n_5291),
.C(n_5285),
.Y(n_7169)
);

AOI22xp33_ASAP7_75t_L g7170 ( 
.A1(n_6086),
.A2(n_5178),
.B1(n_5244),
.B2(n_5177),
.Y(n_7170)
);

AND2x2_ASAP7_75t_SL g7171 ( 
.A(n_5938),
.B(n_4705),
.Y(n_7171)
);

INVx5_ASAP7_75t_L g7172 ( 
.A(n_6468),
.Y(n_7172)
);

INVx3_ASAP7_75t_L g7173 ( 
.A(n_5806),
.Y(n_7173)
);

BUFx2_ASAP7_75t_L g7174 ( 
.A(n_5741),
.Y(n_7174)
);

AOI22xp33_ASAP7_75t_L g7175 ( 
.A1(n_6086),
.A2(n_5252),
.B1(n_5255),
.B2(n_5244),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_6012),
.B(n_4769),
.Y(n_7176)
);

OR2x2_ASAP7_75t_SL g7177 ( 
.A(n_6127),
.B(n_4485),
.Y(n_7177)
);

INVx2_ASAP7_75t_L g7178 ( 
.A(n_6766),
.Y(n_7178)
);

XNOR2xp5_ASAP7_75t_L g7179 ( 
.A(n_5995),
.B(n_5510),
.Y(n_7179)
);

OR2x2_ASAP7_75t_L g7180 ( 
.A(n_6407),
.B(n_4992),
.Y(n_7180)
);

INVx4_ASAP7_75t_L g7181 ( 
.A(n_6066),
.Y(n_7181)
);

INVx2_ASAP7_75t_SL g7182 ( 
.A(n_6721),
.Y(n_7182)
);

INVx1_ASAP7_75t_SL g7183 ( 
.A(n_6554),
.Y(n_7183)
);

NAND2xp5_ASAP7_75t_L g7184 ( 
.A(n_6276),
.B(n_4881),
.Y(n_7184)
);

OAI22xp5_ASAP7_75t_L g7185 ( 
.A1(n_5901),
.A2(n_5281),
.B1(n_4918),
.B2(n_4793),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6766),
.Y(n_7186)
);

INVx1_ASAP7_75t_SL g7187 ( 
.A(n_6554),
.Y(n_7187)
);

AND2x2_ASAP7_75t_L g7188 ( 
.A(n_6012),
.B(n_4769),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_6012),
.B(n_4769),
.Y(n_7189)
);

INVx2_ASAP7_75t_L g7190 ( 
.A(n_6769),
.Y(n_7190)
);

AOI21xp5_ASAP7_75t_L g7191 ( 
.A1(n_6089),
.A2(n_5710),
.B(n_5714),
.Y(n_7191)
);

BUFx2_ASAP7_75t_L g7192 ( 
.A(n_5768),
.Y(n_7192)
);

AOI21xp5_ASAP7_75t_L g7193 ( 
.A1(n_6089),
.A2(n_5719),
.B(n_5714),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_6407),
.B(n_4881),
.Y(n_7194)
);

AOI22xp33_ASAP7_75t_L g7195 ( 
.A1(n_6241),
.A2(n_5252),
.B1(n_5258),
.B2(n_5255),
.Y(n_7195)
);

BUFx6f_ASAP7_75t_L g7196 ( 
.A(n_5762),
.Y(n_7196)
);

INVx2_ASAP7_75t_SL g7197 ( 
.A(n_6721),
.Y(n_7197)
);

INVx2_ASAP7_75t_L g7198 ( 
.A(n_6769),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_5809),
.Y(n_7199)
);

AOI22xp33_ASAP7_75t_L g7200 ( 
.A1(n_6241),
.A2(n_5252),
.B1(n_5258),
.B2(n_5255),
.Y(n_7200)
);

INVx2_ASAP7_75t_L g7201 ( 
.A(n_6769),
.Y(n_7201)
);

NOR2xp33_ASAP7_75t_SL g7202 ( 
.A(n_6212),
.B(n_6175),
.Y(n_7202)
);

AOI22xp5_ASAP7_75t_L g7203 ( 
.A1(n_6099),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7203)
);

AOI22xp33_ASAP7_75t_SL g7204 ( 
.A1(n_6342),
.A2(n_5252),
.B1(n_5255),
.B2(n_5244),
.Y(n_7204)
);

OR2x2_ASAP7_75t_L g7205 ( 
.A(n_6413),
.B(n_4997),
.Y(n_7205)
);

INVxp67_ASAP7_75t_L g7206 ( 
.A(n_6563),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_5809),
.Y(n_7207)
);

NAND2xp5_ASAP7_75t_L g7208 ( 
.A(n_6413),
.B(n_4890),
.Y(n_7208)
);

NAND2xp5_ASAP7_75t_L g7209 ( 
.A(n_6413),
.B(n_4890),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6598),
.B(n_4890),
.Y(n_7210)
);

BUFx6f_ASAP7_75t_L g7211 ( 
.A(n_5762),
.Y(n_7211)
);

AND2x4_ASAP7_75t_L g7212 ( 
.A(n_6256),
.B(n_6273),
.Y(n_7212)
);

AOI21xp5_ASAP7_75t_L g7213 ( 
.A1(n_6107),
.A2(n_5719),
.B(n_5709),
.Y(n_7213)
);

BUFx12f_ASAP7_75t_L g7214 ( 
.A(n_5851),
.Y(n_7214)
);

OR2x2_ASAP7_75t_L g7215 ( 
.A(n_6037),
.B(n_4997),
.Y(n_7215)
);

BUFx10_ASAP7_75t_L g7216 ( 
.A(n_6767),
.Y(n_7216)
);

INVx4_ASAP7_75t_L g7217 ( 
.A(n_6066),
.Y(n_7217)
);

AOI22xp33_ASAP7_75t_L g7218 ( 
.A1(n_6042),
.A2(n_5255),
.B1(n_5258),
.B2(n_5244),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_6598),
.B(n_4894),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6769),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_5954),
.B(n_4894),
.Y(n_7221)
);

OR2x2_ASAP7_75t_L g7222 ( 
.A(n_6037),
.B(n_5014),
.Y(n_7222)
);

AOI21xp5_ASAP7_75t_L g7223 ( 
.A1(n_6107),
.A2(n_5709),
.B(n_4791),
.Y(n_7223)
);

INVx2_ASAP7_75t_SL g7224 ( 
.A(n_6256),
.Y(n_7224)
);

BUFx6f_ASAP7_75t_L g7225 ( 
.A(n_5762),
.Y(n_7225)
);

NAND2xp5_ASAP7_75t_L g7226 ( 
.A(n_5954),
.B(n_4894),
.Y(n_7226)
);

O2A1O1Ixp5_ASAP7_75t_L g7227 ( 
.A1(n_5960),
.A2(n_4900),
.B(n_4904),
.C(n_4898),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_L g7228 ( 
.A(n_5981),
.B(n_4898),
.Y(n_7228)
);

AOI21xp5_ASAP7_75t_L g7229 ( 
.A1(n_6174),
.A2(n_4791),
.B(n_4774),
.Y(n_7229)
);

BUFx6f_ASAP7_75t_L g7230 ( 
.A(n_5762),
.Y(n_7230)
);

INVx5_ASAP7_75t_L g7231 ( 
.A(n_6468),
.Y(n_7231)
);

INVx3_ASAP7_75t_SL g7232 ( 
.A(n_6262),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_5821),
.Y(n_7233)
);

BUFx2_ASAP7_75t_L g7234 ( 
.A(n_5768),
.Y(n_7234)
);

CKINVDCx20_ASAP7_75t_R g7235 ( 
.A(n_6059),
.Y(n_7235)
);

AOI21xp5_ASAP7_75t_L g7236 ( 
.A1(n_6174),
.A2(n_4791),
.B(n_4774),
.Y(n_7236)
);

AOI21xp5_ASAP7_75t_L g7237 ( 
.A1(n_6176),
.A2(n_4805),
.B(n_4774),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_5821),
.Y(n_7238)
);

BUFx2_ASAP7_75t_L g7239 ( 
.A(n_5768),
.Y(n_7239)
);

BUFx3_ASAP7_75t_L g7240 ( 
.A(n_6824),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_5822),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_5822),
.Y(n_7242)
);

INVx1_ASAP7_75t_L g7243 ( 
.A(n_5823),
.Y(n_7243)
);

INVx2_ASAP7_75t_SL g7244 ( 
.A(n_5784),
.Y(n_7244)
);

BUFx6f_ASAP7_75t_L g7245 ( 
.A(n_5816),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_5823),
.Y(n_7246)
);

OAI22xp5_ASAP7_75t_L g7247 ( 
.A1(n_5901),
.A2(n_4918),
.B1(n_4793),
.B2(n_5003),
.Y(n_7247)
);

AOI21x1_ASAP7_75t_L g7248 ( 
.A1(n_6295),
.A2(n_5202),
.B(n_5195),
.Y(n_7248)
);

OR2x2_ASAP7_75t_L g7249 ( 
.A(n_6037),
.B(n_5001),
.Y(n_7249)
);

AOI22xp33_ASAP7_75t_L g7250 ( 
.A1(n_6204),
.A2(n_5255),
.B1(n_5258),
.B2(n_5252),
.Y(n_7250)
);

OAI22xp5_ASAP7_75t_L g7251 ( 
.A1(n_6141),
.A2(n_6112),
.B1(n_6053),
.B2(n_6149),
.Y(n_7251)
);

OAI22xp33_ASAP7_75t_L g7252 ( 
.A1(n_6087),
.A2(n_5375),
.B1(n_5393),
.B2(n_5334),
.Y(n_7252)
);

NOR2xp33_ASAP7_75t_L g7253 ( 
.A(n_5881),
.B(n_5482),
.Y(n_7253)
);

AND2x2_ASAP7_75t_L g7254 ( 
.A(n_6035),
.B(n_6547),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_5981),
.B(n_4898),
.Y(n_7255)
);

AOI21xp5_ASAP7_75t_L g7256 ( 
.A1(n_6176),
.A2(n_4816),
.B(n_4811),
.Y(n_7256)
);

AO31x2_ASAP7_75t_L g7257 ( 
.A1(n_6260),
.A2(n_5600),
.A3(n_5606),
.B(n_5595),
.Y(n_7257)
);

INVx2_ASAP7_75t_SL g7258 ( 
.A(n_5784),
.Y(n_7258)
);

INVx2_ASAP7_75t_SL g7259 ( 
.A(n_5784),
.Y(n_7259)
);

HAxp5_ASAP7_75t_L g7260 ( 
.A(n_6123),
.B(n_5196),
.CON(n_7260),
.SN(n_7260)
);

AOI22xp33_ASAP7_75t_L g7261 ( 
.A1(n_6204),
.A2(n_5258),
.B1(n_5266),
.B2(n_5252),
.Y(n_7261)
);

BUFx2_ASAP7_75t_L g7262 ( 
.A(n_6573),
.Y(n_7262)
);

AOI22xp33_ASAP7_75t_L g7263 ( 
.A1(n_6162),
.A2(n_5258),
.B1(n_5266),
.B2(n_5252),
.Y(n_7263)
);

BUFx3_ASAP7_75t_L g7264 ( 
.A(n_6824),
.Y(n_7264)
);

HB1xp67_ASAP7_75t_L g7265 ( 
.A(n_6005),
.Y(n_7265)
);

BUFx2_ASAP7_75t_L g7266 ( 
.A(n_6573),
.Y(n_7266)
);

INVx3_ASAP7_75t_L g7267 ( 
.A(n_5806),
.Y(n_7267)
);

AOI21xp5_ASAP7_75t_L g7268 ( 
.A1(n_6186),
.A2(n_4824),
.B(n_4822),
.Y(n_7268)
);

AOI21xp5_ASAP7_75t_L g7269 ( 
.A1(n_6186),
.A2(n_4824),
.B(n_4822),
.Y(n_7269)
);

AOI22xp5_ASAP7_75t_L g7270 ( 
.A1(n_6087),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7270)
);

NAND2xp5_ASAP7_75t_L g7271 ( 
.A(n_6046),
.B(n_4900),
.Y(n_7271)
);

AOI22xp33_ASAP7_75t_L g7272 ( 
.A1(n_6162),
.A2(n_5258),
.B1(n_5326),
.B2(n_5255),
.Y(n_7272)
);

INVx2_ASAP7_75t_SL g7273 ( 
.A(n_5748),
.Y(n_7273)
);

NAND2x1p5_ASAP7_75t_L g7274 ( 
.A(n_6459),
.B(n_5676),
.Y(n_7274)
);

CKINVDCx20_ASAP7_75t_R g7275 ( 
.A(n_6059),
.Y(n_7275)
);

INVx3_ASAP7_75t_L g7276 ( 
.A(n_5840),
.Y(n_7276)
);

AOI22xp33_ASAP7_75t_L g7277 ( 
.A1(n_6217),
.A2(n_5258),
.B1(n_5326),
.B2(n_5255),
.Y(n_7277)
);

INVx2_ASAP7_75t_SL g7278 ( 
.A(n_5748),
.Y(n_7278)
);

OAI22xp5_ASAP7_75t_L g7279 ( 
.A1(n_6141),
.A2(n_4918),
.B1(n_4793),
.B2(n_5067),
.Y(n_7279)
);

CKINVDCx11_ASAP7_75t_R g7280 ( 
.A(n_6801),
.Y(n_7280)
);

NOR2xp33_ASAP7_75t_L g7281 ( 
.A(n_6085),
.B(n_5482),
.Y(n_7281)
);

BUFx12f_ASAP7_75t_L g7282 ( 
.A(n_5859),
.Y(n_7282)
);

BUFx12f_ASAP7_75t_L g7283 ( 
.A(n_5859),
.Y(n_7283)
);

INVx2_ASAP7_75t_SL g7284 ( 
.A(n_5748),
.Y(n_7284)
);

INVx1_ASAP7_75t_SL g7285 ( 
.A(n_6554),
.Y(n_7285)
);

BUFx6f_ASAP7_75t_L g7286 ( 
.A(n_5816),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_6046),
.B(n_4900),
.Y(n_7287)
);

NAND2xp5_ASAP7_75t_L g7288 ( 
.A(n_6062),
.B(n_6071),
.Y(n_7288)
);

CKINVDCx12_ASAP7_75t_R g7289 ( 
.A(n_6764),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_5828),
.Y(n_7290)
);

AND2x2_ASAP7_75t_SL g7291 ( 
.A(n_5938),
.B(n_5108),
.Y(n_7291)
);

NOR2xp33_ASAP7_75t_SL g7292 ( 
.A(n_6212),
.B(n_5028),
.Y(n_7292)
);

O2A1O1Ixp33_ASAP7_75t_L g7293 ( 
.A1(n_5894),
.A2(n_5291),
.B(n_5142),
.C(n_5014),
.Y(n_7293)
);

HB1xp67_ASAP7_75t_L g7294 ( 
.A(n_6039),
.Y(n_7294)
);

INVxp67_ASAP7_75t_L g7295 ( 
.A(n_6675),
.Y(n_7295)
);

BUFx6f_ASAP7_75t_L g7296 ( 
.A(n_5816),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_5828),
.Y(n_7297)
);

OR2x6_ASAP7_75t_L g7298 ( 
.A(n_6388),
.B(n_5689),
.Y(n_7298)
);

OA21x2_ASAP7_75t_L g7299 ( 
.A1(n_6454),
.A2(n_5211),
.B(n_5209),
.Y(n_7299)
);

INVx4_ASAP7_75t_L g7300 ( 
.A(n_6066),
.Y(n_7300)
);

BUFx10_ASAP7_75t_L g7301 ( 
.A(n_6767),
.Y(n_7301)
);

INVx3_ASAP7_75t_L g7302 ( 
.A(n_5840),
.Y(n_7302)
);

INVx3_ASAP7_75t_L g7303 ( 
.A(n_5840),
.Y(n_7303)
);

OAI22xp5_ASAP7_75t_L g7304 ( 
.A1(n_6112),
.A2(n_4918),
.B1(n_4793),
.B2(n_5224),
.Y(n_7304)
);

NAND2x2_ASAP7_75t_L g7305 ( 
.A(n_6708),
.B(n_5665),
.Y(n_7305)
);

NAND2xp5_ASAP7_75t_L g7306 ( 
.A(n_6062),
.B(n_4904),
.Y(n_7306)
);

A2O1A1Ixp33_ASAP7_75t_L g7307 ( 
.A1(n_5960),
.A2(n_5402),
.B(n_5440),
.C(n_5393),
.Y(n_7307)
);

NOR2xp33_ASAP7_75t_L g7308 ( 
.A(n_6085),
.B(n_5482),
.Y(n_7308)
);

BUFx2_ASAP7_75t_L g7309 ( 
.A(n_6573),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_5838),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_L g7311 ( 
.A(n_6071),
.B(n_4904),
.Y(n_7311)
);

BUFx12f_ASAP7_75t_L g7312 ( 
.A(n_5859),
.Y(n_7312)
);

AOI22xp33_ASAP7_75t_L g7313 ( 
.A1(n_6217),
.A2(n_5326),
.B1(n_5374),
.B2(n_5266),
.Y(n_7313)
);

OAI22xp33_ASAP7_75t_L g7314 ( 
.A1(n_6165),
.A2(n_5402),
.B1(n_5440),
.B2(n_5393),
.Y(n_7314)
);

INVx3_ASAP7_75t_L g7315 ( 
.A(n_5840),
.Y(n_7315)
);

INVxp67_ASAP7_75t_SL g7316 ( 
.A(n_6558),
.Y(n_7316)
);

BUFx4f_ASAP7_75t_L g7317 ( 
.A(n_6444),
.Y(n_7317)
);

AOI22xp33_ASAP7_75t_L g7318 ( 
.A1(n_6408),
.A2(n_5326),
.B1(n_5374),
.B2(n_5266),
.Y(n_7318)
);

AOI22xp33_ASAP7_75t_L g7319 ( 
.A1(n_6408),
.A2(n_5326),
.B1(n_5374),
.B2(n_5266),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_6250),
.B(n_4911),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_5838),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_5839),
.Y(n_7322)
);

OR2x6_ASAP7_75t_L g7323 ( 
.A(n_6388),
.B(n_5689),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_6250),
.B(n_4911),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_L g7325 ( 
.A(n_6255),
.B(n_4911),
.Y(n_7325)
);

BUFx12f_ASAP7_75t_L g7326 ( 
.A(n_5865),
.Y(n_7326)
);

INVx2_ASAP7_75t_L g7327 ( 
.A(n_6566),
.Y(n_7327)
);

OAI22xp5_ASAP7_75t_L g7328 ( 
.A1(n_6053),
.A2(n_4918),
.B1(n_4793),
.B2(n_5031),
.Y(n_7328)
);

NAND2xp5_ASAP7_75t_L g7329 ( 
.A(n_6255),
.B(n_4917),
.Y(n_7329)
);

NAND2xp5_ASAP7_75t_L g7330 ( 
.A(n_6265),
.B(n_4917),
.Y(n_7330)
);

AO21x2_ASAP7_75t_L g7331 ( 
.A1(n_6260),
.A2(n_6274),
.B(n_6454),
.Y(n_7331)
);

BUFx6f_ASAP7_75t_L g7332 ( 
.A(n_5816),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_5839),
.Y(n_7333)
);

AOI21xp5_ASAP7_75t_L g7334 ( 
.A1(n_6187),
.A2(n_4831),
.B(n_4829),
.Y(n_7334)
);

BUFx2_ASAP7_75t_L g7335 ( 
.A(n_6619),
.Y(n_7335)
);

NAND2xp5_ASAP7_75t_SL g7336 ( 
.A(n_5959),
.B(n_4485),
.Y(n_7336)
);

NAND2xp5_ASAP7_75t_L g7337 ( 
.A(n_6265),
.B(n_4917),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_5846),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6566),
.Y(n_7339)
);

INVx4_ASAP7_75t_L g7340 ( 
.A(n_6431),
.Y(n_7340)
);

NOR2xp67_ASAP7_75t_L g7341 ( 
.A(n_5761),
.B(n_5051),
.Y(n_7341)
);

INVx1_ASAP7_75t_SL g7342 ( 
.A(n_6558),
.Y(n_7342)
);

NAND2xp5_ASAP7_75t_L g7343 ( 
.A(n_6370),
.B(n_4924),
.Y(n_7343)
);

OR2x6_ASAP7_75t_L g7344 ( 
.A(n_6179),
.B(n_6485),
.Y(n_7344)
);

AOI222xp33_ASAP7_75t_L g7345 ( 
.A1(n_6096),
.A2(n_5079),
.B1(n_5708),
.B2(n_5707),
.C1(n_5505),
.C2(n_5517),
.Y(n_7345)
);

BUFx2_ASAP7_75t_L g7346 ( 
.A(n_6619),
.Y(n_7346)
);

AOI21xp5_ASAP7_75t_L g7347 ( 
.A1(n_6187),
.A2(n_4844),
.B(n_4831),
.Y(n_7347)
);

AND2x2_ASAP7_75t_SL g7348 ( 
.A(n_5938),
.B(n_5108),
.Y(n_7348)
);

NOR2xp33_ASAP7_75t_L g7349 ( 
.A(n_6100),
.B(n_6104),
.Y(n_7349)
);

CKINVDCx5p33_ASAP7_75t_R g7350 ( 
.A(n_6493),
.Y(n_7350)
);

OR2x6_ASAP7_75t_L g7351 ( 
.A(n_6179),
.B(n_5689),
.Y(n_7351)
);

HB1xp67_ASAP7_75t_L g7352 ( 
.A(n_6039),
.Y(n_7352)
);

INVxp67_ASAP7_75t_L g7353 ( 
.A(n_6675),
.Y(n_7353)
);

AOI21xp5_ASAP7_75t_L g7354 ( 
.A1(n_6211),
.A2(n_4848),
.B(n_4844),
.Y(n_7354)
);

INVx3_ASAP7_75t_SL g7355 ( 
.A(n_6794),
.Y(n_7355)
);

OR2x6_ASAP7_75t_L g7356 ( 
.A(n_6179),
.B(n_5689),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_5846),
.Y(n_7357)
);

NOR2xp33_ASAP7_75t_SL g7358 ( 
.A(n_6459),
.B(n_5028),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_5853),
.Y(n_7359)
);

AOI22xp33_ASAP7_75t_L g7360 ( 
.A1(n_5995),
.A2(n_5326),
.B1(n_5374),
.B2(n_5266),
.Y(n_7360)
);

BUFx3_ASAP7_75t_L g7361 ( 
.A(n_6827),
.Y(n_7361)
);

NOR2x1_ASAP7_75t_SL g7362 ( 
.A(n_5841),
.B(n_4485),
.Y(n_7362)
);

NAND2xp5_ASAP7_75t_L g7363 ( 
.A(n_6370),
.B(n_4924),
.Y(n_7363)
);

INVx2_ASAP7_75t_L g7364 ( 
.A(n_6566),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_5853),
.Y(n_7365)
);

OR2x6_ASAP7_75t_L g7366 ( 
.A(n_6179),
.B(n_5689),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_6245),
.B(n_4924),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_L g7368 ( 
.A(n_6245),
.B(n_4925),
.Y(n_7368)
);

INVx1_ASAP7_75t_SL g7369 ( 
.A(n_6558),
.Y(n_7369)
);

BUFx4f_ASAP7_75t_SL g7370 ( 
.A(n_6801),
.Y(n_7370)
);

OAI22xp5_ASAP7_75t_L g7371 ( 
.A1(n_6149),
.A2(n_4918),
.B1(n_4793),
.B2(n_5003),
.Y(n_7371)
);

BUFx6f_ASAP7_75t_L g7372 ( 
.A(n_5816),
.Y(n_7372)
);

A2O1A1Ixp33_ASAP7_75t_SL g7373 ( 
.A1(n_6106),
.A2(n_5695),
.B(n_5675),
.C(n_5583),
.Y(n_7373)
);

INVx5_ASAP7_75t_L g7374 ( 
.A(n_6468),
.Y(n_7374)
);

HB1xp67_ASAP7_75t_L g7375 ( 
.A(n_6040),
.Y(n_7375)
);

CKINVDCx12_ASAP7_75t_R g7376 ( 
.A(n_6764),
.Y(n_7376)
);

INVxp67_ASAP7_75t_L g7377 ( 
.A(n_6770),
.Y(n_7377)
);

INVx2_ASAP7_75t_SL g7378 ( 
.A(n_5748),
.Y(n_7378)
);

BUFx4_ASAP7_75t_SL g7379 ( 
.A(n_6830),
.Y(n_7379)
);

BUFx6f_ASAP7_75t_L g7380 ( 
.A(n_5816),
.Y(n_7380)
);

CKINVDCx5p33_ASAP7_75t_R g7381 ( 
.A(n_6493),
.Y(n_7381)
);

BUFx12f_ASAP7_75t_L g7382 ( 
.A(n_5865),
.Y(n_7382)
);

BUFx3_ASAP7_75t_L g7383 ( 
.A(n_6827),
.Y(n_7383)
);

O2A1O1Ixp5_ASAP7_75t_L g7384 ( 
.A1(n_6169),
.A2(n_4932),
.B(n_4934),
.C(n_4925),
.Y(n_7384)
);

O2A1O1Ixp5_ASAP7_75t_L g7385 ( 
.A1(n_6169),
.A2(n_4932),
.B(n_4934),
.C(n_4925),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_5882),
.Y(n_7386)
);

BUFx6f_ASAP7_75t_L g7387 ( 
.A(n_5816),
.Y(n_7387)
);

BUFx6f_ASAP7_75t_L g7388 ( 
.A(n_5991),
.Y(n_7388)
);

INVx2_ASAP7_75t_SL g7389 ( 
.A(n_6072),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_L g7390 ( 
.A(n_6133),
.B(n_4932),
.Y(n_7390)
);

NAND2xp5_ASAP7_75t_L g7391 ( 
.A(n_6133),
.B(n_6148),
.Y(n_7391)
);

INVx4_ASAP7_75t_L g7392 ( 
.A(n_6431),
.Y(n_7392)
);

AND2x6_ASAP7_75t_L g7393 ( 
.A(n_6215),
.B(n_4486),
.Y(n_7393)
);

INVx1_ASAP7_75t_SL g7394 ( 
.A(n_6619),
.Y(n_7394)
);

NAND2xp5_ASAP7_75t_SL g7395 ( 
.A(n_6154),
.B(n_4485),
.Y(n_7395)
);

BUFx6f_ASAP7_75t_L g7396 ( 
.A(n_5991),
.Y(n_7396)
);

AOI22xp33_ASAP7_75t_L g7397 ( 
.A1(n_6277),
.A2(n_6342),
.B1(n_6154),
.B2(n_6127),
.Y(n_7397)
);

HB1xp67_ASAP7_75t_L g7398 ( 
.A(n_6040),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_5882),
.Y(n_7399)
);

AOI21x1_ASAP7_75t_L g7400 ( 
.A1(n_6295),
.A2(n_5211),
.B(n_5209),
.Y(n_7400)
);

OR2x2_ASAP7_75t_L g7401 ( 
.A(n_6157),
.B(n_5001),
.Y(n_7401)
);

NOR2x1_ASAP7_75t_SL g7402 ( 
.A(n_5841),
.B(n_4485),
.Y(n_7402)
);

BUFx2_ASAP7_75t_L g7403 ( 
.A(n_6635),
.Y(n_7403)
);

INVx5_ASAP7_75t_L g7404 ( 
.A(n_6468),
.Y(n_7404)
);

INVxp67_ASAP7_75t_L g7405 ( 
.A(n_6770),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_5885),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_L g7407 ( 
.A(n_6148),
.B(n_4934),
.Y(n_7407)
);

AOI21xp5_ASAP7_75t_L g7408 ( 
.A1(n_6232),
.A2(n_4861),
.B(n_4848),
.Y(n_7408)
);

AOI22xp5_ASAP7_75t_L g7409 ( 
.A1(n_6234),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7409)
);

NAND2xp5_ASAP7_75t_L g7410 ( 
.A(n_6599),
.B(n_6600),
.Y(n_7410)
);

NOR2xp33_ASAP7_75t_L g7411 ( 
.A(n_6100),
.B(n_5488),
.Y(n_7411)
);

INVx5_ASAP7_75t_L g7412 ( 
.A(n_6468),
.Y(n_7412)
);

BUFx2_ASAP7_75t_R g7413 ( 
.A(n_5866),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_L g7414 ( 
.A(n_6599),
.B(n_4940),
.Y(n_7414)
);

AOI21xp5_ASAP7_75t_L g7415 ( 
.A1(n_6232),
.A2(n_4876),
.B(n_4861),
.Y(n_7415)
);

BUFx2_ASAP7_75t_L g7416 ( 
.A(n_6635),
.Y(n_7416)
);

AOI22xp5_ASAP7_75t_L g7417 ( 
.A1(n_6234),
.A2(n_4666),
.B1(n_4807),
.B2(n_4660),
.Y(n_7417)
);

BUFx2_ASAP7_75t_L g7418 ( 
.A(n_6635),
.Y(n_7418)
);

HB1xp67_ASAP7_75t_L g7419 ( 
.A(n_6220),
.Y(n_7419)
);

O2A1O1Ixp5_ASAP7_75t_L g7420 ( 
.A1(n_6129),
.A2(n_4950),
.B(n_4958),
.C(n_4940),
.Y(n_7420)
);

CKINVDCx20_ASAP7_75t_R g7421 ( 
.A(n_6830),
.Y(n_7421)
);

CKINVDCx20_ASAP7_75t_R g7422 ( 
.A(n_6880),
.Y(n_7422)
);

OAI22xp5_ASAP7_75t_L g7423 ( 
.A1(n_6104),
.A2(n_4918),
.B1(n_4793),
.B2(n_5003),
.Y(n_7423)
);

BUFx10_ASAP7_75t_L g7424 ( 
.A(n_6767),
.Y(n_7424)
);

NAND2xp5_ASAP7_75t_L g7425 ( 
.A(n_6600),
.B(n_4940),
.Y(n_7425)
);

AOI22xp33_ASAP7_75t_SL g7426 ( 
.A1(n_6266),
.A2(n_5300),
.B1(n_5326),
.B2(n_5266),
.Y(n_7426)
);

OAI21xp5_ASAP7_75t_L g7427 ( 
.A1(n_5974),
.A2(n_5400),
.B(n_4561),
.Y(n_7427)
);

NOR2xp33_ASAP7_75t_L g7428 ( 
.A(n_6108),
.B(n_5488),
.Y(n_7428)
);

HB1xp67_ASAP7_75t_L g7429 ( 
.A(n_6220),
.Y(n_7429)
);

INVx1_ASAP7_75t_L g7430 ( 
.A(n_5885),
.Y(n_7430)
);

NAND2xp5_ASAP7_75t_SL g7431 ( 
.A(n_6152),
.B(n_4485),
.Y(n_7431)
);

BUFx2_ASAP7_75t_L g7432 ( 
.A(n_6636),
.Y(n_7432)
);

CKINVDCx11_ASAP7_75t_R g7433 ( 
.A(n_6880),
.Y(n_7433)
);

HB1xp67_ASAP7_75t_L g7434 ( 
.A(n_6269),
.Y(n_7434)
);

INVxp67_ASAP7_75t_SL g7435 ( 
.A(n_6777),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_5891),
.Y(n_7436)
);

HB1xp67_ASAP7_75t_L g7437 ( 
.A(n_6269),
.Y(n_7437)
);

INVxp67_ASAP7_75t_SL g7438 ( 
.A(n_6777),
.Y(n_7438)
);

O2A1O1Ixp33_ASAP7_75t_L g7439 ( 
.A1(n_6029),
.A2(n_5142),
.B(n_5016),
.C(n_5029),
.Y(n_7439)
);

NOR2xp33_ASAP7_75t_L g7440 ( 
.A(n_6108),
.B(n_5488),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_SL g7441 ( 
.A(n_6152),
.B(n_4485),
.Y(n_7441)
);

HB1xp67_ASAP7_75t_L g7442 ( 
.A(n_6290),
.Y(n_7442)
);

CKINVDCx5p33_ASAP7_75t_R g7443 ( 
.A(n_6761),
.Y(n_7443)
);

OAI22xp5_ASAP7_75t_L g7444 ( 
.A1(n_6116),
.A2(n_5031),
.B1(n_5067),
.B2(n_5003),
.Y(n_7444)
);

CKINVDCx5p33_ASAP7_75t_R g7445 ( 
.A(n_6761),
.Y(n_7445)
);

OR2x2_ASAP7_75t_L g7446 ( 
.A(n_6157),
.B(n_5015),
.Y(n_7446)
);

NAND2xp5_ASAP7_75t_L g7447 ( 
.A(n_6409),
.B(n_4950),
.Y(n_7447)
);

OAI21x1_ASAP7_75t_L g7448 ( 
.A1(n_6166),
.A2(n_4561),
.B(n_5600),
.Y(n_7448)
);

INVx2_ASAP7_75t_SL g7449 ( 
.A(n_6072),
.Y(n_7449)
);

OR2x2_ASAP7_75t_L g7450 ( 
.A(n_6157),
.B(n_5015),
.Y(n_7450)
);

INVxp67_ASAP7_75t_L g7451 ( 
.A(n_5873),
.Y(n_7451)
);

AOI22xp5_ASAP7_75t_L g7452 ( 
.A1(n_6165),
.A2(n_4945),
.B1(n_4954),
.B2(n_4807),
.Y(n_7452)
);

INVx1_ASAP7_75t_L g7453 ( 
.A(n_5891),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_5917),
.Y(n_7454)
);

AOI21xp5_ASAP7_75t_L g7455 ( 
.A1(n_6237),
.A2(n_4879),
.B(n_4876),
.Y(n_7455)
);

NAND2xp5_ASAP7_75t_L g7456 ( 
.A(n_6409),
.B(n_4950),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_5917),
.Y(n_7457)
);

OR2x2_ASAP7_75t_SL g7458 ( 
.A(n_6384),
.B(n_4507),
.Y(n_7458)
);

NOR2x1_ASAP7_75t_L g7459 ( 
.A(n_6163),
.B(n_4958),
.Y(n_7459)
);

INVxp67_ASAP7_75t_L g7460 ( 
.A(n_5873),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_5923),
.Y(n_7461)
);

AOI22xp5_ASAP7_75t_L g7462 ( 
.A1(n_6343),
.A2(n_4945),
.B1(n_4954),
.B2(n_4807),
.Y(n_7462)
);

NAND2xp5_ASAP7_75t_L g7463 ( 
.A(n_6312),
.B(n_4958),
.Y(n_7463)
);

INVx2_ASAP7_75t_SL g7464 ( 
.A(n_6072),
.Y(n_7464)
);

AOI21xp5_ASAP7_75t_L g7465 ( 
.A1(n_6240),
.A2(n_6284),
.B(n_6249),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_5923),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_5943),
.Y(n_7467)
);

INVx4_ASAP7_75t_L g7468 ( 
.A(n_6431),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_5943),
.Y(n_7469)
);

OAI22xp5_ASAP7_75t_L g7470 ( 
.A1(n_6116),
.A2(n_5031),
.B1(n_5067),
.B2(n_5003),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_5948),
.Y(n_7471)
);

OAI21x1_ASAP7_75t_L g7472 ( 
.A1(n_6166),
.A2(n_6465),
.B(n_6249),
.Y(n_7472)
);

INVx1_ASAP7_75t_L g7473 ( 
.A(n_5948),
.Y(n_7473)
);

AOI21xp5_ASAP7_75t_L g7474 ( 
.A1(n_6240),
.A2(n_4923),
.B(n_4905),
.Y(n_7474)
);

NAND2xp5_ASAP7_75t_L g7475 ( 
.A(n_6312),
.B(n_6382),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_5958),
.Y(n_7476)
);

BUFx2_ASAP7_75t_L g7477 ( 
.A(n_6636),
.Y(n_7477)
);

INVx4_ASAP7_75t_L g7478 ( 
.A(n_6431),
.Y(n_7478)
);

AOI21xp5_ASAP7_75t_L g7479 ( 
.A1(n_6284),
.A2(n_6306),
.B(n_6304),
.Y(n_7479)
);

NOR2xp33_ASAP7_75t_L g7480 ( 
.A(n_6192),
.B(n_5503),
.Y(n_7480)
);

INVx1_ASAP7_75t_L g7481 ( 
.A(n_5958),
.Y(n_7481)
);

AND2x2_ASAP7_75t_SL g7482 ( 
.A(n_5938),
.B(n_5108),
.Y(n_7482)
);

INVx5_ASAP7_75t_L g7483 ( 
.A(n_6468),
.Y(n_7483)
);

AOI21xp5_ASAP7_75t_L g7484 ( 
.A1(n_6304),
.A2(n_4935),
.B(n_4927),
.Y(n_7484)
);

CKINVDCx5p33_ASAP7_75t_R g7485 ( 
.A(n_5922),
.Y(n_7485)
);

AND2x4_ASAP7_75t_L g7486 ( 
.A(n_6038),
.B(n_6055),
.Y(n_7486)
);

AOI21xp5_ASAP7_75t_L g7487 ( 
.A1(n_6306),
.A2(n_4935),
.B(n_4927),
.Y(n_7487)
);

AOI22xp33_ASAP7_75t_L g7488 ( 
.A1(n_6277),
.A2(n_5300),
.B1(n_5326),
.B2(n_5266),
.Y(n_7488)
);

OAI22xp33_ASAP7_75t_L g7489 ( 
.A1(n_6305),
.A2(n_5402),
.B1(n_5456),
.B2(n_5440),
.Y(n_7489)
);

AOI22xp33_ASAP7_75t_L g7490 ( 
.A1(n_6466),
.A2(n_5374),
.B1(n_5388),
.B2(n_5300),
.Y(n_7490)
);

CKINVDCx14_ASAP7_75t_R g7491 ( 
.A(n_6446),
.Y(n_7491)
);

A2O1A1Ixp33_ASAP7_75t_L g7492 ( 
.A1(n_6092),
.A2(n_5440),
.B(n_5456),
.C(n_5402),
.Y(n_7492)
);

CKINVDCx5p33_ASAP7_75t_R g7493 ( 
.A(n_5922),
.Y(n_7493)
);

NOR2xp67_ASAP7_75t_L g7494 ( 
.A(n_5761),
.B(n_5124),
.Y(n_7494)
);

INVxp67_ASAP7_75t_SL g7495 ( 
.A(n_6380),
.Y(n_7495)
);

AO31x2_ASAP7_75t_L g7496 ( 
.A1(n_6274),
.A2(n_5606),
.A3(n_5211),
.B(n_5220),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_5963),
.Y(n_7497)
);

AOI21xp5_ASAP7_75t_L g7498 ( 
.A1(n_6316),
.A2(n_4935),
.B(n_4927),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_5963),
.Y(n_7499)
);

NAND2xp5_ASAP7_75t_L g7500 ( 
.A(n_6312),
.B(n_4961),
.Y(n_7500)
);

CKINVDCx5p33_ASAP7_75t_R g7501 ( 
.A(n_6402),
.Y(n_7501)
);

BUFx2_ASAP7_75t_L g7502 ( 
.A(n_6636),
.Y(n_7502)
);

AOI21xp5_ASAP7_75t_L g7503 ( 
.A1(n_6316),
.A2(n_4960),
.B(n_4956),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_5967),
.Y(n_7504)
);

AOI221xp5_ASAP7_75t_L g7505 ( 
.A1(n_6096),
.A2(n_4969),
.B1(n_4970),
.B2(n_4962),
.C(n_4961),
.Y(n_7505)
);

HB1xp67_ASAP7_75t_L g7506 ( 
.A(n_6290),
.Y(n_7506)
);

HB1xp67_ASAP7_75t_L g7507 ( 
.A(n_6356),
.Y(n_7507)
);

AOI22xp33_ASAP7_75t_SL g7508 ( 
.A1(n_6266),
.A2(n_5374),
.B1(n_5388),
.B2(n_5300),
.Y(n_7508)
);

AND2x2_ASAP7_75t_SL g7509 ( 
.A(n_5837),
.B(n_5108),
.Y(n_7509)
);

AOI21xp5_ASAP7_75t_L g7510 ( 
.A1(n_6334),
.A2(n_4960),
.B(n_4956),
.Y(n_7510)
);

HB1xp67_ASAP7_75t_L g7511 ( 
.A(n_6356),
.Y(n_7511)
);

BUFx10_ASAP7_75t_L g7512 ( 
.A(n_6767),
.Y(n_7512)
);

OAI22xp5_ASAP7_75t_L g7513 ( 
.A1(n_6192),
.A2(n_5031),
.B1(n_5067),
.B2(n_5003),
.Y(n_7513)
);

BUFx3_ASAP7_75t_L g7514 ( 
.A(n_6851),
.Y(n_7514)
);

AOI22xp33_ASAP7_75t_L g7515 ( 
.A1(n_6466),
.A2(n_5374),
.B1(n_5388),
.B2(n_5300),
.Y(n_7515)
);

INVx2_ASAP7_75t_SL g7516 ( 
.A(n_6072),
.Y(n_7516)
);

AOI22xp5_ASAP7_75t_L g7517 ( 
.A1(n_6343),
.A2(n_4945),
.B1(n_4954),
.B2(n_4807),
.Y(n_7517)
);

NAND2xp5_ASAP7_75t_L g7518 ( 
.A(n_6382),
.B(n_6150),
.Y(n_7518)
);

BUFx2_ASAP7_75t_L g7519 ( 
.A(n_6645),
.Y(n_7519)
);

AOI22xp33_ASAP7_75t_L g7520 ( 
.A1(n_6197),
.A2(n_5374),
.B1(n_5388),
.B2(n_5300),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_5967),
.Y(n_7521)
);

NOR2xp33_ASAP7_75t_L g7522 ( 
.A(n_6197),
.B(n_5503),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_5968),
.Y(n_7523)
);

NAND2xp5_ASAP7_75t_L g7524 ( 
.A(n_6382),
.B(n_4961),
.Y(n_7524)
);

INVx4_ASAP7_75t_L g7525 ( 
.A(n_6431),
.Y(n_7525)
);

INVx2_ASAP7_75t_SL g7526 ( 
.A(n_6072),
.Y(n_7526)
);

CKINVDCx20_ASAP7_75t_R g7527 ( 
.A(n_6601),
.Y(n_7527)
);

NAND3xp33_ASAP7_75t_L g7528 ( 
.A(n_5974),
.B(n_4969),
.C(n_4962),
.Y(n_7528)
);

INVx1_ASAP7_75t_L g7529 ( 
.A(n_5968),
.Y(n_7529)
);

A2O1A1Ixp33_ASAP7_75t_L g7530 ( 
.A1(n_6092),
.A2(n_5472),
.B(n_5487),
.C(n_5456),
.Y(n_7530)
);

CKINVDCx20_ASAP7_75t_R g7531 ( 
.A(n_6601),
.Y(n_7531)
);

NAND2x1_ASAP7_75t_L g7532 ( 
.A(n_6055),
.B(n_5686),
.Y(n_7532)
);

OAI22xp5_ASAP7_75t_L g7533 ( 
.A1(n_6305),
.A2(n_5067),
.B1(n_5109),
.B2(n_5031),
.Y(n_7533)
);

BUFx2_ASAP7_75t_L g7534 ( 
.A(n_6645),
.Y(n_7534)
);

BUFx2_ASAP7_75t_L g7535 ( 
.A(n_6645),
.Y(n_7535)
);

CKINVDCx5p33_ASAP7_75t_R g7536 ( 
.A(n_6803),
.Y(n_7536)
);

OAI22xp5_ASAP7_75t_L g7537 ( 
.A1(n_6289),
.A2(n_6136),
.B1(n_6357),
.B2(n_6065),
.Y(n_7537)
);

NAND2xp5_ASAP7_75t_L g7538 ( 
.A(n_6150),
.B(n_4962),
.Y(n_7538)
);

NAND2xp5_ASAP7_75t_L g7539 ( 
.A(n_6160),
.B(n_4969),
.Y(n_7539)
);

NAND2x1_ASAP7_75t_L g7540 ( 
.A(n_6055),
.B(n_6630),
.Y(n_7540)
);

NAND2x1_ASAP7_75t_L g7541 ( 
.A(n_6055),
.B(n_5686),
.Y(n_7541)
);

INVx4_ASAP7_75t_L g7542 ( 
.A(n_6579),
.Y(n_7542)
);

INVx3_ASAP7_75t_SL g7543 ( 
.A(n_6794),
.Y(n_7543)
);

OR2x2_ASAP7_75t_L g7544 ( 
.A(n_6474),
.B(n_6500),
.Y(n_7544)
);

BUFx4f_ASAP7_75t_SL g7545 ( 
.A(n_5865),
.Y(n_7545)
);

OAI22xp5_ASAP7_75t_L g7546 ( 
.A1(n_6289),
.A2(n_6136),
.B1(n_6357),
.B2(n_6065),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_5970),
.Y(n_7547)
);

NAND2xp5_ASAP7_75t_L g7548 ( 
.A(n_6160),
.B(n_4970),
.Y(n_7548)
);

BUFx12f_ASAP7_75t_L g7549 ( 
.A(n_5876),
.Y(n_7549)
);

A2O1A1Ixp33_ASAP7_75t_SL g7550 ( 
.A1(n_6106),
.A2(n_5962),
.B(n_6281),
.C(n_5952),
.Y(n_7550)
);

AOI222xp33_ASAP7_75t_L g7551 ( 
.A1(n_6111),
.A2(n_5708),
.B1(n_5505),
.B2(n_5517),
.C1(n_5521),
.C2(n_5518),
.Y(n_7551)
);

INVx4_ASAP7_75t_L g7552 ( 
.A(n_6579),
.Y(n_7552)
);

INVx4_ASAP7_75t_SL g7553 ( 
.A(n_5998),
.Y(n_7553)
);

BUFx2_ASAP7_75t_L g7554 ( 
.A(n_6649),
.Y(n_7554)
);

BUFx2_ASAP7_75t_L g7555 ( 
.A(n_6649),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_5970),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_5971),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_5971),
.Y(n_7558)
);

BUFx3_ASAP7_75t_L g7559 ( 
.A(n_6851),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_6504),
.B(n_4970),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_5980),
.Y(n_7561)
);

NOR2xp33_ASAP7_75t_L g7562 ( 
.A(n_6078),
.B(n_5503),
.Y(n_7562)
);

OAI21x1_ASAP7_75t_L g7563 ( 
.A1(n_6166),
.A2(n_5703),
.B(n_5220),
.Y(n_7563)
);

BUFx12f_ASAP7_75t_L g7564 ( 
.A(n_5876),
.Y(n_7564)
);

INVx1_ASAP7_75t_SL g7565 ( 
.A(n_6649),
.Y(n_7565)
);

INVx1_ASAP7_75t_L g7566 ( 
.A(n_5980),
.Y(n_7566)
);

NAND2xp5_ASAP7_75t_L g7567 ( 
.A(n_6504),
.B(n_4971),
.Y(n_7567)
);

BUFx8_ASAP7_75t_L g7568 ( 
.A(n_6057),
.Y(n_7568)
);

INVxp67_ASAP7_75t_SL g7569 ( 
.A(n_6380),
.Y(n_7569)
);

CKINVDCx5p33_ASAP7_75t_R g7570 ( 
.A(n_6803),
.Y(n_7570)
);

AOI22xp33_ASAP7_75t_L g7571 ( 
.A1(n_6301),
.A2(n_5388),
.B1(n_5407),
.B2(n_5300),
.Y(n_7571)
);

AOI21x1_ASAP7_75t_L g7572 ( 
.A1(n_6298),
.A2(n_5220),
.B(n_5209),
.Y(n_7572)
);

NAND2x1_ASAP7_75t_L g7573 ( 
.A(n_6630),
.B(n_5686),
.Y(n_7573)
);

NOR2xp33_ASAP7_75t_L g7574 ( 
.A(n_6078),
.B(n_5505),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_5982),
.Y(n_7575)
);

BUFx3_ASAP7_75t_L g7576 ( 
.A(n_6851),
.Y(n_7576)
);

AND2x4_ASAP7_75t_L g7577 ( 
.A(n_6868),
.B(n_6851),
.Y(n_7577)
);

INVxp67_ASAP7_75t_SL g7578 ( 
.A(n_6564),
.Y(n_7578)
);

INVx2_ASAP7_75t_SL g7579 ( 
.A(n_6081),
.Y(n_7579)
);

AND2x2_ASAP7_75t_SL g7580 ( 
.A(n_5837),
.B(n_5031),
.Y(n_7580)
);

INVx1_ASAP7_75t_SL g7581 ( 
.A(n_6652),
.Y(n_7581)
);

INVx1_ASAP7_75t_L g7582 ( 
.A(n_5982),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_5986),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_5986),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_5987),
.Y(n_7585)
);

HB1xp67_ASAP7_75t_L g7586 ( 
.A(n_6379),
.Y(n_7586)
);

BUFx2_ASAP7_75t_L g7587 ( 
.A(n_6652),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_5987),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_5988),
.Y(n_7589)
);

INVx1_ASAP7_75t_L g7590 ( 
.A(n_5988),
.Y(n_7590)
);

BUFx2_ASAP7_75t_L g7591 ( 
.A(n_6652),
.Y(n_7591)
);

HB1xp67_ASAP7_75t_L g7592 ( 
.A(n_6379),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_6001),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_6001),
.Y(n_7594)
);

NOR2xp33_ASAP7_75t_L g7595 ( 
.A(n_6360),
.B(n_5517),
.Y(n_7595)
);

INVx1_ASAP7_75t_L g7596 ( 
.A(n_6003),
.Y(n_7596)
);

AOI221xp5_ASAP7_75t_L g7597 ( 
.A1(n_6022),
.A2(n_4975),
.B1(n_4982),
.B2(n_4972),
.C(n_4971),
.Y(n_7597)
);

AO22x1_ASAP7_75t_L g7598 ( 
.A1(n_6207),
.A2(n_5890),
.B1(n_5883),
.B2(n_5929),
.Y(n_7598)
);

OR2x2_ASAP7_75t_L g7599 ( 
.A(n_6474),
.B(n_5016),
.Y(n_7599)
);

BUFx3_ASAP7_75t_L g7600 ( 
.A(n_6868),
.Y(n_7600)
);

INVx1_ASAP7_75t_L g7601 ( 
.A(n_6003),
.Y(n_7601)
);

OAI22xp5_ASAP7_75t_L g7602 ( 
.A1(n_6207),
.A2(n_5067),
.B1(n_5224),
.B2(n_5109),
.Y(n_7602)
);

NAND2xp5_ASAP7_75t_SL g7603 ( 
.A(n_6301),
.B(n_4507),
.Y(n_7603)
);

INVx4_ASAP7_75t_L g7604 ( 
.A(n_6579),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_6564),
.B(n_4971),
.Y(n_7605)
);

INVx6_ASAP7_75t_L g7606 ( 
.A(n_5893),
.Y(n_7606)
);

BUFx2_ASAP7_75t_L g7607 ( 
.A(n_6668),
.Y(n_7607)
);

AOI21x1_ASAP7_75t_SL g7608 ( 
.A1(n_5834),
.A2(n_5574),
.B(n_5273),
.Y(n_7608)
);

CKINVDCx20_ASAP7_75t_R g7609 ( 
.A(n_6602),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_6027),
.Y(n_7610)
);

AOI22xp33_ASAP7_75t_L g7611 ( 
.A1(n_6257),
.A2(n_5388),
.B1(n_5407),
.B2(n_5300),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_6027),
.Y(n_7612)
);

O2A1O1Ixp5_ASAP7_75t_L g7613 ( 
.A1(n_6129),
.A2(n_4975),
.B(n_4982),
.C(n_4972),
.Y(n_7613)
);

AOI21xp5_ASAP7_75t_L g7614 ( 
.A1(n_6341),
.A2(n_6394),
.B(n_6363),
.Y(n_7614)
);

NOR2x1_ASAP7_75t_L g7615 ( 
.A(n_6163),
.B(n_6178),
.Y(n_7615)
);

INVx6_ASAP7_75t_L g7616 ( 
.A(n_5893),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6045),
.Y(n_7617)
);

INVx1_ASAP7_75t_L g7618 ( 
.A(n_6045),
.Y(n_7618)
);

OR2x2_ASAP7_75t_L g7619 ( 
.A(n_6474),
.B(n_5029),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_6597),
.B(n_6679),
.Y(n_7620)
);

OAI22xp33_ASAP7_75t_L g7621 ( 
.A1(n_6469),
.A2(n_5472),
.B1(n_5487),
.B2(n_5456),
.Y(n_7621)
);

AOI22xp33_ASAP7_75t_L g7622 ( 
.A1(n_6257),
.A2(n_5407),
.B1(n_5388),
.B2(n_4954),
.Y(n_7622)
);

OR2x2_ASAP7_75t_L g7623 ( 
.A(n_6500),
.B(n_5033),
.Y(n_7623)
);

NAND2xp33_ASAP7_75t_L g7624 ( 
.A(n_6478),
.B(n_5755),
.Y(n_7624)
);

INVxp67_ASAP7_75t_SL g7625 ( 
.A(n_6597),
.Y(n_7625)
);

BUFx2_ASAP7_75t_L g7626 ( 
.A(n_6668),
.Y(n_7626)
);

NAND2xp5_ASAP7_75t_L g7627 ( 
.A(n_6679),
.B(n_4972),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_6047),
.Y(n_7628)
);

O2A1O1Ixp33_ASAP7_75t_L g7629 ( 
.A1(n_6029),
.A2(n_5036),
.B(n_5037),
.C(n_5033),
.Y(n_7629)
);

O2A1O1Ixp33_ASAP7_75t_L g7630 ( 
.A1(n_5962),
.A2(n_5037),
.B(n_5048),
.C(n_5036),
.Y(n_7630)
);

AND2x4_ASAP7_75t_SL g7631 ( 
.A(n_5989),
.B(n_5109),
.Y(n_7631)
);

AND2x4_ASAP7_75t_L g7632 ( 
.A(n_6875),
.B(n_6900),
.Y(n_7632)
);

AOI21xp5_ASAP7_75t_L g7633 ( 
.A1(n_6363),
.A2(n_5088),
.B(n_5082),
.Y(n_7633)
);

INVxp67_ASAP7_75t_L g7634 ( 
.A(n_6070),
.Y(n_7634)
);

AOI21xp5_ASAP7_75t_L g7635 ( 
.A1(n_6394),
.A2(n_5088),
.B(n_5082),
.Y(n_7635)
);

BUFx4f_ASAP7_75t_L g7636 ( 
.A(n_6444),
.Y(n_7636)
);

INVxp67_ASAP7_75t_L g7637 ( 
.A(n_6070),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_6047),
.Y(n_7638)
);

INVx4_ASAP7_75t_L g7639 ( 
.A(n_6579),
.Y(n_7639)
);

HB1xp67_ASAP7_75t_L g7640 ( 
.A(n_6417),
.Y(n_7640)
);

AOI21xp5_ASAP7_75t_L g7641 ( 
.A1(n_6400),
.A2(n_5130),
.B(n_5111),
.Y(n_7641)
);

BUFx2_ASAP7_75t_L g7642 ( 
.A(n_6668),
.Y(n_7642)
);

INVx1_ASAP7_75t_L g7643 ( 
.A(n_6048),
.Y(n_7643)
);

CKINVDCx11_ASAP7_75t_R g7644 ( 
.A(n_6602),
.Y(n_7644)
);

AND2x4_ASAP7_75t_L g7645 ( 
.A(n_6875),
.B(n_6900),
.Y(n_7645)
);

AOI22xp5_ASAP7_75t_L g7646 ( 
.A1(n_5929),
.A2(n_4954),
.B1(n_4945),
.B2(n_5518),
.Y(n_7646)
);

AOI21xp5_ASAP7_75t_L g7647 ( 
.A1(n_6465),
.A2(n_5130),
.B(n_5111),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_6048),
.Y(n_7648)
);

AOI21x1_ASAP7_75t_L g7649 ( 
.A1(n_6298),
.A2(n_6365),
.B(n_6781),
.Y(n_7649)
);

BUFx5_ASAP7_75t_L g7650 ( 
.A(n_6444),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_6064),
.Y(n_7651)
);

BUFx4_ASAP7_75t_SL g7652 ( 
.A(n_6686),
.Y(n_7652)
);

AOI221x1_ASAP7_75t_L g7653 ( 
.A1(n_5985),
.A2(n_5703),
.B1(n_4987),
.B2(n_4988),
.C(n_4982),
.Y(n_7653)
);

AOI21xp5_ASAP7_75t_L g7654 ( 
.A1(n_6011),
.A2(n_5205),
.B(n_5139),
.Y(n_7654)
);

OAI22xp5_ASAP7_75t_L g7655 ( 
.A1(n_5945),
.A2(n_5109),
.B1(n_5225),
.B2(n_5224),
.Y(n_7655)
);

INVx1_ASAP7_75t_L g7656 ( 
.A(n_6064),
.Y(n_7656)
);

AOI21xp5_ASAP7_75t_L g7657 ( 
.A1(n_6011),
.A2(n_6488),
.B(n_6506),
.Y(n_7657)
);

NOR2xp33_ASAP7_75t_L g7658 ( 
.A(n_6360),
.B(n_6111),
.Y(n_7658)
);

AOI21xp5_ASAP7_75t_L g7659 ( 
.A1(n_6488),
.A2(n_6506),
.B(n_6428),
.Y(n_7659)
);

NAND2xp5_ASAP7_75t_L g7660 ( 
.A(n_6271),
.B(n_4975),
.Y(n_7660)
);

BUFx2_ASAP7_75t_L g7661 ( 
.A(n_6670),
.Y(n_7661)
);

A2O1A1Ixp33_ASAP7_75t_L g7662 ( 
.A1(n_6143),
.A2(n_5487),
.B(n_5532),
.C(n_5472),
.Y(n_7662)
);

HB1xp67_ASAP7_75t_L g7663 ( 
.A(n_6417),
.Y(n_7663)
);

AOI22xp33_ASAP7_75t_L g7664 ( 
.A1(n_5942),
.A2(n_5407),
.B1(n_5388),
.B2(n_4954),
.Y(n_7664)
);

BUFx3_ASAP7_75t_L g7665 ( 
.A(n_6914),
.Y(n_7665)
);

CKINVDCx5p33_ASAP7_75t_R g7666 ( 
.A(n_5774),
.Y(n_7666)
);

OAI22xp5_ASAP7_75t_L g7667 ( 
.A1(n_5945),
.A2(n_5109),
.B1(n_5225),
.B2(n_5224),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_6084),
.Y(n_7668)
);

OAI222xp33_ASAP7_75t_SL g7669 ( 
.A1(n_6866),
.A2(n_5357),
.B1(n_5454),
.B2(n_5224),
.C1(n_5109),
.C2(n_5292),
.Y(n_7669)
);

CKINVDCx20_ASAP7_75t_R g7670 ( 
.A(n_6686),
.Y(n_7670)
);

CKINVDCx5p33_ASAP7_75t_R g7671 ( 
.A(n_5961),
.Y(n_7671)
);

AOI21xp5_ASAP7_75t_L g7672 ( 
.A1(n_6403),
.A2(n_5205),
.B(n_5139),
.Y(n_7672)
);

AOI21xp5_ASAP7_75t_L g7673 ( 
.A1(n_6403),
.A2(n_5208),
.B(n_5205),
.Y(n_7673)
);

BUFx2_ASAP7_75t_R g7674 ( 
.A(n_5866),
.Y(n_7674)
);

NAND2xp5_ASAP7_75t_L g7675 ( 
.A(n_6271),
.B(n_4987),
.Y(n_7675)
);

AOI21x1_ASAP7_75t_L g7676 ( 
.A1(n_6298),
.A2(n_5242),
.B(n_5228),
.Y(n_7676)
);

NAND2xp5_ASAP7_75t_L g7677 ( 
.A(n_6054),
.B(n_4987),
.Y(n_7677)
);

CKINVDCx11_ASAP7_75t_R g7678 ( 
.A(n_6695),
.Y(n_7678)
);

HAxp5_ASAP7_75t_L g7679 ( 
.A(n_6123),
.B(n_5196),
.CON(n_7679),
.SN(n_7679)
);

A2O1A1Ixp33_ASAP7_75t_SL g7680 ( 
.A1(n_6281),
.A2(n_5695),
.B(n_5675),
.C(n_5576),
.Y(n_7680)
);

OAI221xp5_ASAP7_75t_L g7681 ( 
.A1(n_6143),
.A2(n_5487),
.B1(n_5532),
.B2(n_5472),
.C(n_5028),
.Y(n_7681)
);

INVx2_ASAP7_75t_SL g7682 ( 
.A(n_6081),
.Y(n_7682)
);

NAND2xp5_ASAP7_75t_L g7683 ( 
.A(n_6054),
.B(n_4988),
.Y(n_7683)
);

OAI22xp5_ASAP7_75t_L g7684 ( 
.A1(n_6491),
.A2(n_6022),
.B1(n_6025),
.B2(n_6348),
.Y(n_7684)
);

NAND2xp5_ASAP7_75t_L g7685 ( 
.A(n_6611),
.B(n_4988),
.Y(n_7685)
);

BUFx2_ASAP7_75t_L g7686 ( 
.A(n_6670),
.Y(n_7686)
);

BUFx3_ASAP7_75t_L g7687 ( 
.A(n_6914),
.Y(n_7687)
);

OAI22xp5_ASAP7_75t_L g7688 ( 
.A1(n_6491),
.A2(n_5225),
.B1(n_5276),
.B2(n_5224),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_6084),
.Y(n_7689)
);

BUFx2_ASAP7_75t_L g7690 ( 
.A(n_6670),
.Y(n_7690)
);

INVx1_ASAP7_75t_L g7691 ( 
.A(n_6747),
.Y(n_7691)
);

OAI22xp5_ASAP7_75t_SL g7692 ( 
.A1(n_6695),
.A2(n_6471),
.B1(n_6446),
.B2(n_5735),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_6747),
.Y(n_7693)
);

BUFx3_ASAP7_75t_L g7694 ( 
.A(n_5799),
.Y(n_7694)
);

INVx1_ASAP7_75t_L g7695 ( 
.A(n_6753),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_6753),
.Y(n_7696)
);

INVx1_ASAP7_75t_SL g7697 ( 
.A(n_6729),
.Y(n_7697)
);

INVx1_ASAP7_75t_SL g7698 ( 
.A(n_6729),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_6754),
.Y(n_7699)
);

BUFx2_ASAP7_75t_L g7700 ( 
.A(n_6729),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_6754),
.Y(n_7701)
);

AOI22xp33_ASAP7_75t_L g7702 ( 
.A1(n_5942),
.A2(n_5407),
.B1(n_4954),
.B2(n_4945),
.Y(n_7702)
);

CKINVDCx6p67_ASAP7_75t_R g7703 ( 
.A(n_6794),
.Y(n_7703)
);

INVx4_ASAP7_75t_L g7704 ( 
.A(n_6579),
.Y(n_7704)
);

OR2x2_ASAP7_75t_L g7705 ( 
.A(n_6500),
.B(n_6525),
.Y(n_7705)
);

INVx2_ASAP7_75t_SL g7706 ( 
.A(n_6081),
.Y(n_7706)
);

AOI22xp33_ASAP7_75t_L g7707 ( 
.A1(n_5934),
.A2(n_5407),
.B1(n_4954),
.B2(n_4945),
.Y(n_7707)
);

NAND2x1_ASAP7_75t_L g7708 ( 
.A(n_6630),
.B(n_5700),
.Y(n_7708)
);

AOI22xp33_ASAP7_75t_L g7709 ( 
.A1(n_5934),
.A2(n_5407),
.B1(n_4954),
.B2(n_4945),
.Y(n_7709)
);

AOI22xp33_ASAP7_75t_L g7710 ( 
.A1(n_6390),
.A2(n_5407),
.B1(n_4954),
.B2(n_4945),
.Y(n_7710)
);

HB1xp67_ASAP7_75t_L g7711 ( 
.A(n_6424),
.Y(n_7711)
);

AOI22xp33_ASAP7_75t_L g7712 ( 
.A1(n_6390),
.A2(n_4954),
.B1(n_4945),
.B2(n_4989),
.Y(n_7712)
);

AOI22xp33_ASAP7_75t_L g7713 ( 
.A1(n_6443),
.A2(n_4945),
.B1(n_4994),
.B2(n_4989),
.Y(n_7713)
);

INVx1_ASAP7_75t_SL g7714 ( 
.A(n_6780),
.Y(n_7714)
);

AOI21xp5_ASAP7_75t_L g7715 ( 
.A1(n_6428),
.A2(n_6569),
.B(n_6478),
.Y(n_7715)
);

O2A1O1Ixp5_ASAP7_75t_SL g7716 ( 
.A1(n_5985),
.A2(n_5242),
.B(n_5228),
.C(n_5395),
.Y(n_7716)
);

NAND2xp5_ASAP7_75t_L g7717 ( 
.A(n_6611),
.B(n_4989),
.Y(n_7717)
);

AOI21xp5_ASAP7_75t_L g7718 ( 
.A1(n_6569),
.A2(n_5234),
.B(n_5230),
.Y(n_7718)
);

AOI22xp5_ASAP7_75t_L g7719 ( 
.A1(n_6422),
.A2(n_4945),
.B1(n_5521),
.B2(n_5518),
.Y(n_7719)
);

NAND2xp5_ASAP7_75t_SL g7720 ( 
.A(n_5735),
.B(n_4508),
.Y(n_7720)
);

AOI21xp5_ASAP7_75t_L g7721 ( 
.A1(n_6067),
.A2(n_5234),
.B(n_5230),
.Y(n_7721)
);

BUFx12f_ASAP7_75t_L g7722 ( 
.A(n_5876),
.Y(n_7722)
);

NAND2x1_ASAP7_75t_L g7723 ( 
.A(n_6630),
.B(n_5700),
.Y(n_7723)
);

INVx1_ASAP7_75t_SL g7724 ( 
.A(n_6780),
.Y(n_7724)
);

BUFx3_ASAP7_75t_L g7725 ( 
.A(n_5799),
.Y(n_7725)
);

NOR2xp33_ASAP7_75t_L g7726 ( 
.A(n_6103),
.B(n_5521),
.Y(n_7726)
);

NAND2xp5_ASAP7_75t_L g7727 ( 
.A(n_6608),
.B(n_4994),
.Y(n_7727)
);

INVx4_ASAP7_75t_L g7728 ( 
.A(n_6588),
.Y(n_7728)
);

NOR2xp33_ASAP7_75t_R g7729 ( 
.A(n_6886),
.B(n_4880),
.Y(n_7729)
);

CKINVDCx8_ASAP7_75t_R g7730 ( 
.A(n_6068),
.Y(n_7730)
);

BUFx2_ASAP7_75t_L g7731 ( 
.A(n_6780),
.Y(n_7731)
);

INVx2_ASAP7_75t_SL g7732 ( 
.A(n_6081),
.Y(n_7732)
);

HB1xp67_ASAP7_75t_L g7733 ( 
.A(n_6424),
.Y(n_7733)
);

NAND2xp5_ASAP7_75t_L g7734 ( 
.A(n_6608),
.B(n_4994),
.Y(n_7734)
);

AOI22xp5_ASAP7_75t_L g7735 ( 
.A1(n_6422),
.A2(n_6443),
.B1(n_6469),
.B2(n_6494),
.Y(n_7735)
);

BUFx6f_ASAP7_75t_L g7736 ( 
.A(n_6444),
.Y(n_7736)
);

BUFx2_ASAP7_75t_L g7737 ( 
.A(n_6782),
.Y(n_7737)
);

AOI21xp5_ASAP7_75t_L g7738 ( 
.A1(n_6067),
.A2(n_5265),
.B(n_5234),
.Y(n_7738)
);

INVx5_ASAP7_75t_L g7739 ( 
.A(n_6221),
.Y(n_7739)
);

BUFx2_ASAP7_75t_L g7740 ( 
.A(n_6782),
.Y(n_7740)
);

OR2x2_ASAP7_75t_L g7741 ( 
.A(n_6525),
.B(n_5048),
.Y(n_7741)
);

A2O1A1Ixp33_ASAP7_75t_L g7742 ( 
.A1(n_6025),
.A2(n_5532),
.B(n_4496),
.C(n_4592),
.Y(n_7742)
);

BUFx6f_ASAP7_75t_L g7743 ( 
.A(n_6545),
.Y(n_7743)
);

AOI21xp5_ASAP7_75t_L g7744 ( 
.A1(n_6498),
.A2(n_6511),
.B(n_6503),
.Y(n_7744)
);

OAI21xp33_ASAP7_75t_L g7745 ( 
.A1(n_5952),
.A2(n_5574),
.B(n_5053),
.Y(n_7745)
);

CKINVDCx5p33_ASAP7_75t_R g7746 ( 
.A(n_5975),
.Y(n_7746)
);

CKINVDCx5p33_ASAP7_75t_R g7747 ( 
.A(n_5916),
.Y(n_7747)
);

AOI21xp5_ASAP7_75t_L g7748 ( 
.A1(n_6498),
.A2(n_5272),
.B(n_5265),
.Y(n_7748)
);

OAI22xp5_ASAP7_75t_L g7749 ( 
.A1(n_6348),
.A2(n_5276),
.B1(n_5292),
.B2(n_5225),
.Y(n_7749)
);

BUFx2_ASAP7_75t_L g7750 ( 
.A(n_6782),
.Y(n_7750)
);

OAI22xp5_ASAP7_75t_L g7751 ( 
.A1(n_6120),
.A2(n_5276),
.B1(n_5292),
.B2(n_5225),
.Y(n_7751)
);

HB1xp67_ASAP7_75t_L g7752 ( 
.A(n_6432),
.Y(n_7752)
);

NOR2xp33_ASAP7_75t_R g7753 ( 
.A(n_6384),
.B(n_5553),
.Y(n_7753)
);

NAND2xp5_ASAP7_75t_L g7754 ( 
.A(n_6609),
.B(n_6628),
.Y(n_7754)
);

NAND2xp5_ASAP7_75t_L g7755 ( 
.A(n_6609),
.B(n_5002),
.Y(n_7755)
);

BUFx6f_ASAP7_75t_L g7756 ( 
.A(n_6545),
.Y(n_7756)
);

BUFx6f_ASAP7_75t_L g7757 ( 
.A(n_6545),
.Y(n_7757)
);

BUFx3_ASAP7_75t_L g7758 ( 
.A(n_5799),
.Y(n_7758)
);

INVx2_ASAP7_75t_SL g7759 ( 
.A(n_6081),
.Y(n_7759)
);

AOI22xp33_ASAP7_75t_L g7760 ( 
.A1(n_6350),
.A2(n_5005),
.B1(n_5007),
.B2(n_5002),
.Y(n_7760)
);

AOI21xp5_ASAP7_75t_L g7761 ( 
.A1(n_6511),
.A2(n_5307),
.B(n_5272),
.Y(n_7761)
);

NAND2xp5_ASAP7_75t_L g7762 ( 
.A(n_6628),
.B(n_5002),
.Y(n_7762)
);

A2O1A1Ixp33_ASAP7_75t_L g7763 ( 
.A1(n_6103),
.A2(n_5532),
.B(n_4496),
.C(n_4592),
.Y(n_7763)
);

INVx4_ASAP7_75t_L g7764 ( 
.A(n_6588),
.Y(n_7764)
);

BUFx2_ASAP7_75t_L g7765 ( 
.A(n_6870),
.Y(n_7765)
);

INVx4_ASAP7_75t_L g7766 ( 
.A(n_6588),
.Y(n_7766)
);

AOI22xp33_ASAP7_75t_SL g7767 ( 
.A1(n_5890),
.A2(n_4518),
.B1(n_4532),
.B2(n_4508),
.Y(n_7767)
);

AOI22xp5_ASAP7_75t_L g7768 ( 
.A1(n_6494),
.A2(n_5534),
.B1(n_5543),
.B2(n_5526),
.Y(n_7768)
);

AOI21xp5_ASAP7_75t_L g7769 ( 
.A1(n_6503),
.A2(n_5315),
.B(n_5307),
.Y(n_7769)
);

AOI22xp5_ASAP7_75t_L g7770 ( 
.A1(n_5927),
.A2(n_5534),
.B1(n_5543),
.B2(n_5526),
.Y(n_7770)
);

BUFx2_ASAP7_75t_L g7771 ( 
.A(n_6870),
.Y(n_7771)
);

NAND2xp5_ASAP7_75t_L g7772 ( 
.A(n_6395),
.B(n_5005),
.Y(n_7772)
);

BUFx3_ASAP7_75t_L g7773 ( 
.A(n_5799),
.Y(n_7773)
);

NOR2xp33_ASAP7_75t_L g7774 ( 
.A(n_6120),
.B(n_5526),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_6395),
.B(n_5005),
.Y(n_7775)
);

CKINVDCx20_ASAP7_75t_R g7776 ( 
.A(n_6346),
.Y(n_7776)
);

BUFx12f_ASAP7_75t_L g7777 ( 
.A(n_5916),
.Y(n_7777)
);

AOI21xp5_ASAP7_75t_L g7778 ( 
.A1(n_6026),
.A2(n_5315),
.B(n_5307),
.Y(n_7778)
);

BUFx6f_ASAP7_75t_L g7779 ( 
.A(n_6545),
.Y(n_7779)
);

A2O1A1Ixp33_ASAP7_75t_L g7780 ( 
.A1(n_6383),
.A2(n_4496),
.B(n_4592),
.C(n_4503),
.Y(n_7780)
);

AOI22xp33_ASAP7_75t_L g7781 ( 
.A1(n_6350),
.A2(n_5731),
.B1(n_6010),
.B2(n_5897),
.Y(n_7781)
);

INVx3_ASAP7_75t_SL g7782 ( 
.A(n_6139),
.Y(n_7782)
);

HB1xp67_ASAP7_75t_L g7783 ( 
.A(n_6432),
.Y(n_7783)
);

AOI22xp33_ASAP7_75t_L g7784 ( 
.A1(n_5731),
.A2(n_5008),
.B1(n_5011),
.B2(n_5007),
.Y(n_7784)
);

INVxp33_ASAP7_75t_L g7785 ( 
.A(n_5883),
.Y(n_7785)
);

AOI22xp5_ASAP7_75t_L g7786 ( 
.A1(n_5927),
.A2(n_5543),
.B1(n_5544),
.B2(n_5534),
.Y(n_7786)
);

BUFx3_ASAP7_75t_L g7787 ( 
.A(n_5826),
.Y(n_7787)
);

BUFx12f_ASAP7_75t_L g7788 ( 
.A(n_5916),
.Y(n_7788)
);

NAND2xp5_ASAP7_75t_L g7789 ( 
.A(n_6410),
.B(n_5007),
.Y(n_7789)
);

AOI22xp5_ASAP7_75t_L g7790 ( 
.A1(n_6383),
.A2(n_5548),
.B1(n_5550),
.B2(n_5544),
.Y(n_7790)
);

AOI21xp5_ASAP7_75t_L g7791 ( 
.A1(n_6060),
.A2(n_5373),
.B(n_5242),
.Y(n_7791)
);

INVxp67_ASAP7_75t_L g7792 ( 
.A(n_6534),
.Y(n_7792)
);

AOI21xp5_ASAP7_75t_L g7793 ( 
.A1(n_6060),
.A2(n_5228),
.B(n_5671),
.Y(n_7793)
);

NAND2xp5_ASAP7_75t_L g7794 ( 
.A(n_6410),
.B(n_5008),
.Y(n_7794)
);

INVx5_ASAP7_75t_SL g7795 ( 
.A(n_5735),
.Y(n_7795)
);

INVx3_ASAP7_75t_SL g7796 ( 
.A(n_6139),
.Y(n_7796)
);

BUFx6f_ASAP7_75t_L g7797 ( 
.A(n_6365),
.Y(n_7797)
);

BUFx2_ASAP7_75t_SL g7798 ( 
.A(n_6097),
.Y(n_7798)
);

INVx1_ASAP7_75t_SL g7799 ( 
.A(n_6870),
.Y(n_7799)
);

INVx2_ASAP7_75t_SL g7800 ( 
.A(n_6083),
.Y(n_7800)
);

INVx4_ASAP7_75t_L g7801 ( 
.A(n_6588),
.Y(n_7801)
);

AOI22xp5_ASAP7_75t_L g7802 ( 
.A1(n_6386),
.A2(n_5548),
.B1(n_5550),
.B2(n_5544),
.Y(n_7802)
);

BUFx3_ASAP7_75t_L g7803 ( 
.A(n_5826),
.Y(n_7803)
);

NAND2x1p5_ASAP7_75t_L g7804 ( 
.A(n_6481),
.B(n_5700),
.Y(n_7804)
);

INVx2_ASAP7_75t_SL g7805 ( 
.A(n_6083),
.Y(n_7805)
);

OAI22xp5_ASAP7_75t_L g7806 ( 
.A1(n_6146),
.A2(n_5276),
.B1(n_5292),
.B2(n_5225),
.Y(n_7806)
);

AOI22xp33_ASAP7_75t_L g7807 ( 
.A1(n_6010),
.A2(n_5011),
.B1(n_5019),
.B2(n_5008),
.Y(n_7807)
);

OAI22xp5_ASAP7_75t_SL g7808 ( 
.A1(n_6471),
.A2(n_5560),
.B1(n_5588),
.B2(n_5553),
.Y(n_7808)
);

BUFx6f_ASAP7_75t_L g7809 ( 
.A(n_6365),
.Y(n_7809)
);

INVx2_ASAP7_75t_SL g7810 ( 
.A(n_6083),
.Y(n_7810)
);

INVx1_ASAP7_75t_SL g7811 ( 
.A(n_6890),
.Y(n_7811)
);

OA21x2_ASAP7_75t_L g7812 ( 
.A1(n_6907),
.A2(n_5679),
.B(n_5053),
.Y(n_7812)
);

NAND2xp5_ASAP7_75t_L g7813 ( 
.A(n_6034),
.B(n_6331),
.Y(n_7813)
);

AOI21xp5_ASAP7_75t_L g7814 ( 
.A1(n_6026),
.A2(n_5692),
.B(n_5671),
.Y(n_7814)
);

NAND2xp5_ASAP7_75t_L g7815 ( 
.A(n_6034),
.B(n_5011),
.Y(n_7815)
);

BUFx8_ASAP7_75t_SL g7816 ( 
.A(n_6082),
.Y(n_7816)
);

BUFx2_ASAP7_75t_L g7817 ( 
.A(n_6890),
.Y(n_7817)
);

OAI22xp5_ASAP7_75t_L g7818 ( 
.A1(n_6146),
.A2(n_5292),
.B1(n_5308),
.B2(n_5276),
.Y(n_7818)
);

BUFx6f_ASAP7_75t_L g7819 ( 
.A(n_6097),
.Y(n_7819)
);

NAND2xp5_ASAP7_75t_L g7820 ( 
.A(n_6034),
.B(n_5019),
.Y(n_7820)
);

BUFx6f_ASAP7_75t_L g7821 ( 
.A(n_6228),
.Y(n_7821)
);

AOI22xp5_ASAP7_75t_L g7822 ( 
.A1(n_6386),
.A2(n_5550),
.B1(n_5551),
.B2(n_5548),
.Y(n_7822)
);

BUFx2_ASAP7_75t_L g7823 ( 
.A(n_6890),
.Y(n_7823)
);

AOI22xp5_ASAP7_75t_L g7824 ( 
.A1(n_6378),
.A2(n_5557),
.B1(n_5551),
.B2(n_5720),
.Y(n_7824)
);

AND2x2_ASAP7_75t_SL g7825 ( 
.A(n_5837),
.B(n_5276),
.Y(n_7825)
);

CKINVDCx5p33_ASAP7_75t_R g7826 ( 
.A(n_6082),
.Y(n_7826)
);

NAND2xp5_ASAP7_75t_L g7827 ( 
.A(n_6331),
.B(n_6392),
.Y(n_7827)
);

OAI22xp5_ASAP7_75t_L g7828 ( 
.A1(n_5796),
.A2(n_5308),
.B1(n_5369),
.B2(n_5292),
.Y(n_7828)
);

BUFx2_ASAP7_75t_L g7829 ( 
.A(n_6906),
.Y(n_7829)
);

AOI21xp5_ASAP7_75t_L g7830 ( 
.A1(n_6036),
.A2(n_5692),
.B(n_5671),
.Y(n_7830)
);

BUFx2_ASAP7_75t_SL g7831 ( 
.A(n_6228),
.Y(n_7831)
);

CKINVDCx5p33_ASAP7_75t_R g7832 ( 
.A(n_6082),
.Y(n_7832)
);

INVx1_ASAP7_75t_SL g7833 ( 
.A(n_6906),
.Y(n_7833)
);

BUFx6f_ASAP7_75t_L g7834 ( 
.A(n_6228),
.Y(n_7834)
);

AOI22xp33_ASAP7_75t_L g7835 ( 
.A1(n_5897),
.A2(n_5021),
.B1(n_5035),
.B2(n_5019),
.Y(n_7835)
);

BUFx2_ASAP7_75t_L g7836 ( 
.A(n_6906),
.Y(n_7836)
);

AOI21xp5_ASAP7_75t_L g7837 ( 
.A1(n_6036),
.A2(n_5692),
.B(n_5632),
.Y(n_7837)
);

INVx2_ASAP7_75t_SL g7838 ( 
.A(n_6083),
.Y(n_7838)
);

BUFx3_ASAP7_75t_L g7839 ( 
.A(n_5826),
.Y(n_7839)
);

CKINVDCx6p67_ASAP7_75t_R g7840 ( 
.A(n_6881),
.Y(n_7840)
);

BUFx3_ASAP7_75t_L g7841 ( 
.A(n_5826),
.Y(n_7841)
);

OR2x2_ASAP7_75t_L g7842 ( 
.A(n_6525),
.B(n_5049),
.Y(n_7842)
);

NAND2x1p5_ASAP7_75t_L g7843 ( 
.A(n_6481),
.B(n_5700),
.Y(n_7843)
);

NOR2xp67_ASAP7_75t_L g7844 ( 
.A(n_5761),
.B(n_5124),
.Y(n_7844)
);

AOI21xp5_ASAP7_75t_L g7845 ( 
.A1(n_6061),
.A2(n_5632),
.B(n_5630),
.Y(n_7845)
);

INVx2_ASAP7_75t_SL g7846 ( 
.A(n_6083),
.Y(n_7846)
);

NAND2xp5_ASAP7_75t_L g7847 ( 
.A(n_6392),
.B(n_5021),
.Y(n_7847)
);

NOR2xp33_ASAP7_75t_SL g7848 ( 
.A(n_5866),
.B(n_5190),
.Y(n_7848)
);

AOI22xp5_ASAP7_75t_L g7849 ( 
.A1(n_6378),
.A2(n_5557),
.B1(n_5551),
.B2(n_5720),
.Y(n_7849)
);

AOI22xp33_ASAP7_75t_L g7850 ( 
.A1(n_5921),
.A2(n_5035),
.B1(n_5038),
.B2(n_5021),
.Y(n_7850)
);

AO21x1_ASAP7_75t_L g7851 ( 
.A1(n_6244),
.A2(n_5054),
.B(n_5049),
.Y(n_7851)
);

OAI22xp5_ASAP7_75t_L g7852 ( 
.A1(n_5796),
.A2(n_5369),
.B1(n_5418),
.B2(n_5308),
.Y(n_7852)
);

AOI21xp5_ASAP7_75t_L g7853 ( 
.A1(n_6052),
.A2(n_6061),
.B(n_6501),
.Y(n_7853)
);

INVx2_ASAP7_75t_SL g7854 ( 
.A(n_6115),
.Y(n_7854)
);

BUFx2_ASAP7_75t_L g7855 ( 
.A(n_6908),
.Y(n_7855)
);

BUFx12f_ASAP7_75t_L g7856 ( 
.A(n_6109),
.Y(n_7856)
);

INVx2_ASAP7_75t_SL g7857 ( 
.A(n_6115),
.Y(n_7857)
);

INVxp67_ASAP7_75t_L g7858 ( 
.A(n_6534),
.Y(n_7858)
);

AOI22x1_ASAP7_75t_L g7859 ( 
.A1(n_6052),
.A2(n_5588),
.B1(n_5594),
.B2(n_5560),
.Y(n_7859)
);

OA21x2_ASAP7_75t_L g7860 ( 
.A1(n_6907),
.A2(n_5679),
.B(n_5055),
.Y(n_7860)
);

CKINVDCx5p33_ASAP7_75t_R g7861 ( 
.A(n_6109),
.Y(n_7861)
);

BUFx2_ASAP7_75t_L g7862 ( 
.A(n_6908),
.Y(n_7862)
);

OAI22xp5_ASAP7_75t_L g7863 ( 
.A1(n_5829),
.A2(n_5369),
.B1(n_5418),
.B2(n_5308),
.Y(n_7863)
);

AOI221xp5_ASAP7_75t_L g7864 ( 
.A1(n_6200),
.A2(n_5039),
.B1(n_5042),
.B2(n_5038),
.C(n_5035),
.Y(n_7864)
);

NAND2xp5_ASAP7_75t_L g7865 ( 
.A(n_6401),
.B(n_5038),
.Y(n_7865)
);

INVx5_ASAP7_75t_L g7866 ( 
.A(n_6221),
.Y(n_7866)
);

HB1xp67_ASAP7_75t_L g7867 ( 
.A(n_6531),
.Y(n_7867)
);

BUFx4_ASAP7_75t_SL g7868 ( 
.A(n_6235),
.Y(n_7868)
);

NAND2xp5_ASAP7_75t_L g7869 ( 
.A(n_6401),
.B(n_6439),
.Y(n_7869)
);

AOI21x1_ASAP7_75t_L g7870 ( 
.A1(n_6781),
.A2(n_5604),
.B(n_5615),
.Y(n_7870)
);

INVx5_ASAP7_75t_L g7871 ( 
.A(n_6221),
.Y(n_7871)
);

AOI22xp33_ASAP7_75t_L g7872 ( 
.A1(n_5921),
.A2(n_5042),
.B1(n_5045),
.B2(n_5039),
.Y(n_7872)
);

OAI22xp5_ASAP7_75t_L g7873 ( 
.A1(n_5829),
.A2(n_5369),
.B1(n_5418),
.B2(n_5308),
.Y(n_7873)
);

NOR2xp33_ASAP7_75t_L g7874 ( 
.A(n_6013),
.B(n_5557),
.Y(n_7874)
);

AOI22xp33_ASAP7_75t_L g7875 ( 
.A1(n_6013),
.A2(n_5042),
.B1(n_5045),
.B2(n_5039),
.Y(n_7875)
);

NAND2x1p5_ASAP7_75t_L g7876 ( 
.A(n_6389),
.B(n_5124),
.Y(n_7876)
);

BUFx3_ASAP7_75t_L g7877 ( 
.A(n_5836),
.Y(n_7877)
);

NAND2xp5_ASAP7_75t_L g7878 ( 
.A(n_6439),
.B(n_5045),
.Y(n_7878)
);

AOI22xp5_ASAP7_75t_L g7879 ( 
.A1(n_6580),
.A2(n_5720),
.B1(n_4522),
.B2(n_4528),
.Y(n_7879)
);

NOR2xp33_ASAP7_75t_L g7880 ( 
.A(n_6015),
.B(n_6028),
.Y(n_7880)
);

INVx2_ASAP7_75t_SL g7881 ( 
.A(n_6115),
.Y(n_7881)
);

NAND2xp5_ASAP7_75t_L g7882 ( 
.A(n_6200),
.B(n_6629),
.Y(n_7882)
);

O2A1O1Ixp33_ASAP7_75t_L g7883 ( 
.A1(n_6123),
.A2(n_5055),
.B(n_5058),
.C(n_5054),
.Y(n_7883)
);

NAND2xp5_ASAP7_75t_L g7884 ( 
.A(n_6629),
.B(n_6639),
.Y(n_7884)
);

AOI21xp5_ASAP7_75t_L g7885 ( 
.A1(n_6501),
.A2(n_5632),
.B(n_5630),
.Y(n_7885)
);

BUFx2_ASAP7_75t_L g7886 ( 
.A(n_6908),
.Y(n_7886)
);

INVx2_ASAP7_75t_SL g7887 ( 
.A(n_6115),
.Y(n_7887)
);

INVx1_ASAP7_75t_SL g7888 ( 
.A(n_6916),
.Y(n_7888)
);

BUFx6f_ASAP7_75t_L g7889 ( 
.A(n_6634),
.Y(n_7889)
);

INVx6_ASAP7_75t_L g7890 ( 
.A(n_5893),
.Y(n_7890)
);

OAI22xp33_ASAP7_75t_L g7891 ( 
.A1(n_6580),
.A2(n_5124),
.B1(n_5243),
.B2(n_5190),
.Y(n_7891)
);

AOI222xp33_ASAP7_75t_L g7892 ( 
.A1(n_6015),
.A2(n_5060),
.B1(n_5052),
.B2(n_5063),
.C1(n_5056),
.C2(n_5050),
.Y(n_7892)
);

AOI21xp5_ASAP7_75t_L g7893 ( 
.A1(n_6502),
.A2(n_5632),
.B(n_5630),
.Y(n_7893)
);

BUFx3_ASAP7_75t_L g7894 ( 
.A(n_5836),
.Y(n_7894)
);

OAI321xp33_ASAP7_75t_L g7895 ( 
.A1(n_6181),
.A2(n_5367),
.A3(n_5364),
.B1(n_5368),
.B2(n_5365),
.C(n_5359),
.Y(n_7895)
);

AOI21xp5_ASAP7_75t_L g7896 ( 
.A1(n_6502),
.A2(n_5632),
.B(n_5630),
.Y(n_7896)
);

INVxp67_ASAP7_75t_L g7897 ( 
.A(n_6561),
.Y(n_7897)
);

OAI21x1_ASAP7_75t_L g7898 ( 
.A1(n_6724),
.A2(n_4517),
.B(n_4516),
.Y(n_7898)
);

CKINVDCx20_ASAP7_75t_R g7899 ( 
.A(n_6346),
.Y(n_7899)
);

AOI22xp33_ASAP7_75t_L g7900 ( 
.A1(n_6028),
.A2(n_5052),
.B1(n_5056),
.B2(n_5050),
.Y(n_7900)
);

INVx1_ASAP7_75t_SL g7901 ( 
.A(n_6916),
.Y(n_7901)
);

NOR2xp33_ASAP7_75t_L g7902 ( 
.A(n_6049),
.B(n_5050),
.Y(n_7902)
);

CKINVDCx5p33_ASAP7_75t_R g7903 ( 
.A(n_6109),
.Y(n_7903)
);

BUFx2_ASAP7_75t_L g7904 ( 
.A(n_6916),
.Y(n_7904)
);

A2O1A1Ixp33_ASAP7_75t_L g7905 ( 
.A1(n_6542),
.A2(n_4503),
.B(n_4599),
.C(n_4522),
.Y(n_7905)
);

INVx3_ASAP7_75t_SL g7906 ( 
.A(n_6630),
.Y(n_7906)
);

CKINVDCx5p33_ASAP7_75t_R g7907 ( 
.A(n_6349),
.Y(n_7907)
);

CKINVDCx6p67_ASAP7_75t_R g7908 ( 
.A(n_6881),
.Y(n_7908)
);

INVx5_ASAP7_75t_L g7909 ( 
.A(n_6221),
.Y(n_7909)
);

NAND2xp5_ASAP7_75t_L g7910 ( 
.A(n_6639),
.B(n_5052),
.Y(n_7910)
);

INVx1_ASAP7_75t_SL g7911 ( 
.A(n_5813),
.Y(n_7911)
);

INVxp67_ASAP7_75t_SL g7912 ( 
.A(n_6877),
.Y(n_7912)
);

BUFx2_ASAP7_75t_L g7913 ( 
.A(n_5919),
.Y(n_7913)
);

A2O1A1Ixp33_ASAP7_75t_L g7914 ( 
.A1(n_6542),
.A2(n_4503),
.B(n_4599),
.C(n_4522),
.Y(n_7914)
);

BUFx8_ASAP7_75t_L g7915 ( 
.A(n_6057),
.Y(n_7915)
);

NAND2xp5_ASAP7_75t_L g7916 ( 
.A(n_6641),
.B(n_5056),
.Y(n_7916)
);

CKINVDCx20_ASAP7_75t_R g7917 ( 
.A(n_6785),
.Y(n_7917)
);

BUFx6f_ASAP7_75t_L g7918 ( 
.A(n_6634),
.Y(n_7918)
);

INVx2_ASAP7_75t_SL g7919 ( 
.A(n_6115),
.Y(n_7919)
);

OAI21x1_ASAP7_75t_L g7920 ( 
.A1(n_6724),
.A2(n_4517),
.B(n_4516),
.Y(n_7920)
);

OR2x2_ASAP7_75t_L g7921 ( 
.A(n_6559),
.B(n_5058),
.Y(n_7921)
);

AOI21x1_ASAP7_75t_L g7922 ( 
.A1(n_6781),
.A2(n_5604),
.B(n_5615),
.Y(n_7922)
);

OAI22xp5_ASAP7_75t_L g7923 ( 
.A1(n_6049),
.A2(n_5369),
.B1(n_5418),
.B2(n_5308),
.Y(n_7923)
);

HB1xp67_ASAP7_75t_L g7924 ( 
.A(n_6531),
.Y(n_7924)
);

BUFx2_ASAP7_75t_L g7925 ( 
.A(n_5919),
.Y(n_7925)
);

O2A1O1Ixp33_ASAP7_75t_L g7926 ( 
.A1(n_6123),
.A2(n_5065),
.B(n_5070),
.C(n_5064),
.Y(n_7926)
);

INVx4_ASAP7_75t_L g7927 ( 
.A(n_6588),
.Y(n_7927)
);

AOI21xp5_ASAP7_75t_L g7928 ( 
.A1(n_6508),
.A2(n_5632),
.B(n_5630),
.Y(n_7928)
);

CKINVDCx20_ASAP7_75t_R g7929 ( 
.A(n_6785),
.Y(n_7929)
);

AO32x2_ASAP7_75t_L g7930 ( 
.A1(n_6616),
.A2(n_4658),
.A3(n_4720),
.B1(n_4624),
.B2(n_4599),
.Y(n_7930)
);

INVx3_ASAP7_75t_SL g7931 ( 
.A(n_6672),
.Y(n_7931)
);

CKINVDCx16_ASAP7_75t_R g7932 ( 
.A(n_6412),
.Y(n_7932)
);

INVx1_ASAP7_75t_SL g7933 ( 
.A(n_5813),
.Y(n_7933)
);

NAND2xp5_ASAP7_75t_SL g7934 ( 
.A(n_5735),
.B(n_4508),
.Y(n_7934)
);

BUFx2_ASAP7_75t_L g7935 ( 
.A(n_5949),
.Y(n_7935)
);

AOI22xp5_ASAP7_75t_L g7936 ( 
.A1(n_6051),
.A2(n_5720),
.B1(n_4505),
.B2(n_4528),
.Y(n_7936)
);

AOI21xp5_ASAP7_75t_L g7937 ( 
.A1(n_6508),
.A2(n_6555),
.B(n_6517),
.Y(n_7937)
);

OR2x2_ASAP7_75t_L g7938 ( 
.A(n_6559),
.B(n_5064),
.Y(n_7938)
);

INVx3_ASAP7_75t_SL g7939 ( 
.A(n_6672),
.Y(n_7939)
);

INVx1_ASAP7_75t_SL g7940 ( 
.A(n_5813),
.Y(n_7940)
);

HB1xp67_ASAP7_75t_L g7941 ( 
.A(n_6535),
.Y(n_7941)
);

AOI22xp33_ASAP7_75t_L g7942 ( 
.A1(n_6051),
.A2(n_5063),
.B1(n_5073),
.B2(n_5060),
.Y(n_7942)
);

NAND2xp5_ASAP7_75t_L g7943 ( 
.A(n_6641),
.B(n_5060),
.Y(n_7943)
);

NOR2xp33_ASAP7_75t_L g7944 ( 
.A(n_5863),
.B(n_5063),
.Y(n_7944)
);

HB1xp67_ASAP7_75t_L g7945 ( 
.A(n_6535),
.Y(n_7945)
);

CKINVDCx11_ASAP7_75t_R g7946 ( 
.A(n_6349),
.Y(n_7946)
);

AOI21xp5_ASAP7_75t_L g7947 ( 
.A1(n_6555),
.A2(n_5630),
.B(n_5583),
.Y(n_7947)
);

AOI21x1_ASAP7_75t_L g7948 ( 
.A1(n_6726),
.A2(n_5706),
.B(n_5399),
.Y(n_7948)
);

INVx2_ASAP7_75t_SL g7949 ( 
.A(n_6117),
.Y(n_7949)
);

BUFx3_ASAP7_75t_L g7950 ( 
.A(n_5836),
.Y(n_7950)
);

AOI22xp33_ASAP7_75t_L g7951 ( 
.A1(n_6296),
.A2(n_5075),
.B1(n_5081),
.B2(n_5073),
.Y(n_7951)
);

NAND2xp5_ASAP7_75t_L g7952 ( 
.A(n_6646),
.B(n_6748),
.Y(n_7952)
);

OAI22xp5_ASAP7_75t_SL g7953 ( 
.A1(n_6450),
.A2(n_5682),
.B1(n_5684),
.B2(n_5594),
.Y(n_7953)
);

OR2x2_ASAP7_75t_SL g7954 ( 
.A(n_6895),
.B(n_4508),
.Y(n_7954)
);

INVx2_ASAP7_75t_SL g7955 ( 
.A(n_6117),
.Y(n_7955)
);

CKINVDCx5p33_ASAP7_75t_R g7956 ( 
.A(n_6349),
.Y(n_7956)
);

BUFx6f_ASAP7_75t_L g7957 ( 
.A(n_6634),
.Y(n_7957)
);

AOI21xp5_ASAP7_75t_L g7958 ( 
.A1(n_6555),
.A2(n_5583),
.B(n_5576),
.Y(n_7958)
);

NOR2xp33_ASAP7_75t_L g7959 ( 
.A(n_5863),
.B(n_5073),
.Y(n_7959)
);

NAND2xp5_ASAP7_75t_L g7960 ( 
.A(n_6646),
.B(n_5075),
.Y(n_7960)
);

AOI21xp5_ASAP7_75t_L g7961 ( 
.A1(n_6555),
.A2(n_5614),
.B(n_5611),
.Y(n_7961)
);

INVx1_ASAP7_75t_SL g7962 ( 
.A(n_5847),
.Y(n_7962)
);

NAND2xp5_ASAP7_75t_L g7963 ( 
.A(n_6748),
.B(n_5075),
.Y(n_7963)
);

INVxp67_ASAP7_75t_SL g7964 ( 
.A(n_6877),
.Y(n_7964)
);

O2A1O1Ixp5_ASAP7_75t_L g7965 ( 
.A1(n_6292),
.A2(n_5087),
.B(n_5093),
.C(n_5081),
.Y(n_7965)
);

BUFx2_ASAP7_75t_L g7966 ( 
.A(n_5949),
.Y(n_7966)
);

AND2x2_ASAP7_75t_L g7967 ( 
.A(n_6489),
.B(n_4995),
.Y(n_7967)
);

NAND2xp5_ASAP7_75t_L g7968 ( 
.A(n_6763),
.B(n_5081),
.Y(n_7968)
);

OAI22xp5_ASAP7_75t_L g7969 ( 
.A1(n_5856),
.A2(n_5418),
.B1(n_5369),
.B2(n_5070),
.Y(n_7969)
);

NAND2xp5_ASAP7_75t_L g7970 ( 
.A(n_6763),
.B(n_5087),
.Y(n_7970)
);

NOR2xp33_ASAP7_75t_L g7971 ( 
.A(n_5747),
.B(n_5743),
.Y(n_7971)
);

OAI22xp5_ASAP7_75t_L g7972 ( 
.A1(n_5856),
.A2(n_5418),
.B1(n_5076),
.B2(n_5085),
.Y(n_7972)
);

INVxp67_ASAP7_75t_L g7973 ( 
.A(n_6561),
.Y(n_7973)
);

OAI221xp5_ASAP7_75t_L g7974 ( 
.A1(n_6153),
.A2(n_5094),
.B1(n_5097),
.B2(n_5093),
.C(n_5087),
.Y(n_7974)
);

BUFx4f_ASAP7_75t_L g7975 ( 
.A(n_6385),
.Y(n_7975)
);

BUFx6f_ASAP7_75t_L g7976 ( 
.A(n_6032),
.Y(n_7976)
);

OAI21xp33_ASAP7_75t_SL g7977 ( 
.A1(n_6181),
.A2(n_4658),
.B(n_4624),
.Y(n_7977)
);

CKINVDCx16_ASAP7_75t_R g7978 ( 
.A(n_6412),
.Y(n_7978)
);

BUFx4f_ASAP7_75t_L g7979 ( 
.A(n_6385),
.Y(n_7979)
);

AO21x1_ASAP7_75t_L g7980 ( 
.A1(n_6244),
.A2(n_5076),
.B(n_5065),
.Y(n_7980)
);

OAI22xp33_ASAP7_75t_L g7981 ( 
.A1(n_6532),
.A2(n_5124),
.B1(n_5243),
.B2(n_5190),
.Y(n_7981)
);

NAND2xp5_ASAP7_75t_L g7982 ( 
.A(n_6796),
.B(n_6815),
.Y(n_7982)
);

OR2x2_ASAP7_75t_L g7983 ( 
.A(n_5747),
.B(n_5085),
.Y(n_7983)
);

INVx2_ASAP7_75t_SL g7984 ( 
.A(n_6117),
.Y(n_7984)
);

NAND2xp5_ASAP7_75t_L g7985 ( 
.A(n_6796),
.B(n_5093),
.Y(n_7985)
);

AO21x1_ASAP7_75t_L g7986 ( 
.A1(n_6178),
.A2(n_5089),
.B(n_5086),
.Y(n_7986)
);

NOR2xp33_ASAP7_75t_L g7987 ( 
.A(n_5747),
.B(n_5743),
.Y(n_7987)
);

NAND2xp5_ASAP7_75t_L g7988 ( 
.A(n_6815),
.B(n_5094),
.Y(n_7988)
);

NOR2x1_ASAP7_75t_L g7989 ( 
.A(n_5739),
.B(n_5094),
.Y(n_7989)
);

AOI22xp5_ASAP7_75t_L g7990 ( 
.A1(n_6374),
.A2(n_5720),
.B1(n_4522),
.B2(n_4528),
.Y(n_7990)
);

NAND2xp5_ASAP7_75t_SL g7991 ( 
.A(n_6728),
.B(n_4518),
.Y(n_7991)
);

HB1xp67_ASAP7_75t_L g7992 ( 
.A(n_6551),
.Y(n_7992)
);

AOI22xp33_ASAP7_75t_L g7993 ( 
.A1(n_6296),
.A2(n_5099),
.B1(n_5110),
.B2(n_5097),
.Y(n_7993)
);

AOI21xp5_ASAP7_75t_L g7994 ( 
.A1(n_6555),
.A2(n_5614),
.B(n_5611),
.Y(n_7994)
);

BUFx6f_ASAP7_75t_L g7995 ( 
.A(n_6032),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_L g7996 ( 
.A(n_6833),
.B(n_5097),
.Y(n_7996)
);

OAI22xp33_ASAP7_75t_L g7997 ( 
.A1(n_6532),
.A2(n_5124),
.B1(n_5243),
.B2(n_5190),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_6833),
.B(n_5099),
.Y(n_7998)
);

BUFx12f_ASAP7_75t_L g7999 ( 
.A(n_6364),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_L g8000 ( 
.A(n_6839),
.B(n_5099),
.Y(n_8000)
);

OAI22xp33_ASAP7_75t_L g8001 ( 
.A1(n_5977),
.A2(n_5124),
.B1(n_5245),
.B2(n_5243),
.Y(n_8001)
);

BUFx6f_ASAP7_75t_L g8002 ( 
.A(n_6032),
.Y(n_8002)
);

OR2x2_ASAP7_75t_L g8003 ( 
.A(n_6791),
.B(n_5086),
.Y(n_8003)
);

BUFx12f_ASAP7_75t_L g8004 ( 
.A(n_6364),
.Y(n_8004)
);

OAI22xp5_ASAP7_75t_L g8005 ( 
.A1(n_6327),
.A2(n_5095),
.B1(n_5102),
.B2(n_5089),
.Y(n_8005)
);

OR2x2_ASAP7_75t_L g8006 ( 
.A(n_6791),
.B(n_5095),
.Y(n_8006)
);

AOI22xp33_ASAP7_75t_L g8007 ( 
.A1(n_6302),
.A2(n_5113),
.B1(n_5110),
.B2(n_5245),
.Y(n_8007)
);

AOI21xp5_ASAP7_75t_L g8008 ( 
.A1(n_6555),
.A2(n_5614),
.B(n_4658),
.Y(n_8008)
);

AOI22xp5_ASAP7_75t_L g8009 ( 
.A1(n_6374),
.A2(n_5720),
.B1(n_4522),
.B2(n_4528),
.Y(n_8009)
);

AOI21xp5_ASAP7_75t_L g8010 ( 
.A1(n_6555),
.A2(n_4720),
.B(n_4624),
.Y(n_8010)
);

INVxp67_ASAP7_75t_L g8011 ( 
.A(n_6427),
.Y(n_8011)
);

NAND2x1p5_ASAP7_75t_L g8012 ( 
.A(n_6389),
.B(n_5124),
.Y(n_8012)
);

NAND2xp5_ASAP7_75t_SL g8013 ( 
.A(n_6728),
.B(n_4518),
.Y(n_8013)
);

BUFx12f_ASAP7_75t_L g8014 ( 
.A(n_6364),
.Y(n_8014)
);

OAI22xp33_ASAP7_75t_L g8015 ( 
.A1(n_5977),
.A2(n_5124),
.B1(n_5245),
.B2(n_4518),
.Y(n_8015)
);

OA21x2_ASAP7_75t_L g8016 ( 
.A1(n_6726),
.A2(n_5103),
.B(n_5102),
.Y(n_8016)
);

AOI21xp5_ASAP7_75t_L g8017 ( 
.A1(n_6512),
.A2(n_4720),
.B(n_5603),
.Y(n_8017)
);

INVx2_ASAP7_75t_SL g8018 ( 
.A(n_6117),
.Y(n_8018)
);

NAND2x1p5_ASAP7_75t_L g8019 ( 
.A(n_6389),
.B(n_5431),
.Y(n_8019)
);

AOI21xp33_ASAP7_75t_L g8020 ( 
.A1(n_6153),
.A2(n_5113),
.B(n_5110),
.Y(n_8020)
);

BUFx6f_ASAP7_75t_L g8021 ( 
.A(n_6032),
.Y(n_8021)
);

NAND2xp5_ASAP7_75t_SL g8022 ( 
.A(n_6692),
.B(n_4518),
.Y(n_8022)
);

AOI22xp5_ASAP7_75t_L g8023 ( 
.A1(n_6122),
.A2(n_5720),
.B1(n_4528),
.B2(n_4556),
.Y(n_8023)
);

OAI22xp5_ASAP7_75t_L g8024 ( 
.A1(n_6327),
.A2(n_5104),
.B1(n_5107),
.B2(n_5103),
.Y(n_8024)
);

BUFx2_ASAP7_75t_L g8025 ( 
.A(n_5847),
.Y(n_8025)
);

NAND2xp5_ASAP7_75t_L g8026 ( 
.A(n_6839),
.B(n_5113),
.Y(n_8026)
);

BUFx3_ASAP7_75t_L g8027 ( 
.A(n_5836),
.Y(n_8027)
);

BUFx2_ASAP7_75t_L g8028 ( 
.A(n_5847),
.Y(n_8028)
);

AOI21xp5_ASAP7_75t_L g8029 ( 
.A1(n_6512),
.A2(n_5612),
.B(n_5603),
.Y(n_8029)
);

NAND2xp5_ASAP7_75t_L g8030 ( 
.A(n_6842),
.B(n_5104),
.Y(n_8030)
);

HAxp5_ASAP7_75t_L g8031 ( 
.A(n_5895),
.B(n_5273),
.CON(n_8031),
.SN(n_8031)
);

HB1xp67_ASAP7_75t_L g8032 ( 
.A(n_6551),
.Y(n_8032)
);

NOR2xp67_ASAP7_75t_L g8033 ( 
.A(n_5761),
.B(n_6105),
.Y(n_8033)
);

OAI21xp33_ASAP7_75t_L g8034 ( 
.A1(n_5755),
.A2(n_5112),
.B(n_5107),
.Y(n_8034)
);

NAND2xp5_ASAP7_75t_L g8035 ( 
.A(n_6842),
.B(n_5112),
.Y(n_8035)
);

OAI22xp5_ASAP7_75t_L g8036 ( 
.A1(n_6327),
.A2(n_5123),
.B1(n_5126),
.B2(n_5114),
.Y(n_8036)
);

INVx2_ASAP7_75t_SL g8037 ( 
.A(n_6117),
.Y(n_8037)
);

AND2x2_ASAP7_75t_L g8038 ( 
.A(n_6489),
.B(n_4995),
.Y(n_8038)
);

AOI22xp33_ASAP7_75t_L g8039 ( 
.A1(n_6302),
.A2(n_5245),
.B1(n_5713),
.B2(n_5712),
.Y(n_8039)
);

HB1xp67_ASAP7_75t_L g8040 ( 
.A(n_6556),
.Y(n_8040)
);

AOI21xp5_ASAP7_75t_L g8041 ( 
.A1(n_6517),
.A2(n_5612),
.B(n_5603),
.Y(n_8041)
);

INVx2_ASAP7_75t_SL g8042 ( 
.A(n_6118),
.Y(n_8042)
);

OAI22xp5_ASAP7_75t_L g8043 ( 
.A1(n_5733),
.A2(n_5123),
.B1(n_5126),
.B2(n_5114),
.Y(n_8043)
);

CKINVDCx11_ASAP7_75t_R g8044 ( 
.A(n_6568),
.Y(n_8044)
);

BUFx2_ASAP7_75t_L g8045 ( 
.A(n_5857),
.Y(n_8045)
);

AOI22xp33_ASAP7_75t_L g8046 ( 
.A1(n_5754),
.A2(n_5713),
.B1(n_5723),
.B2(n_5712),
.Y(n_8046)
);

A2O1A1Ixp33_ASAP7_75t_L g8047 ( 
.A1(n_5913),
.A2(n_4556),
.B(n_4604),
.C(n_4505),
.Y(n_8047)
);

INVx3_ASAP7_75t_SL g8048 ( 
.A(n_6672),
.Y(n_8048)
);

AOI22xp5_ASAP7_75t_L g8049 ( 
.A1(n_6122),
.A2(n_5720),
.B1(n_4556),
.B2(n_4604),
.Y(n_8049)
);

CKINVDCx16_ASAP7_75t_R g8050 ( 
.A(n_6423),
.Y(n_8050)
);

OR2x2_ASAP7_75t_L g8051 ( 
.A(n_6791),
.B(n_5128),
.Y(n_8051)
);

NAND2xp5_ASAP7_75t_L g8052 ( 
.A(n_6844),
.B(n_5128),
.Y(n_8052)
);

CKINVDCx5p33_ASAP7_75t_R g8053 ( 
.A(n_6568),
.Y(n_8053)
);

BUFx2_ASAP7_75t_L g8054 ( 
.A(n_5857),
.Y(n_8054)
);

AO221x2_ASAP7_75t_L g8055 ( 
.A1(n_6450),
.A2(n_6464),
.B1(n_5733),
.B2(n_5807),
.C(n_5810),
.Y(n_8055)
);

BUFx3_ASAP7_75t_L g8056 ( 
.A(n_5915),
.Y(n_8056)
);

BUFx3_ASAP7_75t_L g8057 ( 
.A(n_5915),
.Y(n_8057)
);

CKINVDCx5p33_ASAP7_75t_R g8058 ( 
.A(n_6568),
.Y(n_8058)
);

INVx1_ASAP7_75t_SL g8059 ( 
.A(n_5857),
.Y(n_8059)
);

HB1xp67_ASAP7_75t_L g8060 ( 
.A(n_6556),
.Y(n_8060)
);

NAND2xp5_ASAP7_75t_L g8061 ( 
.A(n_6844),
.B(n_4621),
.Y(n_8061)
);

AND2x2_ASAP7_75t_L g8062 ( 
.A(n_6489),
.B(n_4995),
.Y(n_8062)
);

CKINVDCx20_ASAP7_75t_R g8063 ( 
.A(n_6275),
.Y(n_8063)
);

BUFx3_ASAP7_75t_L g8064 ( 
.A(n_5915),
.Y(n_8064)
);

OAI22xp5_ASAP7_75t_L g8065 ( 
.A1(n_6464),
.A2(n_5431),
.B1(n_5162),
.B2(n_5174),
.Y(n_8065)
);

HB1xp67_ASAP7_75t_L g8066 ( 
.A(n_6585),
.Y(n_8066)
);

BUFx12f_ASAP7_75t_L g8067 ( 
.A(n_6596),
.Y(n_8067)
);

INVx2_ASAP7_75t_SL g8068 ( 
.A(n_6118),
.Y(n_8068)
);

BUFx6f_ASAP7_75t_L g8069 ( 
.A(n_6607),
.Y(n_8069)
);

INVx4_ASAP7_75t_L g8070 ( 
.A(n_6607),
.Y(n_8070)
);

BUFx12f_ASAP7_75t_L g8071 ( 
.A(n_6596),
.Y(n_8071)
);

CKINVDCx6p67_ASAP7_75t_R g8072 ( 
.A(n_6895),
.Y(n_8072)
);

AOI21xp5_ASAP7_75t_L g8073 ( 
.A1(n_6806),
.A2(n_5622),
.B(n_5612),
.Y(n_8073)
);

AND2x2_ASAP7_75t_L g8074 ( 
.A(n_6287),
.B(n_4998),
.Y(n_8074)
);

O2A1O1Ixp33_ASAP7_75t_SL g8075 ( 
.A1(n_5895),
.A2(n_5357),
.B(n_5694),
.C(n_5454),
.Y(n_8075)
);

BUFx3_ASAP7_75t_L g8076 ( 
.A(n_5915),
.Y(n_8076)
);

NAND2x1_ASAP7_75t_L g8077 ( 
.A(n_6672),
.B(n_4516),
.Y(n_8077)
);

BUFx2_ASAP7_75t_L g8078 ( 
.A(n_5903),
.Y(n_8078)
);

INVx3_ASAP7_75t_SL g8079 ( 
.A(n_6672),
.Y(n_8079)
);

BUFx3_ASAP7_75t_L g8080 ( 
.A(n_5976),
.Y(n_8080)
);

AND2x2_ASAP7_75t_L g8081 ( 
.A(n_6287),
.B(n_6445),
.Y(n_8081)
);

OR2x2_ASAP7_75t_L g8082 ( 
.A(n_5752),
.B(n_5372),
.Y(n_8082)
);

INVx1_ASAP7_75t_SL g8083 ( 
.A(n_5903),
.Y(n_8083)
);

AOI22xp5_ASAP7_75t_L g8084 ( 
.A1(n_5737),
.A2(n_5720),
.B1(n_4556),
.B2(n_4604),
.Y(n_8084)
);

AOI222xp33_ASAP7_75t_L g8085 ( 
.A1(n_5862),
.A2(n_5684),
.B1(n_5699),
.B2(n_5682),
.C1(n_5372),
.C2(n_5720),
.Y(n_8085)
);

A2O1A1Ixp33_ASAP7_75t_SL g8086 ( 
.A1(n_6674),
.A2(n_5680),
.B(n_5685),
.C(n_5673),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_6088),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_6088),
.Y(n_8088)
);

AND2x2_ASAP7_75t_L g8089 ( 
.A(n_6287),
.B(n_4998),
.Y(n_8089)
);

INVx2_ASAP7_75t_SL g8090 ( 
.A(n_6118),
.Y(n_8090)
);

BUFx8_ASAP7_75t_L g8091 ( 
.A(n_6057),
.Y(n_8091)
);

AOI22xp5_ASAP7_75t_L g8092 ( 
.A1(n_5737),
.A2(n_5720),
.B1(n_4556),
.B2(n_4604),
.Y(n_8092)
);

INVx2_ASAP7_75t_SL g8093 ( 
.A(n_6118),
.Y(n_8093)
);

INVx4_ASAP7_75t_L g8094 ( 
.A(n_6613),
.Y(n_8094)
);

NAND2xp5_ASAP7_75t_L g8095 ( 
.A(n_6854),
.B(n_4621),
.Y(n_8095)
);

AOI21xp33_ASAP7_75t_L g8096 ( 
.A1(n_6043),
.A2(n_5672),
.B(n_5140),
.Y(n_8096)
);

NAND2xp5_ASAP7_75t_L g8097 ( 
.A(n_6854),
.B(n_4621),
.Y(n_8097)
);

INVx2_ASAP7_75t_SL g8098 ( 
.A(n_6118),
.Y(n_8098)
);

AND2x2_ASAP7_75t_L g8099 ( 
.A(n_6445),
.B(n_4998),
.Y(n_8099)
);

OAI22xp5_ASAP7_75t_L g8100 ( 
.A1(n_6570),
.A2(n_5431),
.B1(n_5162),
.B2(n_5174),
.Y(n_8100)
);

BUFx2_ASAP7_75t_L g8101 ( 
.A(n_5903),
.Y(n_8101)
);

AOI21xp5_ASAP7_75t_L g8102 ( 
.A1(n_6806),
.A2(n_5634),
.B(n_5622),
.Y(n_8102)
);

AND2x2_ASAP7_75t_L g8103 ( 
.A(n_6445),
.B(n_4998),
.Y(n_8103)
);

BUFx3_ASAP7_75t_L g8104 ( 
.A(n_5976),
.Y(n_8104)
);

NOR2xp33_ASAP7_75t_L g8105 ( 
.A(n_5832),
.B(n_5627),
.Y(n_8105)
);

AOI22xp33_ASAP7_75t_L g8106 ( 
.A1(n_5754),
.A2(n_5713),
.B1(n_5723),
.B2(n_5712),
.Y(n_8106)
);

BUFx2_ASAP7_75t_L g8107 ( 
.A(n_5909),
.Y(n_8107)
);

INVx2_ASAP7_75t_SL g8108 ( 
.A(n_6145),
.Y(n_8108)
);

BUFx2_ASAP7_75t_L g8109 ( 
.A(n_5909),
.Y(n_8109)
);

OR2x6_ASAP7_75t_L g8110 ( 
.A(n_6640),
.B(n_6270),
.Y(n_8110)
);

INVx1_ASAP7_75t_L g8111 ( 
.A(n_6090),
.Y(n_8111)
);

AOI221xp5_ASAP7_75t_L g8112 ( 
.A1(n_5727),
.A2(n_5372),
.B1(n_5174),
.B2(n_5176),
.C(n_5169),
.Y(n_8112)
);

AOI22xp5_ASAP7_75t_L g8113 ( 
.A1(n_5862),
.A2(n_4556),
.B1(n_4604),
.B2(n_4505),
.Y(n_8113)
);

AND2x2_ASAP7_75t_L g8114 ( 
.A(n_6455),
.B(n_5024),
.Y(n_8114)
);

INVx1_ASAP7_75t_SL g8115 ( 
.A(n_5909),
.Y(n_8115)
);

CKINVDCx6p67_ASAP7_75t_R g8116 ( 
.A(n_6901),
.Y(n_8116)
);

BUFx2_ASAP7_75t_L g8117 ( 
.A(n_5910),
.Y(n_8117)
);

NAND2x1p5_ASAP7_75t_L g8118 ( 
.A(n_6389),
.B(n_6416),
.Y(n_8118)
);

AND2x2_ASAP7_75t_SL g8119 ( 
.A(n_5837),
.B(n_4505),
.Y(n_8119)
);

NOR3xp33_ASAP7_75t_L g8120 ( 
.A(n_6292),
.B(n_5143),
.C(n_5138),
.Y(n_8120)
);

NAND2xp5_ASAP7_75t_L g8121 ( 
.A(n_6867),
.B(n_4621),
.Y(n_8121)
);

BUFx2_ASAP7_75t_L g8122 ( 
.A(n_5910),
.Y(n_8122)
);

AND2x2_ASAP7_75t_L g8123 ( 
.A(n_6455),
.B(n_5024),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_L g8124 ( 
.A(n_6867),
.B(n_4629),
.Y(n_8124)
);

OR2x2_ASAP7_75t_L g8125 ( 
.A(n_5752),
.B(n_5140),
.Y(n_8125)
);

O2A1O1Ixp33_ASAP7_75t_L g8126 ( 
.A1(n_5924),
.A2(n_6438),
.B(n_5913),
.C(n_5727),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_6208),
.B(n_4629),
.Y(n_8127)
);

O2A1O1Ixp33_ASAP7_75t_SL g8128 ( 
.A1(n_6404),
.A2(n_5694),
.B(n_5649),
.C(n_5399),
.Y(n_8128)
);

A2O1A1Ixp33_ASAP7_75t_L g8129 ( 
.A1(n_7202),
.A2(n_8126),
.B(n_7056),
.C(n_7546),
.Y(n_8129)
);

OAI21xp5_ASAP7_75t_L g8130 ( 
.A1(n_7202),
.A2(n_6438),
.B(n_6194),
.Y(n_8130)
);

NAND2xp5_ASAP7_75t_L g8131 ( 
.A(n_6985),
.B(n_6202),
.Y(n_8131)
);

OAI21x1_ASAP7_75t_L g8132 ( 
.A1(n_7051),
.A2(n_6738),
.B(n_6734),
.Y(n_8132)
);

NAND3xp33_ASAP7_75t_L g8133 ( 
.A(n_7202),
.B(n_6194),
.C(n_5787),
.Y(n_8133)
);

OR2x2_ASAP7_75t_L g8134 ( 
.A(n_7079),
.B(n_6031),
.Y(n_8134)
);

INVx1_ASAP7_75t_L g8135 ( 
.A(n_8087),
.Y(n_8135)
);

OAI21x1_ASAP7_75t_L g8136 ( 
.A1(n_7051),
.A2(n_6738),
.B(n_6734),
.Y(n_8136)
);

NOR2x1_ASAP7_75t_L g8137 ( 
.A(n_6997),
.B(n_6560),
.Y(n_8137)
);

OA21x2_ASAP7_75t_L g8138 ( 
.A1(n_7937),
.A2(n_6915),
.B(n_6909),
.Y(n_8138)
);

INVx1_ASAP7_75t_L g8139 ( 
.A(n_7029),
.Y(n_8139)
);

AO31x2_ASAP7_75t_L g8140 ( 
.A1(n_7095),
.A2(n_6591),
.A3(n_6658),
.B(n_6366),
.Y(n_8140)
);

CKINVDCx5p33_ASAP7_75t_R g8141 ( 
.A(n_6930),
.Y(n_8141)
);

CKINVDCx5p33_ASAP7_75t_R g8142 ( 
.A(n_6930),
.Y(n_8142)
);

OAI21x1_ASAP7_75t_SL g8143 ( 
.A1(n_7095),
.A2(n_5800),
.B(n_6866),
.Y(n_8143)
);

OA21x2_ASAP7_75t_L g8144 ( 
.A1(n_7937),
.A2(n_6915),
.B(n_6909),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_7948),
.Y(n_8145)
);

NAND2xp5_ASAP7_75t_L g8146 ( 
.A(n_6985),
.B(n_6202),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_7029),
.Y(n_8147)
);

NOR2xp33_ASAP7_75t_L g8148 ( 
.A(n_7684),
.B(n_7658),
.Y(n_8148)
);

OAI21x1_ASAP7_75t_L g8149 ( 
.A1(n_7051),
.A2(n_6194),
.B(n_6771),
.Y(n_8149)
);

OA21x2_ASAP7_75t_L g8150 ( 
.A1(n_7937),
.A2(n_6694),
.B(n_6768),
.Y(n_8150)
);

AOI22x1_ASAP7_75t_L g8151 ( 
.A1(n_7079),
.A2(n_6605),
.B1(n_6778),
.B2(n_6596),
.Y(n_8151)
);

INVx2_ASAP7_75t_SL g8152 ( 
.A(n_6997),
.Y(n_8152)
);

OAI22xp5_ASAP7_75t_L g8153 ( 
.A1(n_7251),
.A2(n_5769),
.B1(n_6586),
.B2(n_6526),
.Y(n_8153)
);

INVx1_ASAP7_75t_L g8154 ( 
.A(n_7029),
.Y(n_8154)
);

OAI21x1_ASAP7_75t_L g8155 ( 
.A1(n_7649),
.A2(n_6793),
.B(n_6771),
.Y(n_8155)
);

INVx2_ASAP7_75t_L g8156 ( 
.A(n_7948),
.Y(n_8156)
);

INVx2_ASAP7_75t_L g8157 ( 
.A(n_7948),
.Y(n_8157)
);

INVx3_ASAP7_75t_L g8158 ( 
.A(n_7079),
.Y(n_8158)
);

BUFx12f_ASAP7_75t_L g8159 ( 
.A(n_7946),
.Y(n_8159)
);

BUFx12f_ASAP7_75t_L g8160 ( 
.A(n_7946),
.Y(n_8160)
);

AOI221x1_ASAP7_75t_L g8161 ( 
.A1(n_7251),
.A2(n_7546),
.B1(n_7537),
.B2(n_7684),
.C(n_7391),
.Y(n_8161)
);

A2O1A1Ixp33_ASAP7_75t_L g8162 ( 
.A1(n_8126),
.A2(n_7056),
.B(n_7546),
.C(n_7537),
.Y(n_8162)
);

NAND2xp5_ASAP7_75t_L g8163 ( 
.A(n_6985),
.B(n_6205),
.Y(n_8163)
);

AND2x4_ASAP7_75t_L g8164 ( 
.A(n_7212),
.B(n_6145),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_7327),
.Y(n_8165)
);

OR2x2_ASAP7_75t_L g8166 ( 
.A(n_7115),
.B(n_6997),
.Y(n_8166)
);

OA21x2_ASAP7_75t_L g8167 ( 
.A1(n_7657),
.A2(n_6694),
.B(n_6768),
.Y(n_8167)
);

INVx2_ASAP7_75t_L g8168 ( 
.A(n_7327),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7036),
.Y(n_8169)
);

HB1xp67_ASAP7_75t_L g8170 ( 
.A(n_7038),
.Y(n_8170)
);

CKINVDCx5p33_ASAP7_75t_R g8171 ( 
.A(n_7280),
.Y(n_8171)
);

NAND2x1p5_ASAP7_75t_L g8172 ( 
.A(n_7317),
.B(n_6389),
.Y(n_8172)
);

O2A1O1Ixp33_ASAP7_75t_SL g8173 ( 
.A1(n_7550),
.A2(n_6404),
.B(n_6553),
.C(n_6557),
.Y(n_8173)
);

NAND2xp5_ASAP7_75t_L g8174 ( 
.A(n_7083),
.B(n_6205),
.Y(n_8174)
);

NAND2xp5_ASAP7_75t_SL g8175 ( 
.A(n_7038),
.B(n_6821),
.Y(n_8175)
);

INVx2_ASAP7_75t_SL g8176 ( 
.A(n_7038),
.Y(n_8176)
);

BUFx3_ASAP7_75t_L g8177 ( 
.A(n_7115),
.Y(n_8177)
);

OAI21x1_ASAP7_75t_L g8178 ( 
.A1(n_7649),
.A2(n_6793),
.B(n_6713),
.Y(n_8178)
);

AOI21x1_ASAP7_75t_L g8179 ( 
.A1(n_7649),
.A2(n_6737),
.B(n_6713),
.Y(n_8179)
);

BUFx12f_ASAP7_75t_L g8180 ( 
.A(n_8044),
.Y(n_8180)
);

AOI22xp33_ASAP7_75t_SL g8181 ( 
.A1(n_7537),
.A2(n_6043),
.B1(n_6406),
.B2(n_6515),
.Y(n_8181)
);

OA21x2_ASAP7_75t_L g8182 ( 
.A1(n_7657),
.A2(n_7659),
.B(n_7472),
.Y(n_8182)
);

AO21x2_ASAP7_75t_L g8183 ( 
.A1(n_7657),
.A2(n_6449),
.B(n_6043),
.Y(n_8183)
);

INVx1_ASAP7_75t_L g8184 ( 
.A(n_7036),
.Y(n_8184)
);

OAI21x1_ASAP7_75t_L g8185 ( 
.A1(n_7472),
.A2(n_6789),
.B(n_6872),
.Y(n_8185)
);

INVx2_ASAP7_75t_L g8186 ( 
.A(n_7327),
.Y(n_8186)
);

AO31x2_ASAP7_75t_L g8187 ( 
.A1(n_7095),
.A2(n_6591),
.A3(n_6658),
.B(n_6366),
.Y(n_8187)
);

NAND2xp5_ASAP7_75t_SL g8188 ( 
.A(n_7019),
.B(n_6821),
.Y(n_8188)
);

OAI21x1_ASAP7_75t_L g8189 ( 
.A1(n_7472),
.A2(n_6789),
.B(n_6872),
.Y(n_8189)
);

OAI21xp5_ASAP7_75t_L g8190 ( 
.A1(n_7251),
.A2(n_5790),
.B(n_5914),
.Y(n_8190)
);

BUFx3_ASAP7_75t_L g8191 ( 
.A(n_7115),
.Y(n_8191)
);

AOI22xp33_ASAP7_75t_L g8192 ( 
.A1(n_7397),
.A2(n_6043),
.B1(n_6482),
.B2(n_6505),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7036),
.Y(n_8193)
);

NOR2xp33_ASAP7_75t_L g8194 ( 
.A(n_7684),
.B(n_5908),
.Y(n_8194)
);

AOI21xp5_ASAP7_75t_L g8195 ( 
.A1(n_7624),
.A2(n_7744),
.B(n_7715),
.Y(n_8195)
);

OAI21xp5_ASAP7_75t_L g8196 ( 
.A1(n_7056),
.A2(n_5790),
.B(n_5914),
.Y(n_8196)
);

NAND2x1p5_ASAP7_75t_L g8197 ( 
.A(n_7317),
.B(n_6389),
.Y(n_8197)
);

AOI22xp33_ASAP7_75t_L g8198 ( 
.A1(n_7397),
.A2(n_6043),
.B1(n_6482),
.B2(n_6505),
.Y(n_8198)
);

AOI21xp5_ASAP7_75t_L g8199 ( 
.A1(n_7624),
.A2(n_6896),
.B(n_6894),
.Y(n_8199)
);

CKINVDCx8_ASAP7_75t_R g8200 ( 
.A(n_6928),
.Y(n_8200)
);

INVx1_ASAP7_75t_L g8201 ( 
.A(n_7046),
.Y(n_8201)
);

OR2x6_ASAP7_75t_L g8202 ( 
.A(n_8110),
.B(n_6640),
.Y(n_8202)
);

AND2x4_ASAP7_75t_L g8203 ( 
.A(n_7212),
.B(n_6145),
.Y(n_8203)
);

INVx2_ASAP7_75t_SL g8204 ( 
.A(n_7212),
.Y(n_8204)
);

INVx2_ASAP7_75t_L g8205 ( 
.A(n_7327),
.Y(n_8205)
);

OR2x6_ASAP7_75t_L g8206 ( 
.A(n_8110),
.B(n_6640),
.Y(n_8206)
);

OAI21xp5_ASAP7_75t_L g8207 ( 
.A1(n_7658),
.A2(n_5914),
.B(n_5843),
.Y(n_8207)
);

OAI21x1_ASAP7_75t_L g8208 ( 
.A1(n_7472),
.A2(n_6789),
.B(n_6872),
.Y(n_8208)
);

BUFx2_ASAP7_75t_L g8209 ( 
.A(n_7930),
.Y(n_8209)
);

OAI21x1_ASAP7_75t_L g8210 ( 
.A1(n_7647),
.A2(n_7744),
.B(n_7748),
.Y(n_8210)
);

BUFx6f_ASAP7_75t_L g8211 ( 
.A(n_6926),
.Y(n_8211)
);

OAI21x1_ASAP7_75t_L g8212 ( 
.A1(n_7647),
.A2(n_6663),
.B(n_6701),
.Y(n_8212)
);

AND2x2_ASAP7_75t_L g8213 ( 
.A(n_8081),
.B(n_6455),
.Y(n_8213)
);

AO21x2_ASAP7_75t_L g8214 ( 
.A1(n_7744),
.A2(n_6449),
.B(n_6732),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_8087),
.Y(n_8215)
);

AND2x4_ASAP7_75t_L g8216 ( 
.A(n_7212),
.B(n_6145),
.Y(n_8216)
);

BUFx2_ASAP7_75t_L g8217 ( 
.A(n_7930),
.Y(n_8217)
);

AO31x2_ASAP7_75t_L g8218 ( 
.A1(n_7095),
.A2(n_6526),
.A3(n_6528),
.B(n_6515),
.Y(n_8218)
);

OAI21x1_ASAP7_75t_L g8219 ( 
.A1(n_7647),
.A2(n_7748),
.B(n_7128),
.Y(n_8219)
);

OAI21x1_ASAP7_75t_L g8220 ( 
.A1(n_7748),
.A2(n_6663),
.B(n_6701),
.Y(n_8220)
);

HB1xp67_ASAP7_75t_L g8221 ( 
.A(n_7419),
.Y(n_8221)
);

AOI22xp33_ASAP7_75t_L g8222 ( 
.A1(n_7345),
.A2(n_6183),
.B1(n_5770),
.B2(n_5787),
.Y(n_8222)
);

INVxp67_ASAP7_75t_L g8223 ( 
.A(n_7615),
.Y(n_8223)
);

OAI21x1_ASAP7_75t_L g8224 ( 
.A1(n_7128),
.A2(n_7659),
.B(n_7958),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_8087),
.Y(n_8225)
);

AO21x2_ASAP7_75t_L g8226 ( 
.A1(n_7659),
.A2(n_6732),
.B(n_6834),
.Y(n_8226)
);

INVx2_ASAP7_75t_L g8227 ( 
.A(n_7339),
.Y(n_8227)
);

INVx1_ASAP7_75t_L g8228 ( 
.A(n_8088),
.Y(n_8228)
);

NAND3xp33_ASAP7_75t_L g8229 ( 
.A(n_7391),
.B(n_5770),
.C(n_5769),
.Y(n_8229)
);

NAND2xp5_ASAP7_75t_L g8230 ( 
.A(n_7083),
.B(n_6031),
.Y(n_8230)
);

OAI221xp5_ASAP7_75t_L g8231 ( 
.A1(n_7735),
.A2(n_6509),
.B1(n_5843),
.B2(n_5751),
.C(n_6582),
.Y(n_8231)
);

INVx5_ASAP7_75t_L g8232 ( 
.A(n_7819),
.Y(n_8232)
);

OAI21xp5_ASAP7_75t_L g8233 ( 
.A1(n_7528),
.A2(n_7391),
.B(n_7735),
.Y(n_8233)
);

INVx2_ASAP7_75t_L g8234 ( 
.A(n_7339),
.Y(n_8234)
);

INVx1_ASAP7_75t_L g8235 ( 
.A(n_7046),
.Y(n_8235)
);

HB1xp67_ASAP7_75t_L g8236 ( 
.A(n_7419),
.Y(n_8236)
);

OAI21x1_ASAP7_75t_L g8237 ( 
.A1(n_7128),
.A2(n_6707),
.B(n_6544),
.Y(n_8237)
);

AND2x4_ASAP7_75t_L g8238 ( 
.A(n_7212),
.B(n_6145),
.Y(n_8238)
);

INVx2_ASAP7_75t_SL g8239 ( 
.A(n_7212),
.Y(n_8239)
);

INVx1_ASAP7_75t_SL g8240 ( 
.A(n_7652),
.Y(n_8240)
);

OAI22xp5_ASAP7_75t_L g8241 ( 
.A1(n_6975),
.A2(n_6586),
.B1(n_6528),
.B2(n_6509),
.Y(n_8241)
);

NAND2xp5_ASAP7_75t_SL g8242 ( 
.A(n_7019),
.B(n_6831),
.Y(n_8242)
);

OAI21x1_ASAP7_75t_L g8243 ( 
.A1(n_7958),
.A2(n_7994),
.B(n_7961),
.Y(n_8243)
);

INVx2_ASAP7_75t_L g8244 ( 
.A(n_7339),
.Y(n_8244)
);

OA21x2_ASAP7_75t_L g8245 ( 
.A1(n_7853),
.A2(n_6442),
.B(n_6896),
.Y(n_8245)
);

BUFx3_ASAP7_75t_L g8246 ( 
.A(n_7458),
.Y(n_8246)
);

INVx2_ASAP7_75t_L g8247 ( 
.A(n_7339),
.Y(n_8247)
);

INVx1_ASAP7_75t_L g8248 ( 
.A(n_7046),
.Y(n_8248)
);

OAI21x1_ASAP7_75t_L g8249 ( 
.A1(n_7958),
.A2(n_6707),
.B(n_6544),
.Y(n_8249)
);

OAI21x1_ASAP7_75t_L g8250 ( 
.A1(n_7961),
.A2(n_6689),
.B(n_6680),
.Y(n_8250)
);

AOI21xp5_ASAP7_75t_L g8251 ( 
.A1(n_7715),
.A2(n_6894),
.B(n_6582),
.Y(n_8251)
);

OAI21x1_ASAP7_75t_L g8252 ( 
.A1(n_7961),
.A2(n_6689),
.B(n_6680),
.Y(n_8252)
);

INVx1_ASAP7_75t_L g8253 ( 
.A(n_7059),
.Y(n_8253)
);

OAI21x1_ASAP7_75t_L g8254 ( 
.A1(n_7994),
.A2(n_6497),
.B(n_6480),
.Y(n_8254)
);

OAI21x1_ASAP7_75t_L g8255 ( 
.A1(n_7994),
.A2(n_6497),
.B(n_6480),
.Y(n_8255)
);

AND2x4_ASAP7_75t_L g8256 ( 
.A(n_7212),
.B(n_6190),
.Y(n_8256)
);

CKINVDCx16_ASAP7_75t_R g8257 ( 
.A(n_7022),
.Y(n_8257)
);

OAI21x1_ASAP7_75t_L g8258 ( 
.A1(n_7853),
.A2(n_6536),
.B(n_6527),
.Y(n_8258)
);

BUFx3_ASAP7_75t_L g8259 ( 
.A(n_7458),
.Y(n_8259)
);

OAI21x1_ASAP7_75t_SL g8260 ( 
.A1(n_7087),
.A2(n_5800),
.B(n_6878),
.Y(n_8260)
);

INVx1_ASAP7_75t_L g8261 ( 
.A(n_7059),
.Y(n_8261)
);

NOR2xp67_ASAP7_75t_L g8262 ( 
.A(n_7977),
.B(n_5761),
.Y(n_8262)
);

BUFx2_ASAP7_75t_L g8263 ( 
.A(n_7930),
.Y(n_8263)
);

OAI21x1_ASAP7_75t_L g8264 ( 
.A1(n_7853),
.A2(n_6536),
.B(n_6527),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_7059),
.Y(n_8265)
);

OAI21x1_ASAP7_75t_L g8266 ( 
.A1(n_7020),
.A2(n_7035),
.B(n_7033),
.Y(n_8266)
);

NOR2xp33_ASAP7_75t_L g8267 ( 
.A(n_7083),
.B(n_7880),
.Y(n_8267)
);

OAI22xp5_ASAP7_75t_L g8268 ( 
.A1(n_6975),
.A2(n_5854),
.B1(n_5888),
.B2(n_5789),
.Y(n_8268)
);

CKINVDCx5p33_ASAP7_75t_R g8269 ( 
.A(n_7280),
.Y(n_8269)
);

OAI21x1_ASAP7_75t_L g8270 ( 
.A1(n_7020),
.A2(n_5738),
.B(n_6712),
.Y(n_8270)
);

AOI22xp33_ASAP7_75t_L g8271 ( 
.A1(n_7345),
.A2(n_6183),
.B1(n_5924),
.B2(n_5833),
.Y(n_8271)
);

INVx1_ASAP7_75t_SL g8272 ( 
.A(n_7652),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_7077),
.Y(n_8273)
);

OAI21x1_ASAP7_75t_L g8274 ( 
.A1(n_7020),
.A2(n_5738),
.B(n_6712),
.Y(n_8274)
);

A2O1A1Ixp33_ASAP7_75t_L g8275 ( 
.A1(n_7735),
.A2(n_5751),
.B(n_6647),
.C(n_5745),
.Y(n_8275)
);

OA21x2_ASAP7_75t_L g8276 ( 
.A1(n_7465),
.A2(n_6442),
.B(n_6647),
.Y(n_8276)
);

OAI21x1_ASAP7_75t_L g8277 ( 
.A1(n_7033),
.A2(n_5738),
.B(n_6594),
.Y(n_8277)
);

AOI21xp5_ASAP7_75t_L g8278 ( 
.A1(n_7715),
.A2(n_6864),
.B(n_6692),
.Y(n_8278)
);

INVx2_ASAP7_75t_L g8279 ( 
.A(n_7364),
.Y(n_8279)
);

INVxp67_ASAP7_75t_L g8280 ( 
.A(n_7615),
.Y(n_8280)
);

OAI21x1_ASAP7_75t_L g8281 ( 
.A1(n_7033),
.A2(n_6594),
.B(n_6702),
.Y(n_8281)
);

OAI21x1_ASAP7_75t_L g8282 ( 
.A1(n_7035),
.A2(n_6702),
.B(n_6487),
.Y(n_8282)
);

INVx1_ASAP7_75t_L g8283 ( 
.A(n_7077),
.Y(n_8283)
);

AOI22xp33_ASAP7_75t_SL g8284 ( 
.A1(n_8055),
.A2(n_6406),
.B1(n_6423),
.B2(n_5892),
.Y(n_8284)
);

NAND3xp33_ASAP7_75t_L g8285 ( 
.A(n_7550),
.B(n_7569),
.C(n_7495),
.Y(n_8285)
);

AOI22xp5_ASAP7_75t_L g8286 ( 
.A1(n_7345),
.A2(n_5888),
.B1(n_5912),
.B2(n_5776),
.Y(n_8286)
);

NAND3xp33_ASAP7_75t_L g8287 ( 
.A(n_7495),
.B(n_6560),
.C(n_6520),
.Y(n_8287)
);

AND2x2_ASAP7_75t_L g8288 ( 
.A(n_8081),
.B(n_7254),
.Y(n_8288)
);

INVx2_ASAP7_75t_L g8289 ( 
.A(n_7364),
.Y(n_8289)
);

OAI22xp33_ASAP7_75t_L g8290 ( 
.A1(n_7292),
.A2(n_6618),
.B1(n_6248),
.B2(n_6667),
.Y(n_8290)
);

OA21x2_ASAP7_75t_L g8291 ( 
.A1(n_7465),
.A2(n_6882),
.B(n_6825),
.Y(n_8291)
);

HB1xp67_ASAP7_75t_L g8292 ( 
.A(n_7429),
.Y(n_8292)
);

INVx1_ASAP7_75t_L g8293 ( 
.A(n_8088),
.Y(n_8293)
);

NAND2xp5_ASAP7_75t_L g8294 ( 
.A(n_7031),
.B(n_6050),
.Y(n_8294)
);

AO21x2_ASAP7_75t_L g8295 ( 
.A1(n_7110),
.A2(n_6834),
.B(n_6737),
.Y(n_8295)
);

INVx3_ASAP7_75t_L g8296 ( 
.A(n_7039),
.Y(n_8296)
);

OA21x2_ASAP7_75t_L g8297 ( 
.A1(n_7465),
.A2(n_7614),
.B(n_7479),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_7077),
.Y(n_8298)
);

INVxp67_ASAP7_75t_L g8299 ( 
.A(n_7615),
.Y(n_8299)
);

INVx2_ASAP7_75t_L g8300 ( 
.A(n_7364),
.Y(n_8300)
);

NAND2xp5_ASAP7_75t_L g8301 ( 
.A(n_7031),
.B(n_6050),
.Y(n_8301)
);

AOI22x1_ASAP7_75t_L g8302 ( 
.A1(n_7569),
.A2(n_6778),
.B1(n_6876),
.B2(n_6605),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7086),
.Y(n_8303)
);

AOI22xp5_ASAP7_75t_L g8304 ( 
.A1(n_7292),
.A2(n_7331),
.B1(n_8055),
.B2(n_7395),
.Y(n_8304)
);

OAI21x1_ASAP7_75t_L g8305 ( 
.A1(n_7035),
.A2(n_6487),
.B(n_6847),
.Y(n_8305)
);

INVx3_ASAP7_75t_L g8306 ( 
.A(n_7039),
.Y(n_8306)
);

OAI21xp5_ASAP7_75t_L g8307 ( 
.A1(n_7528),
.A2(n_6520),
.B(n_5789),
.Y(n_8307)
);

INVx1_ASAP7_75t_SL g8308 ( 
.A(n_7644),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_8081),
.B(n_6430),
.Y(n_8309)
);

BUFx2_ASAP7_75t_L g8310 ( 
.A(n_7930),
.Y(n_8310)
);

NAND2xp5_ASAP7_75t_L g8311 ( 
.A(n_7031),
.B(n_6056),
.Y(n_8311)
);

AND2x2_ASAP7_75t_L g8312 ( 
.A(n_8081),
.B(n_6430),
.Y(n_8312)
);

INVxp67_ASAP7_75t_L g8313 ( 
.A(n_7459),
.Y(n_8313)
);

NAND2xp5_ASAP7_75t_L g8314 ( 
.A(n_7122),
.B(n_6056),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_8088),
.Y(n_8315)
);

O2A1O1Ixp33_ASAP7_75t_L g8316 ( 
.A1(n_7260),
.A2(n_5924),
.B(n_5941),
.C(n_5908),
.Y(n_8316)
);

AND2x4_ASAP7_75t_L g8317 ( 
.A(n_7039),
.B(n_6190),
.Y(n_8317)
);

NOR2xp67_ASAP7_75t_L g8318 ( 
.A(n_7977),
.B(n_5761),
.Y(n_8318)
);

NOR2xp67_ASAP7_75t_L g8319 ( 
.A(n_7977),
.B(n_7134),
.Y(n_8319)
);

OAI21x1_ASAP7_75t_L g8320 ( 
.A1(n_7057),
.A2(n_6847),
.B(n_6788),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_8111),
.Y(n_8321)
);

AO21x2_ASAP7_75t_L g8322 ( 
.A1(n_7110),
.A2(n_6183),
.B(n_6593),
.Y(n_8322)
);

OAI21x1_ASAP7_75t_L g8323 ( 
.A1(n_7057),
.A2(n_6788),
.B(n_6757),
.Y(n_8323)
);

OAI22xp5_ASAP7_75t_L g8324 ( 
.A1(n_6975),
.A2(n_5854),
.B1(n_5776),
.B2(n_5807),
.Y(n_8324)
);

AO21x1_ASAP7_75t_L g8325 ( 
.A1(n_7050),
.A2(n_6674),
.B(n_6452),
.Y(n_8325)
);

INVx2_ASAP7_75t_SL g8326 ( 
.A(n_7039),
.Y(n_8326)
);

O2A1O1Ixp33_ASAP7_75t_L g8327 ( 
.A1(n_7260),
.A2(n_5924),
.B(n_5941),
.C(n_5745),
.Y(n_8327)
);

INVx2_ASAP7_75t_L g8328 ( 
.A(n_7364),
.Y(n_8328)
);

AOI21xp5_ASAP7_75t_L g8329 ( 
.A1(n_8055),
.A2(n_6864),
.B(n_6621),
.Y(n_8329)
);

NAND2x1p5_ASAP7_75t_L g8330 ( 
.A(n_7317),
.B(n_6389),
.Y(n_8330)
);

NOR2xp67_ASAP7_75t_L g8331 ( 
.A(n_7134),
.B(n_5761),
.Y(n_8331)
);

OAI21x1_ASAP7_75t_L g8332 ( 
.A1(n_7057),
.A2(n_6819),
.B(n_6757),
.Y(n_8332)
);

OAI21x1_ASAP7_75t_L g8333 ( 
.A1(n_7448),
.A2(n_6819),
.B(n_6845),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_7086),
.Y(n_8334)
);

AOI21xp5_ASAP7_75t_L g8335 ( 
.A1(n_8055),
.A2(n_6920),
.B(n_6621),
.Y(n_8335)
);

OR2x6_ASAP7_75t_L g8336 ( 
.A(n_8110),
.B(n_6270),
.Y(n_8336)
);

AOI22xp33_ASAP7_75t_L g8337 ( 
.A1(n_7331),
.A2(n_6183),
.B1(n_5833),
.B2(n_6130),
.Y(n_8337)
);

BUFx2_ASAP7_75t_R g8338 ( 
.A(n_7816),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_7086),
.Y(n_8339)
);

NOR2xp33_ASAP7_75t_L g8340 ( 
.A(n_7880),
.B(n_5832),
.Y(n_8340)
);

INVx2_ASAP7_75t_L g8341 ( 
.A(n_7101),
.Y(n_8341)
);

INVx2_ASAP7_75t_L g8342 ( 
.A(n_7101),
.Y(n_8342)
);

INVx1_ASAP7_75t_L g8343 ( 
.A(n_7088),
.Y(n_8343)
);

INVx2_ASAP7_75t_L g8344 ( 
.A(n_7101),
.Y(n_8344)
);

INVx2_ASAP7_75t_SL g8345 ( 
.A(n_7039),
.Y(n_8345)
);

BUFx3_ASAP7_75t_L g8346 ( 
.A(n_7458),
.Y(n_8346)
);

INVx2_ASAP7_75t_L g8347 ( 
.A(n_7101),
.Y(n_8347)
);

OAI22xp33_ASAP7_75t_L g8348 ( 
.A1(n_7292),
.A2(n_6618),
.B1(n_6248),
.B2(n_6667),
.Y(n_8348)
);

NOR2xp33_ASAP7_75t_L g8349 ( 
.A(n_7349),
.B(n_6612),
.Y(n_8349)
);

OR3x4_ASAP7_75t_SL g8350 ( 
.A(n_7260),
.B(n_6708),
.C(n_6612),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_7088),
.Y(n_8351)
);

INVx2_ASAP7_75t_L g8352 ( 
.A(n_7102),
.Y(n_8352)
);

AO31x2_ASAP7_75t_L g8353 ( 
.A1(n_7851),
.A2(n_6603),
.A3(n_5930),
.B(n_6783),
.Y(n_8353)
);

OA21x2_ASAP7_75t_L g8354 ( 
.A1(n_7479),
.A2(n_6882),
.B(n_6825),
.Y(n_8354)
);

OAI22xp5_ASAP7_75t_L g8355 ( 
.A1(n_6975),
.A2(n_5785),
.B1(n_5810),
.B2(n_6570),
.Y(n_8355)
);

AOI22xp33_ASAP7_75t_L g8356 ( 
.A1(n_7331),
.A2(n_6183),
.B1(n_5993),
.B2(n_6130),
.Y(n_8356)
);

NAND2x1p5_ASAP7_75t_L g8357 ( 
.A(n_7317),
.B(n_6389),
.Y(n_8357)
);

AOI21x1_ASAP7_75t_L g8358 ( 
.A1(n_7572),
.A2(n_7676),
.B(n_7400),
.Y(n_8358)
);

HB1xp67_ASAP7_75t_L g8359 ( 
.A(n_7429),
.Y(n_8359)
);

BUFx6f_ASAP7_75t_L g8360 ( 
.A(n_6926),
.Y(n_8360)
);

CKINVDCx5p33_ASAP7_75t_R g8361 ( 
.A(n_7433),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_8111),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_8111),
.Y(n_8363)
);

AO31x2_ASAP7_75t_L g8364 ( 
.A1(n_7851),
.A2(n_6603),
.A3(n_5930),
.B(n_6783),
.Y(n_8364)
);

OR2x6_ASAP7_75t_L g8365 ( 
.A(n_8110),
.B(n_6270),
.Y(n_8365)
);

BUFx3_ASAP7_75t_L g8366 ( 
.A(n_7458),
.Y(n_8366)
);

INVx2_ASAP7_75t_L g8367 ( 
.A(n_7102),
.Y(n_8367)
);

OAI21x1_ASAP7_75t_L g8368 ( 
.A1(n_7448),
.A2(n_6845),
.B(n_5792),
.Y(n_8368)
);

OAI21x1_ASAP7_75t_L g8369 ( 
.A1(n_7448),
.A2(n_5792),
.B(n_5739),
.Y(n_8369)
);

AOI221xp5_ASAP7_75t_L g8370 ( 
.A1(n_8005),
.A2(n_6593),
.B1(n_6452),
.B2(n_6427),
.C(n_5993),
.Y(n_8370)
);

OAI21x1_ASAP7_75t_L g8371 ( 
.A1(n_7448),
.A2(n_6996),
.B(n_7110),
.Y(n_8371)
);

NOR2x1_ASAP7_75t_SL g8372 ( 
.A(n_7012),
.B(n_5976),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7088),
.Y(n_8373)
);

NOR2xp67_ASAP7_75t_L g8374 ( 
.A(n_7134),
.B(n_6105),
.Y(n_8374)
);

INVx1_ASAP7_75t_L g8375 ( 
.A(n_7096),
.Y(n_8375)
);

OR2x2_ASAP7_75t_L g8376 ( 
.A(n_7019),
.B(n_6076),
.Y(n_8376)
);

INVx3_ASAP7_75t_L g8377 ( 
.A(n_7039),
.Y(n_8377)
);

BUFx3_ASAP7_75t_L g8378 ( 
.A(n_7954),
.Y(n_8378)
);

INVx1_ASAP7_75t_L g8379 ( 
.A(n_7096),
.Y(n_8379)
);

INVx2_ASAP7_75t_L g8380 ( 
.A(n_7102),
.Y(n_8380)
);

AND2x4_ASAP7_75t_L g8381 ( 
.A(n_7039),
.B(n_6190),
.Y(n_8381)
);

INVx2_ASAP7_75t_SL g8382 ( 
.A(n_7081),
.Y(n_8382)
);

OR2x6_ASAP7_75t_L g8383 ( 
.A(n_8110),
.B(n_6270),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_7096),
.Y(n_8384)
);

AND2x4_ASAP7_75t_L g8385 ( 
.A(n_7081),
.B(n_6190),
.Y(n_8385)
);

HB1xp67_ASAP7_75t_L g8386 ( 
.A(n_7434),
.Y(n_8386)
);

AOI21x1_ASAP7_75t_L g8387 ( 
.A1(n_7572),
.A2(n_6419),
.B(n_5889),
.Y(n_8387)
);

OAI21x1_ASAP7_75t_L g8388 ( 
.A1(n_7107),
.A2(n_5804),
.B(n_5880),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7105),
.Y(n_8389)
);

OAI21x1_ASAP7_75t_L g8390 ( 
.A1(n_7107),
.A2(n_5804),
.B(n_5880),
.Y(n_8390)
);

AO21x2_ASAP7_75t_L g8391 ( 
.A1(n_7107),
.A2(n_6899),
.B(n_6550),
.Y(n_8391)
);

OAI21xp5_ASAP7_75t_L g8392 ( 
.A1(n_7528),
.A2(n_5889),
.B(n_6660),
.Y(n_8392)
);

AO21x2_ASAP7_75t_L g8393 ( 
.A1(n_7146),
.A2(n_6899),
.B(n_6550),
.Y(n_8393)
);

AND2x4_ASAP7_75t_L g8394 ( 
.A(n_7081),
.B(n_6190),
.Y(n_8394)
);

AOI22xp33_ASAP7_75t_L g8395 ( 
.A1(n_7331),
.A2(n_5778),
.B1(n_5944),
.B2(n_5912),
.Y(n_8395)
);

OAI21x1_ASAP7_75t_L g8396 ( 
.A1(n_7791),
.A2(n_7163),
.B(n_6991),
.Y(n_8396)
);

AOI21x1_ASAP7_75t_L g8397 ( 
.A1(n_7572),
.A2(n_6419),
.B(n_6813),
.Y(n_8397)
);

INVx1_ASAP7_75t_L g8398 ( 
.A(n_7105),
.Y(n_8398)
);

AOI22xp33_ASAP7_75t_L g8399 ( 
.A1(n_7331),
.A2(n_5778),
.B1(n_5944),
.B2(n_6057),
.Y(n_8399)
);

AOI21xp5_ASAP7_75t_L g8400 ( 
.A1(n_8055),
.A2(n_6920),
.B(n_6814),
.Y(n_8400)
);

INVx5_ASAP7_75t_L g8401 ( 
.A(n_7819),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_7102),
.Y(n_8402)
);

AND2x4_ASAP7_75t_L g8403 ( 
.A(n_7081),
.B(n_6193),
.Y(n_8403)
);

BUFx2_ASAP7_75t_L g8404 ( 
.A(n_7930),
.Y(n_8404)
);

OAI21x1_ASAP7_75t_L g8405 ( 
.A1(n_7791),
.A2(n_6814),
.B(n_6813),
.Y(n_8405)
);

OAI22xp33_ASAP7_75t_L g8406 ( 
.A1(n_7790),
.A2(n_8113),
.B1(n_7782),
.B2(n_7796),
.Y(n_8406)
);

INVx1_ASAP7_75t_SL g8407 ( 
.A(n_7644),
.Y(n_8407)
);

AOI21xp5_ASAP7_75t_SL g8408 ( 
.A1(n_7905),
.A2(n_5892),
.B(n_5902),
.Y(n_8408)
);

INVx2_ASAP7_75t_L g8409 ( 
.A(n_7112),
.Y(n_8409)
);

NOR2xp33_ASAP7_75t_L g8410 ( 
.A(n_7349),
.B(n_5874),
.Y(n_8410)
);

OAI21x1_ASAP7_75t_L g8411 ( 
.A1(n_7791),
.A2(n_5855),
.B(n_6604),
.Y(n_8411)
);

CKINVDCx5p33_ASAP7_75t_R g8412 ( 
.A(n_7433),
.Y(n_8412)
);

AOI22xp33_ASAP7_75t_L g8413 ( 
.A1(n_7331),
.A2(n_6057),
.B1(n_6126),
.B2(n_5785),
.Y(n_8413)
);

INVx2_ASAP7_75t_L g8414 ( 
.A(n_7112),
.Y(n_8414)
);

AOI22xp5_ASAP7_75t_L g8415 ( 
.A1(n_8055),
.A2(n_5845),
.B1(n_5758),
.B2(n_5848),
.Y(n_8415)
);

OAI22xp5_ASAP7_75t_L g8416 ( 
.A1(n_7781),
.A2(n_5902),
.B1(n_5911),
.B2(n_5824),
.Y(n_8416)
);

NAND2xp5_ASAP7_75t_L g8417 ( 
.A(n_7122),
.B(n_6076),
.Y(n_8417)
);

AOI22xp33_ASAP7_75t_L g8418 ( 
.A1(n_8055),
.A2(n_6126),
.B1(n_5734),
.B2(n_6215),
.Y(n_8418)
);

AO31x2_ASAP7_75t_L g8419 ( 
.A1(n_7851),
.A2(n_6604),
.A3(n_6831),
.B(n_6606),
.Y(n_8419)
);

INVx2_ASAP7_75t_L g8420 ( 
.A(n_7112),
.Y(n_8420)
);

INVx2_ASAP7_75t_L g8421 ( 
.A(n_7112),
.Y(n_8421)
);

A2O1A1Ixp33_ASAP7_75t_L g8422 ( 
.A1(n_7227),
.A2(n_5734),
.B(n_5884),
.C(n_6387),
.Y(n_8422)
);

OAI22xp5_ASAP7_75t_L g8423 ( 
.A1(n_7781),
.A2(n_5911),
.B1(n_5824),
.B2(n_5850),
.Y(n_8423)
);

AOI221xp5_ASAP7_75t_L g8424 ( 
.A1(n_8005),
.A2(n_6624),
.B1(n_6683),
.B2(n_6643),
.C(n_6642),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_7125),
.Y(n_8425)
);

OA21x2_ASAP7_75t_L g8426 ( 
.A1(n_7479),
.A2(n_6320),
.B(n_6311),
.Y(n_8426)
);

INVx2_ASAP7_75t_SL g8427 ( 
.A(n_7081),
.Y(n_8427)
);

NAND2x1p5_ASAP7_75t_L g8428 ( 
.A(n_7317),
.B(n_6416),
.Y(n_8428)
);

OAI21x1_ASAP7_75t_L g8429 ( 
.A1(n_7163),
.A2(n_5855),
.B(n_5875),
.Y(n_8429)
);

NAND2xp5_ASAP7_75t_L g8430 ( 
.A(n_7122),
.B(n_6079),
.Y(n_8430)
);

O2A1O1Ixp33_ASAP7_75t_L g8431 ( 
.A1(n_7260),
.A2(n_5884),
.B(n_6666),
.C(n_6660),
.Y(n_8431)
);

OAI21x1_ASAP7_75t_L g8432 ( 
.A1(n_7163),
.A2(n_5877),
.B(n_5875),
.Y(n_8432)
);

INVx2_ASAP7_75t_L g8433 ( 
.A(n_7125),
.Y(n_8433)
);

NAND2xp5_ASAP7_75t_L g8434 ( 
.A(n_7140),
.B(n_6079),
.Y(n_8434)
);

AND2x4_ASAP7_75t_L g8435 ( 
.A(n_7081),
.B(n_6193),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7105),
.Y(n_8436)
);

O2A1O1Ixp33_ASAP7_75t_SL g8437 ( 
.A1(n_7179),
.A2(n_6553),
.B(n_6557),
.C(n_5870),
.Y(n_8437)
);

HB1xp67_ASAP7_75t_L g8438 ( 
.A(n_7434),
.Y(n_8438)
);

NOR2xp33_ASAP7_75t_L g8439 ( 
.A(n_7882),
.B(n_5874),
.Y(n_8439)
);

INVx2_ASAP7_75t_L g8440 ( 
.A(n_7125),
.Y(n_8440)
);

BUFx10_ASAP7_75t_L g8441 ( 
.A(n_7485),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_7114),
.Y(n_8442)
);

CKINVDCx8_ASAP7_75t_R g8443 ( 
.A(n_6928),
.Y(n_8443)
);

OAI21x1_ASAP7_75t_L g8444 ( 
.A1(n_6991),
.A2(n_5877),
.B(n_6606),
.Y(n_8444)
);

OA21x2_ASAP7_75t_L g8445 ( 
.A1(n_7614),
.A2(n_6320),
.B(n_6311),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_7114),
.Y(n_8446)
);

OAI21xp5_ASAP7_75t_L g8447 ( 
.A1(n_7790),
.A2(n_6666),
.B(n_5871),
.Y(n_8447)
);

OAI22xp5_ASAP7_75t_L g8448 ( 
.A1(n_7782),
.A2(n_5850),
.B1(n_6669),
.B2(n_6648),
.Y(n_8448)
);

OAI21x1_ASAP7_75t_L g8449 ( 
.A1(n_6991),
.A2(n_6859),
.B(n_5940),
.Y(n_8449)
);

AND2x4_ASAP7_75t_L g8450 ( 
.A(n_7081),
.B(n_6193),
.Y(n_8450)
);

AOI21xp33_ASAP7_75t_L g8451 ( 
.A1(n_7827),
.A2(n_6919),
.B(n_6889),
.Y(n_8451)
);

CKINVDCx20_ASAP7_75t_R g8452 ( 
.A(n_7421),
.Y(n_8452)
);

OAI21x1_ASAP7_75t_L g8453 ( 
.A1(n_8008),
.A2(n_6859),
.B(n_5940),
.Y(n_8453)
);

AOI21xp5_ASAP7_75t_L g8454 ( 
.A1(n_7851),
.A2(n_6322),
.B(n_6843),
.Y(n_8454)
);

BUFx3_ASAP7_75t_L g8455 ( 
.A(n_7954),
.Y(n_8455)
);

OAI21x1_ASAP7_75t_L g8456 ( 
.A1(n_8008),
.A2(n_5936),
.B(n_6613),
.Y(n_8456)
);

INVx2_ASAP7_75t_L g8457 ( 
.A(n_7125),
.Y(n_8457)
);

INVx2_ASAP7_75t_L g8458 ( 
.A(n_7130),
.Y(n_8458)
);

INVx2_ASAP7_75t_L g8459 ( 
.A(n_7130),
.Y(n_8459)
);

AOI21x1_ASAP7_75t_L g8460 ( 
.A1(n_7676),
.A2(n_6918),
.B(n_6912),
.Y(n_8460)
);

OAI21x1_ASAP7_75t_L g8461 ( 
.A1(n_8008),
.A2(n_8010),
.B(n_7922),
.Y(n_8461)
);

AO32x2_ASAP7_75t_L g8462 ( 
.A1(n_8005),
.A2(n_6643),
.A3(n_6683),
.B1(n_6642),
.B2(n_6624),
.Y(n_8462)
);

OAI21x1_ASAP7_75t_L g8463 ( 
.A1(n_8010),
.A2(n_5936),
.B(n_6613),
.Y(n_8463)
);

OAI21x1_ASAP7_75t_L g8464 ( 
.A1(n_8010),
.A2(n_6843),
.B(n_6041),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7114),
.Y(n_8465)
);

NAND2xp5_ASAP7_75t_L g8466 ( 
.A(n_7140),
.B(n_6094),
.Y(n_8466)
);

O2A1O1Ixp33_ASAP7_75t_L g8467 ( 
.A1(n_7260),
.A2(n_5870),
.B(n_5860),
.C(n_5898),
.Y(n_8467)
);

OR2x2_ASAP7_75t_L g8468 ( 
.A(n_8024),
.B(n_6094),
.Y(n_8468)
);

AND2x4_ASAP7_75t_L g8469 ( 
.A(n_7224),
.B(n_6193),
.Y(n_8469)
);

AOI22xp33_ASAP7_75t_L g8470 ( 
.A1(n_7490),
.A2(n_6215),
.B1(n_5955),
.B2(n_6513),
.Y(n_8470)
);

OA21x2_ASAP7_75t_L g8471 ( 
.A1(n_7614),
.A2(n_6685),
.B(n_6524),
.Y(n_8471)
);

OAI21x1_ASAP7_75t_L g8472 ( 
.A1(n_7870),
.A2(n_6041),
.B(n_6006),
.Y(n_8472)
);

OAI21xp5_ASAP7_75t_L g8473 ( 
.A1(n_7790),
.A2(n_5871),
.B(n_6456),
.Y(n_8473)
);

OA21x2_ASAP7_75t_L g8474 ( 
.A1(n_7947),
.A2(n_6685),
.B(n_6524),
.Y(n_8474)
);

NOR2xp33_ASAP7_75t_L g8475 ( 
.A(n_7882),
.B(n_7140),
.Y(n_8475)
);

OAI21xp5_ASAP7_75t_L g8476 ( 
.A1(n_7227),
.A2(n_6457),
.B(n_6456),
.Y(n_8476)
);

INVx1_ASAP7_75t_L g8477 ( 
.A(n_7120),
.Y(n_8477)
);

OAI21x1_ASAP7_75t_L g8478 ( 
.A1(n_7870),
.A2(n_6041),
.B(n_6006),
.Y(n_8478)
);

AO31x2_ASAP7_75t_L g8479 ( 
.A1(n_7980),
.A2(n_6913),
.A3(n_6904),
.B(n_6698),
.Y(n_8479)
);

AOI22x1_ASAP7_75t_L g8480 ( 
.A1(n_7782),
.A2(n_6778),
.B1(n_6876),
.B2(n_6605),
.Y(n_8480)
);

BUFx3_ASAP7_75t_L g8481 ( 
.A(n_7954),
.Y(n_8481)
);

AND2x2_ASAP7_75t_L g8482 ( 
.A(n_7254),
.B(n_6430),
.Y(n_8482)
);

INVx1_ASAP7_75t_L g8483 ( 
.A(n_7120),
.Y(n_8483)
);

CKINVDCx5p33_ASAP7_75t_R g8484 ( 
.A(n_7379),
.Y(n_8484)
);

NOR2xp33_ASAP7_75t_L g8485 ( 
.A(n_7882),
.B(n_6699),
.Y(n_8485)
);

OAI22x1_ASAP7_75t_L g8486 ( 
.A1(n_7719),
.A2(n_6710),
.B1(n_6744),
.B2(n_6731),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7120),
.Y(n_8487)
);

BUFx3_ASAP7_75t_L g8488 ( 
.A(n_7954),
.Y(n_8488)
);

INVx1_ASAP7_75t_L g8489 ( 
.A(n_7129),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_7254),
.B(n_6201),
.Y(n_8490)
);

OAI21x1_ASAP7_75t_L g8491 ( 
.A1(n_7870),
.A2(n_6041),
.B(n_6006),
.Y(n_8491)
);

INVxp33_ASAP7_75t_L g8492 ( 
.A(n_7753),
.Y(n_8492)
);

NOR2xp67_ASAP7_75t_L g8493 ( 
.A(n_7134),
.B(n_6105),
.Y(n_8493)
);

INVx3_ASAP7_75t_L g8494 ( 
.A(n_7540),
.Y(n_8494)
);

AOI21x1_ASAP7_75t_L g8495 ( 
.A1(n_7676),
.A2(n_6918),
.B(n_6912),
.Y(n_8495)
);

OAI21x1_ASAP7_75t_L g8496 ( 
.A1(n_7922),
.A2(n_6041),
.B(n_6006),
.Y(n_8496)
);

INVx2_ASAP7_75t_L g8497 ( 
.A(n_7130),
.Y(n_8497)
);

BUFx6f_ASAP7_75t_L g8498 ( 
.A(n_6926),
.Y(n_8498)
);

OAI21x1_ASAP7_75t_L g8499 ( 
.A1(n_7922),
.A2(n_6006),
.B(n_6632),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_7129),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7129),
.Y(n_8501)
);

OR2x6_ASAP7_75t_L g8502 ( 
.A(n_8110),
.B(n_6270),
.Y(n_8502)
);

NAND3xp33_ASAP7_75t_L g8503 ( 
.A(n_7827),
.B(n_6919),
.C(n_6889),
.Y(n_8503)
);

CKINVDCx5p33_ASAP7_75t_R g8504 ( 
.A(n_7379),
.Y(n_8504)
);

AO31x2_ASAP7_75t_L g8505 ( 
.A1(n_7980),
.A2(n_6913),
.A3(n_6904),
.B(n_6698),
.Y(n_8505)
);

OAI221xp5_ASAP7_75t_L g8506 ( 
.A1(n_7490),
.A2(n_5845),
.B1(n_6874),
.B2(n_5758),
.C(n_6457),
.Y(n_8506)
);

NOR2x1_ASAP7_75t_L g8507 ( 
.A(n_7012),
.B(n_6433),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_7130),
.Y(n_8508)
);

OAI21x1_ASAP7_75t_L g8509 ( 
.A1(n_7028),
.A2(n_6654),
.B(n_6632),
.Y(n_8509)
);

AND2x2_ASAP7_75t_L g8510 ( 
.A(n_7254),
.B(n_6201),
.Y(n_8510)
);

AOI222xp33_ASAP7_75t_L g8511 ( 
.A1(n_7395),
.A2(n_5920),
.B1(n_5925),
.B2(n_6513),
.C1(n_6510),
.C2(n_6718),
.Y(n_8511)
);

AO21x2_ASAP7_75t_L g8512 ( 
.A1(n_7146),
.A2(n_6749),
.B(n_6644),
.Y(n_8512)
);

OAI21x1_ASAP7_75t_L g8513 ( 
.A1(n_7028),
.A2(n_6654),
.B(n_6720),
.Y(n_8513)
);

INVx3_ASAP7_75t_L g8514 ( 
.A(n_7540),
.Y(n_8514)
);

OAI21x1_ASAP7_75t_L g8515 ( 
.A1(n_7028),
.A2(n_6720),
.B(n_6627),
.Y(n_8515)
);

INVx1_ASAP7_75t_L g8516 ( 
.A(n_7133),
.Y(n_8516)
);

CKINVDCx20_ASAP7_75t_R g8517 ( 
.A(n_7421),
.Y(n_8517)
);

AND2x4_ASAP7_75t_L g8518 ( 
.A(n_7224),
.B(n_6193),
.Y(n_8518)
);

OAI21x1_ASAP7_75t_L g8519 ( 
.A1(n_7947),
.A2(n_6720),
.B(n_6627),
.Y(n_8519)
);

INVxp67_ASAP7_75t_L g8520 ( 
.A(n_7459),
.Y(n_8520)
);

OAI21xp5_ASAP7_75t_L g8521 ( 
.A1(n_7384),
.A2(n_5860),
.B(n_5898),
.Y(n_8521)
);

INVx2_ASAP7_75t_SL g8522 ( 
.A(n_7389),
.Y(n_8522)
);

OAI21x1_ASAP7_75t_L g8523 ( 
.A1(n_7947),
.A2(n_6720),
.B(n_6620),
.Y(n_8523)
);

INVx3_ASAP7_75t_SL g8524 ( 
.A(n_7501),
.Y(n_8524)
);

AND2x2_ASAP7_75t_L g8525 ( 
.A(n_6958),
.B(n_6201),
.Y(n_8525)
);

AOI21xp5_ASAP7_75t_L g8526 ( 
.A1(n_7980),
.A2(n_6322),
.B(n_6725),
.Y(n_8526)
);

OAI21x1_ASAP7_75t_L g8527 ( 
.A1(n_7769),
.A2(n_7793),
.B(n_7563),
.Y(n_8527)
);

OAI21x1_ASAP7_75t_L g8528 ( 
.A1(n_7769),
.A2(n_6620),
.B(n_5937),
.Y(n_8528)
);

AOI21xp5_ASAP7_75t_L g8529 ( 
.A1(n_7980),
.A2(n_6735),
.B(n_6725),
.Y(n_8529)
);

OA21x2_ASAP7_75t_L g8530 ( 
.A1(n_7223),
.A2(n_6749),
.B(n_6773),
.Y(n_8530)
);

INVx2_ASAP7_75t_L g8531 ( 
.A(n_7131),
.Y(n_8531)
);

INVxp67_ASAP7_75t_L g8532 ( 
.A(n_7459),
.Y(n_8532)
);

INVx1_ASAP7_75t_L g8533 ( 
.A(n_7133),
.Y(n_8533)
);

OAI21x1_ASAP7_75t_L g8534 ( 
.A1(n_7769),
.A2(n_5937),
.B(n_6615),
.Y(n_8534)
);

CKINVDCx5p33_ASAP7_75t_R g8535 ( 
.A(n_6941),
.Y(n_8535)
);

AOI21xp5_ASAP7_75t_L g8536 ( 
.A1(n_7050),
.A2(n_7869),
.B(n_7072),
.Y(n_8536)
);

OA21x2_ASAP7_75t_L g8537 ( 
.A1(n_7223),
.A2(n_6798),
.B(n_6773),
.Y(n_8537)
);

AND2x2_ASAP7_75t_L g8538 ( 
.A(n_6958),
.B(n_6203),
.Y(n_8538)
);

OAI21x1_ASAP7_75t_L g8539 ( 
.A1(n_7793),
.A2(n_6615),
.B(n_5831),
.Y(n_8539)
);

INVx1_ASAP7_75t_L g8540 ( 
.A(n_7133),
.Y(n_8540)
);

OAI21x1_ASAP7_75t_L g8541 ( 
.A1(n_7793),
.A2(n_5831),
.B(n_6590),
.Y(n_8541)
);

INVx3_ASAP7_75t_L g8542 ( 
.A(n_7540),
.Y(n_8542)
);

OAI21x1_ASAP7_75t_L g8543 ( 
.A1(n_7563),
.A2(n_6644),
.B(n_6590),
.Y(n_8543)
);

BUFx2_ASAP7_75t_SL g8544 ( 
.A(n_7157),
.Y(n_8544)
);

CKINVDCx20_ASAP7_75t_R g8545 ( 
.A(n_7422),
.Y(n_8545)
);

INVx2_ASAP7_75t_L g8546 ( 
.A(n_7131),
.Y(n_8546)
);

OAI21x1_ASAP7_75t_L g8547 ( 
.A1(n_7563),
.A2(n_6705),
.B(n_6676),
.Y(n_8547)
);

OAI22xp33_ASAP7_75t_L g8548 ( 
.A1(n_8113),
.A2(n_7782),
.B1(n_7796),
.B2(n_7824),
.Y(n_8548)
);

AOI21xp5_ASAP7_75t_L g8549 ( 
.A1(n_7050),
.A2(n_6736),
.B(n_6735),
.Y(n_8549)
);

AO21x2_ASAP7_75t_L g8550 ( 
.A1(n_7146),
.A2(n_6705),
.B(n_6676),
.Y(n_8550)
);

AOI22xp5_ASAP7_75t_L g8551 ( 
.A1(n_7515),
.A2(n_5848),
.B1(n_5925),
.B2(n_5920),
.Y(n_8551)
);

AO21x2_ASAP7_75t_L g8552 ( 
.A1(n_7146),
.A2(n_6758),
.B(n_6756),
.Y(n_8552)
);

INVx1_ASAP7_75t_L g8553 ( 
.A(n_7136),
.Y(n_8553)
);

OAI22xp5_ASAP7_75t_L g8554 ( 
.A1(n_7782),
.A2(n_6669),
.B1(n_6700),
.B2(n_6648),
.Y(n_8554)
);

AND2x4_ASAP7_75t_L g8555 ( 
.A(n_7224),
.B(n_6195),
.Y(n_8555)
);

O2A1O1Ixp33_ASAP7_75t_SL g8556 ( 
.A1(n_7179),
.A2(n_6736),
.B(n_6829),
.C(n_6765),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_7136),
.Y(n_8557)
);

AO21x1_ASAP7_75t_L g8558 ( 
.A1(n_7072),
.A2(n_6239),
.B(n_6236),
.Y(n_8558)
);

AND2x2_ASAP7_75t_L g8559 ( 
.A(n_6958),
.B(n_6203),
.Y(n_8559)
);

OAI21x1_ASAP7_75t_L g8560 ( 
.A1(n_7563),
.A2(n_6758),
.B(n_6756),
.Y(n_8560)
);

OA21x2_ASAP7_75t_L g8561 ( 
.A1(n_7223),
.A2(n_6808),
.B(n_6798),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_7136),
.Y(n_8562)
);

OAI22xp33_ASAP7_75t_L g8563 ( 
.A1(n_8113),
.A2(n_7796),
.B1(n_7849),
.B2(n_7824),
.Y(n_8563)
);

NAND2x1p5_ASAP7_75t_L g8564 ( 
.A(n_7317),
.B(n_6416),
.Y(n_8564)
);

AOI22xp33_ASAP7_75t_L g8565 ( 
.A1(n_7515),
.A2(n_7179),
.B1(n_8112),
.B2(n_7745),
.Y(n_8565)
);

AOI21xp5_ASAP7_75t_L g8566 ( 
.A1(n_7072),
.A2(n_6829),
.B(n_6765),
.Y(n_8566)
);

OAI21x1_ASAP7_75t_L g8567 ( 
.A1(n_7213),
.A2(n_6787),
.B(n_6779),
.Y(n_8567)
);

OAI21x1_ASAP7_75t_L g8568 ( 
.A1(n_7213),
.A2(n_7400),
.B(n_7248),
.Y(n_8568)
);

O2A1O1Ixp33_ASAP7_75t_L g8569 ( 
.A1(n_7679),
.A2(n_5830),
.B(n_5990),
.C(n_5811),
.Y(n_8569)
);

HB1xp67_ASAP7_75t_L g8570 ( 
.A(n_7437),
.Y(n_8570)
);

OA21x2_ASAP7_75t_L g8571 ( 
.A1(n_7653),
.A2(n_6808),
.B(n_6218),
.Y(n_8571)
);

AO31x2_ASAP7_75t_L g8572 ( 
.A1(n_7653),
.A2(n_6743),
.A3(n_6755),
.B(n_6718),
.Y(n_8572)
);

AND2x4_ASAP7_75t_L g8573 ( 
.A(n_7224),
.B(n_6195),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_7151),
.Y(n_8574)
);

OAI21xp5_ASAP7_75t_L g8575 ( 
.A1(n_7384),
.A2(n_6874),
.B(n_5791),
.Y(n_8575)
);

AO31x2_ASAP7_75t_L g8576 ( 
.A1(n_7653),
.A2(n_6755),
.A3(n_6772),
.B(n_6743),
.Y(n_8576)
);

AO32x2_ASAP7_75t_L g8577 ( 
.A1(n_8024),
.A2(n_8036),
.A3(n_6772),
.B1(n_8043),
.B2(n_7182),
.Y(n_8577)
);

INVx2_ASAP7_75t_SL g8578 ( 
.A(n_7389),
.Y(n_8578)
);

NAND2xp5_ASAP7_75t_L g8579 ( 
.A(n_7132),
.B(n_6101),
.Y(n_8579)
);

AOI21xp33_ASAP7_75t_L g8580 ( 
.A1(n_7827),
.A2(n_6258),
.B(n_6110),
.Y(n_8580)
);

AND2x4_ASAP7_75t_L g8581 ( 
.A(n_7389),
.B(n_6195),
.Y(n_8581)
);

OAI22xp5_ASAP7_75t_L g8582 ( 
.A1(n_7796),
.A2(n_6669),
.B1(n_6700),
.B2(n_6648),
.Y(n_8582)
);

OAI21x1_ASAP7_75t_L g8583 ( 
.A1(n_7213),
.A2(n_6787),
.B(n_6779),
.Y(n_8583)
);

NAND2xp5_ASAP7_75t_SL g8584 ( 
.A(n_7932),
.B(n_5910),
.Y(n_8584)
);

OAI21x1_ASAP7_75t_L g8585 ( 
.A1(n_7248),
.A2(n_6507),
.B(n_6385),
.Y(n_8585)
);

OR2x2_ASAP7_75t_L g8586 ( 
.A(n_8024),
.B(n_6101),
.Y(n_8586)
);

BUFx12f_ASAP7_75t_L g8587 ( 
.A(n_8044),
.Y(n_8587)
);

INVx2_ASAP7_75t_SL g8588 ( 
.A(n_7389),
.Y(n_8588)
);

NAND2xp5_ASAP7_75t_L g8589 ( 
.A(n_7132),
.B(n_6114),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_7151),
.Y(n_8590)
);

NAND3xp33_ASAP7_75t_L g8591 ( 
.A(n_7869),
.B(n_6699),
.C(n_6592),
.Y(n_8591)
);

OAI21x1_ASAP7_75t_L g8592 ( 
.A1(n_7248),
.A2(n_6507),
.B(n_6385),
.Y(n_8592)
);

O2A1O1Ixp33_ASAP7_75t_L g8593 ( 
.A1(n_7679),
.A2(n_5830),
.B(n_5990),
.C(n_5811),
.Y(n_8593)
);

INVxp67_ASAP7_75t_SL g8594 ( 
.A(n_7677),
.Y(n_8594)
);

OAI21x1_ASAP7_75t_L g8595 ( 
.A1(n_7400),
.A2(n_6507),
.B(n_6897),
.Y(n_8595)
);

BUFx3_ASAP7_75t_L g8596 ( 
.A(n_7022),
.Y(n_8596)
);

NAND2x1p5_ASAP7_75t_L g8597 ( 
.A(n_7636),
.B(n_6416),
.Y(n_8597)
);

BUFx8_ASAP7_75t_L g8598 ( 
.A(n_7022),
.Y(n_8598)
);

OAI21x1_ASAP7_75t_L g8599 ( 
.A1(n_8017),
.A2(n_7920),
.B(n_7898),
.Y(n_8599)
);

INVx1_ASAP7_75t_L g8600 ( 
.A(n_7151),
.Y(n_8600)
);

INVx1_ASAP7_75t_L g8601 ( 
.A(n_7153),
.Y(n_8601)
);

CKINVDCx9p33_ASAP7_75t_R g8602 ( 
.A(n_7679),
.Y(n_8602)
);

OAI21x1_ASAP7_75t_SL g8603 ( 
.A1(n_7087),
.A2(n_6878),
.B(n_6860),
.Y(n_8603)
);

OAI221xp5_ASAP7_75t_L g8604 ( 
.A1(n_8034),
.A2(n_5772),
.B1(n_6387),
.B2(n_6717),
.C(n_6510),
.Y(n_8604)
);

BUFx3_ASAP7_75t_L g8605 ( 
.A(n_7022),
.Y(n_8605)
);

NOR2xp33_ASAP7_75t_L g8606 ( 
.A(n_7562),
.B(n_5918),
.Y(n_8606)
);

NOR2xp67_ASAP7_75t_L g8607 ( 
.A(n_7154),
.B(n_6105),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_7153),
.Y(n_8608)
);

AOI22xp33_ASAP7_75t_L g8609 ( 
.A1(n_8112),
.A2(n_6215),
.B1(n_5955),
.B2(n_6543),
.Y(n_8609)
);

NAND2x1p5_ASAP7_75t_L g8610 ( 
.A(n_7636),
.B(n_6416),
.Y(n_8610)
);

INVx2_ASAP7_75t_SL g8611 ( 
.A(n_7449),
.Y(n_8611)
);

HB1xp67_ASAP7_75t_L g8612 ( 
.A(n_7437),
.Y(n_8612)
);

OA21x2_ASAP7_75t_L g8613 ( 
.A1(n_8017),
.A2(n_6218),
.B(n_6208),
.Y(n_8613)
);

OAI22xp5_ASAP7_75t_L g8614 ( 
.A1(n_7796),
.A2(n_6700),
.B1(n_6522),
.B2(n_6548),
.Y(n_8614)
);

OAI21x1_ASAP7_75t_L g8615 ( 
.A1(n_8017),
.A2(n_6507),
.B(n_6897),
.Y(n_8615)
);

OAI22xp5_ASAP7_75t_L g8616 ( 
.A1(n_7971),
.A2(n_6522),
.B1(n_6548),
.B2(n_6203),
.Y(n_8616)
);

OAI22x1_ASAP7_75t_L g8617 ( 
.A1(n_7719),
.A2(n_6710),
.B1(n_6744),
.B2(n_6731),
.Y(n_8617)
);

INVx3_ASAP7_75t_L g8618 ( 
.A(n_7797),
.Y(n_8618)
);

INVx3_ASAP7_75t_SL g8619 ( 
.A(n_7501),
.Y(n_8619)
);

OAI21xp5_ASAP7_75t_L g8620 ( 
.A1(n_7385),
.A2(n_5791),
.B(n_5886),
.Y(n_8620)
);

OA21x2_ASAP7_75t_L g8621 ( 
.A1(n_7229),
.A2(n_6018),
.B(n_6236),
.Y(n_8621)
);

AOI22xp5_ASAP7_75t_L g8622 ( 
.A1(n_7692),
.A2(n_5772),
.B1(n_6434),
.B2(n_6475),
.Y(n_8622)
);

INVx3_ASAP7_75t_L g8623 ( 
.A(n_7797),
.Y(n_8623)
);

OAI21xp5_ASAP7_75t_L g8624 ( 
.A1(n_7385),
.A2(n_5886),
.B(n_6008),
.Y(n_8624)
);

OAI21x1_ASAP7_75t_L g8625 ( 
.A1(n_7898),
.A2(n_7920),
.B(n_7718),
.Y(n_8625)
);

INVx2_ASAP7_75t_SL g8626 ( 
.A(n_7449),
.Y(n_8626)
);

INVx4_ASAP7_75t_SL g8627 ( 
.A(n_7393),
.Y(n_8627)
);

NOR2x1_ASAP7_75t_SL g8628 ( 
.A(n_7336),
.B(n_7344),
.Y(n_8628)
);

INVx1_ASAP7_75t_L g8629 ( 
.A(n_7153),
.Y(n_8629)
);

INVx4_ASAP7_75t_L g8630 ( 
.A(n_7138),
.Y(n_8630)
);

INVx2_ASAP7_75t_L g8631 ( 
.A(n_7131),
.Y(n_8631)
);

OR2x2_ASAP7_75t_L g8632 ( 
.A(n_8036),
.B(n_6114),
.Y(n_8632)
);

AND2x2_ASAP7_75t_L g8633 ( 
.A(n_6958),
.B(n_6140),
.Y(n_8633)
);

AOI21xp33_ASAP7_75t_SL g8634 ( 
.A1(n_6980),
.A2(n_6733),
.B(n_5699),
.Y(n_8634)
);

BUFx2_ASAP7_75t_L g8635 ( 
.A(n_7930),
.Y(n_8635)
);

BUFx2_ASAP7_75t_L g8636 ( 
.A(n_7930),
.Y(n_8636)
);

AOI22xp5_ASAP7_75t_L g8637 ( 
.A1(n_7692),
.A2(n_8112),
.B1(n_7598),
.B2(n_8034),
.Y(n_8637)
);

INVx1_ASAP7_75t_L g8638 ( 
.A(n_7165),
.Y(n_8638)
);

INVx2_ASAP7_75t_L g8639 ( 
.A(n_7131),
.Y(n_8639)
);

OA21x2_ASAP7_75t_L g8640 ( 
.A1(n_7229),
.A2(n_6018),
.B(n_6239),
.Y(n_8640)
);

OAI21x1_ASAP7_75t_L g8641 ( 
.A1(n_7920),
.A2(n_6820),
.B(n_6795),
.Y(n_8641)
);

AOI21xp5_ASAP7_75t_L g8642 ( 
.A1(n_7869),
.A2(n_6871),
.B(n_5750),
.Y(n_8642)
);

AOI22xp5_ASAP7_75t_L g8643 ( 
.A1(n_7692),
.A2(n_6434),
.B1(n_6475),
.B2(n_6576),
.Y(n_8643)
);

CKINVDCx6p67_ASAP7_75t_R g8644 ( 
.A(n_7093),
.Y(n_8644)
);

INVx1_ASAP7_75t_L g8645 ( 
.A(n_7165),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_7165),
.Y(n_8646)
);

NAND3xp33_ASAP7_75t_L g8647 ( 
.A(n_7598),
.B(n_6592),
.C(n_6585),
.Y(n_8647)
);

OAI21x1_ASAP7_75t_L g8648 ( 
.A1(n_7920),
.A2(n_6820),
.B(n_6795),
.Y(n_8648)
);

BUFx4f_ASAP7_75t_L g8649 ( 
.A(n_7093),
.Y(n_8649)
);

OAI21x1_ASAP7_75t_L g8650 ( 
.A1(n_7718),
.A2(n_6887),
.B(n_6852),
.Y(n_8650)
);

CKINVDCx5p33_ASAP7_75t_R g8651 ( 
.A(n_6941),
.Y(n_8651)
);

AO31x2_ASAP7_75t_L g8652 ( 
.A1(n_7986),
.A2(n_6247),
.A3(n_6259),
.B(n_6246),
.Y(n_8652)
);

OAI221xp5_ASAP7_75t_L g8653 ( 
.A1(n_8034),
.A2(n_6717),
.B1(n_6745),
.B2(n_6543),
.C(n_6014),
.Y(n_8653)
);

INVx2_ASAP7_75t_SL g8654 ( 
.A(n_7449),
.Y(n_8654)
);

OAI21x1_ASAP7_75t_L g8655 ( 
.A1(n_7718),
.A2(n_6887),
.B(n_6852),
.Y(n_8655)
);

AOI22xp33_ASAP7_75t_L g8656 ( 
.A1(n_7745),
.A2(n_5955),
.B1(n_6543),
.B2(n_6270),
.Y(n_8656)
);

AOI22xp33_ASAP7_75t_L g8657 ( 
.A1(n_7745),
.A2(n_5955),
.B1(n_6543),
.B2(n_6270),
.Y(n_8657)
);

A2O1A1Ixp33_ASAP7_75t_L g8658 ( 
.A1(n_7044),
.A2(n_6252),
.B(n_5764),
.C(n_6017),
.Y(n_8658)
);

OA21x2_ASAP7_75t_L g8659 ( 
.A1(n_7229),
.A2(n_6247),
.B(n_6246),
.Y(n_8659)
);

INVx1_ASAP7_75t_L g8660 ( 
.A(n_7168),
.Y(n_8660)
);

OAI22xp5_ASAP7_75t_L g8661 ( 
.A1(n_7971),
.A2(n_6155),
.B1(n_6189),
.B2(n_6140),
.Y(n_8661)
);

AOI22xp33_ASAP7_75t_L g8662 ( 
.A1(n_7431),
.A2(n_5955),
.B1(n_6543),
.B2(n_6230),
.Y(n_8662)
);

OA21x2_ASAP7_75t_L g8663 ( 
.A1(n_7236),
.A2(n_6288),
.B(n_6259),
.Y(n_8663)
);

INVx1_ASAP7_75t_SL g8664 ( 
.A(n_7678),
.Y(n_8664)
);

AOI221xp5_ASAP7_75t_L g8665 ( 
.A1(n_8036),
.A2(n_6014),
.B1(n_6008),
.B2(n_6293),
.C(n_6288),
.Y(n_8665)
);

OR2x6_ASAP7_75t_L g8666 ( 
.A(n_8110),
.B(n_6332),
.Y(n_8666)
);

OAI21xp5_ASAP7_75t_L g8667 ( 
.A1(n_7974),
.A2(n_5781),
.B(n_5750),
.Y(n_8667)
);

OAI22xp33_ASAP7_75t_L g8668 ( 
.A1(n_7824),
.A2(n_6745),
.B1(n_6810),
.B2(n_6614),
.Y(n_8668)
);

NOR2xp33_ASAP7_75t_L g8669 ( 
.A(n_7562),
.B(n_5918),
.Y(n_8669)
);

INVx1_ASAP7_75t_L g8670 ( 
.A(n_7168),
.Y(n_8670)
);

BUFx4_ASAP7_75t_R g8671 ( 
.A(n_7816),
.Y(n_8671)
);

AND2x6_ASAP7_75t_L g8672 ( 
.A(n_7795),
.B(n_5989),
.Y(n_8672)
);

OR2x6_ASAP7_75t_L g8673 ( 
.A(n_8110),
.B(n_6332),
.Y(n_8673)
);

OAI211xp5_ASAP7_75t_L g8674 ( 
.A1(n_7813),
.A2(n_6910),
.B(n_6733),
.C(n_5939),
.Y(n_8674)
);

BUFx6f_ASAP7_75t_L g8675 ( 
.A(n_6926),
.Y(n_8675)
);

INVx1_ASAP7_75t_L g8676 ( 
.A(n_7168),
.Y(n_8676)
);

HB1xp67_ASAP7_75t_L g8677 ( 
.A(n_7442),
.Y(n_8677)
);

AND2x2_ASAP7_75t_L g8678 ( 
.A(n_6958),
.B(n_6140),
.Y(n_8678)
);

OAI21x1_ASAP7_75t_L g8679 ( 
.A1(n_7654),
.A2(n_6074),
.B(n_6019),
.Y(n_8679)
);

OAI22xp5_ASAP7_75t_L g8680 ( 
.A1(n_7987),
.A2(n_6189),
.B1(n_6155),
.B2(n_6922),
.Y(n_8680)
);

BUFx12f_ASAP7_75t_L g8681 ( 
.A(n_6980),
.Y(n_8681)
);

OAI21x1_ASAP7_75t_L g8682 ( 
.A1(n_7654),
.A2(n_7837),
.B(n_7716),
.Y(n_8682)
);

INVx1_ASAP7_75t_L g8683 ( 
.A(n_7199),
.Y(n_8683)
);

OAI21x1_ASAP7_75t_L g8684 ( 
.A1(n_7654),
.A2(n_6074),
.B(n_6019),
.Y(n_8684)
);

INVx1_ASAP7_75t_L g8685 ( 
.A(n_7199),
.Y(n_8685)
);

AOI21xp5_ASAP7_75t_L g8686 ( 
.A1(n_8086),
.A2(n_6871),
.B(n_5736),
.Y(n_8686)
);

AOI21xp5_ASAP7_75t_L g8687 ( 
.A1(n_8086),
.A2(n_5736),
.B(n_6862),
.Y(n_8687)
);

INVx3_ASAP7_75t_L g8688 ( 
.A(n_7797),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_7199),
.Y(n_8689)
);

AO21x2_ASAP7_75t_L g8690 ( 
.A1(n_7146),
.A2(n_5416),
.B(n_5406),
.Y(n_8690)
);

OA21x2_ASAP7_75t_L g8691 ( 
.A1(n_7236),
.A2(n_7256),
.B(n_7237),
.Y(n_8691)
);

AOI22xp33_ASAP7_75t_SL g8692 ( 
.A1(n_7063),
.A2(n_6319),
.B1(n_6308),
.B2(n_5976),
.Y(n_8692)
);

OAI21x1_ASAP7_75t_L g8693 ( 
.A1(n_7837),
.A2(n_6074),
.B(n_6019),
.Y(n_8693)
);

AO32x2_ASAP7_75t_L g8694 ( 
.A1(n_8043),
.A2(n_5764),
.A3(n_6898),
.B1(n_6816),
.B2(n_6762),
.Y(n_8694)
);

AND2x4_ASAP7_75t_L g8695 ( 
.A(n_7449),
.B(n_6195),
.Y(n_8695)
);

INVx1_ASAP7_75t_L g8696 ( 
.A(n_7207),
.Y(n_8696)
);

NAND2x1p5_ASAP7_75t_L g8697 ( 
.A(n_7636),
.B(n_6416),
.Y(n_8697)
);

INVx3_ASAP7_75t_L g8698 ( 
.A(n_7797),
.Y(n_8698)
);

INVx2_ASAP7_75t_L g8699 ( 
.A(n_7142),
.Y(n_8699)
);

OR2x6_ASAP7_75t_L g8700 ( 
.A(n_8118),
.B(n_6332),
.Y(n_8700)
);

INVx1_ASAP7_75t_L g8701 ( 
.A(n_7207),
.Y(n_8701)
);

INVx1_ASAP7_75t_SL g8702 ( 
.A(n_7678),
.Y(n_8702)
);

OA21x2_ASAP7_75t_L g8703 ( 
.A1(n_7236),
.A2(n_6309),
.B(n_6293),
.Y(n_8703)
);

INVx6_ASAP7_75t_L g8704 ( 
.A(n_7568),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_7142),
.Y(n_8705)
);

OAI21x1_ASAP7_75t_L g8706 ( 
.A1(n_7837),
.A2(n_7716),
.B(n_7814),
.Y(n_8706)
);

A2O1A1Ixp33_ASAP7_75t_L g8707 ( 
.A1(n_7044),
.A2(n_6252),
.B(n_5764),
.C(n_6243),
.Y(n_8707)
);

OAI21x1_ASAP7_75t_L g8708 ( 
.A1(n_7716),
.A2(n_6074),
.B(n_6019),
.Y(n_8708)
);

INVx1_ASAP7_75t_SL g8709 ( 
.A(n_7001),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_7207),
.Y(n_8710)
);

INVx6_ASAP7_75t_L g8711 ( 
.A(n_7568),
.Y(n_8711)
);

INVx2_ASAP7_75t_L g8712 ( 
.A(n_7142),
.Y(n_8712)
);

OAI21x1_ASAP7_75t_L g8713 ( 
.A1(n_7814),
.A2(n_6888),
.B(n_6862),
.Y(n_8713)
);

INVx2_ASAP7_75t_L g8714 ( 
.A(n_7142),
.Y(n_8714)
);

OAI211xp5_ASAP7_75t_L g8715 ( 
.A1(n_7813),
.A2(n_6910),
.B(n_5939),
.C(n_6063),
.Y(n_8715)
);

AOI22xp33_ASAP7_75t_L g8716 ( 
.A1(n_7431),
.A2(n_5955),
.B1(n_6543),
.B2(n_6230),
.Y(n_8716)
);

BUFx3_ASAP7_75t_L g8717 ( 
.A(n_7093),
.Y(n_8717)
);

OAI21xp5_ASAP7_75t_L g8718 ( 
.A1(n_7974),
.A2(n_7965),
.B(n_7293),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_7233),
.Y(n_8719)
);

INVx4_ASAP7_75t_SL g8720 ( 
.A(n_7393),
.Y(n_8720)
);

INVx1_ASAP7_75t_L g8721 ( 
.A(n_7233),
.Y(n_8721)
);

CKINVDCx5p33_ASAP7_75t_R g8722 ( 
.A(n_7729),
.Y(n_8722)
);

INVx1_ASAP7_75t_L g8723 ( 
.A(n_7233),
.Y(n_8723)
);

NOR2xp33_ASAP7_75t_SL g8724 ( 
.A(n_7413),
.B(n_6020),
.Y(n_8724)
);

OAI21x1_ASAP7_75t_L g8725 ( 
.A1(n_7814),
.A2(n_6905),
.B(n_6888),
.Y(n_8725)
);

OAI21x1_ASAP7_75t_L g8726 ( 
.A1(n_7830),
.A2(n_6905),
.B(n_6549),
.Y(n_8726)
);

AOI21xp5_ASAP7_75t_L g8727 ( 
.A1(n_7598),
.A2(n_5781),
.B(n_6230),
.Y(n_8727)
);

NAND2xp5_ASAP7_75t_L g8728 ( 
.A(n_7132),
.B(n_6121),
.Y(n_8728)
);

AO21x2_ASAP7_75t_L g8729 ( 
.A1(n_7146),
.A2(n_5416),
.B(n_5406),
.Y(n_8729)
);

INVx1_ASAP7_75t_L g8730 ( 
.A(n_7238),
.Y(n_8730)
);

OAI21xp5_ASAP7_75t_L g8731 ( 
.A1(n_7974),
.A2(n_6752),
.B(n_6739),
.Y(n_8731)
);

INVx2_ASAP7_75t_L g8732 ( 
.A(n_7152),
.Y(n_8732)
);

AOI22xp33_ASAP7_75t_L g8733 ( 
.A1(n_7441),
.A2(n_5955),
.B1(n_6543),
.B2(n_6230),
.Y(n_8733)
);

OAI21xp5_ASAP7_75t_L g8734 ( 
.A1(n_7965),
.A2(n_6752),
.B(n_6739),
.Y(n_8734)
);

AOI21xp5_ASAP7_75t_L g8735 ( 
.A1(n_7905),
.A2(n_6230),
.B(n_6335),
.Y(n_8735)
);

OAI21x1_ASAP7_75t_L g8736 ( 
.A1(n_7761),
.A2(n_6549),
.B(n_6530),
.Y(n_8736)
);

NAND2xp5_ASAP7_75t_L g8737 ( 
.A(n_7145),
.B(n_6121),
.Y(n_8737)
);

HB1xp67_ASAP7_75t_L g8738 ( 
.A(n_7442),
.Y(n_8738)
);

OAI21x1_ASAP7_75t_L g8739 ( 
.A1(n_7761),
.A2(n_6549),
.B(n_6530),
.Y(n_8739)
);

INVxp67_ASAP7_75t_SL g8740 ( 
.A(n_7677),
.Y(n_8740)
);

OA21x2_ASAP7_75t_L g8741 ( 
.A1(n_7237),
.A2(n_6317),
.B(n_6309),
.Y(n_8741)
);

AND2x4_ASAP7_75t_L g8742 ( 
.A(n_7464),
.B(n_6195),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_7238),
.Y(n_8743)
);

OR2x2_ASAP7_75t_L g8744 ( 
.A(n_7475),
.B(n_7390),
.Y(n_8744)
);

AOI221x1_ASAP7_75t_L g8745 ( 
.A1(n_7063),
.A2(n_5834),
.B1(n_5849),
.B2(n_5842),
.C(n_5835),
.Y(n_8745)
);

AOI22x1_ASAP7_75t_L g8746 ( 
.A1(n_8031),
.A2(n_6876),
.B1(n_6901),
.B2(n_6373),
.Y(n_8746)
);

CKINVDCx11_ASAP7_75t_R g8747 ( 
.A(n_7422),
.Y(n_8747)
);

OAI21x1_ASAP7_75t_L g8748 ( 
.A1(n_7761),
.A2(n_6575),
.B(n_6530),
.Y(n_8748)
);

BUFx2_ASAP7_75t_L g8749 ( 
.A(n_7930),
.Y(n_8749)
);

AOI22xp33_ASAP7_75t_L g8750 ( 
.A1(n_7441),
.A2(n_5955),
.B1(n_6230),
.B2(n_6170),
.Y(n_8750)
);

INVx2_ASAP7_75t_L g8751 ( 
.A(n_7152),
.Y(n_8751)
);

INVx2_ASAP7_75t_L g8752 ( 
.A(n_7152),
.Y(n_8752)
);

O2A1O1Ixp33_ASAP7_75t_SL g8753 ( 
.A1(n_7917),
.A2(n_6472),
.B(n_6484),
.C(n_6458),
.Y(n_8753)
);

OAI21x1_ASAP7_75t_L g8754 ( 
.A1(n_7778),
.A2(n_6577),
.B(n_6575),
.Y(n_8754)
);

NOR2xp33_ASAP7_75t_L g8755 ( 
.A(n_7574),
.B(n_5932),
.Y(n_8755)
);

INVx3_ASAP7_75t_SL g8756 ( 
.A(n_7045),
.Y(n_8756)
);

O2A1O1Ixp33_ASAP7_75t_L g8757 ( 
.A1(n_7679),
.A2(n_8031),
.B(n_7063),
.C(n_7099),
.Y(n_8757)
);

INVx1_ASAP7_75t_L g8758 ( 
.A(n_7238),
.Y(n_8758)
);

BUFx12f_ASAP7_75t_L g8759 ( 
.A(n_6999),
.Y(n_8759)
);

OAI21xp5_ASAP7_75t_L g8760 ( 
.A1(n_7293),
.A2(n_6809),
.B(n_6800),
.Y(n_8760)
);

OAI21xp33_ASAP7_75t_L g8761 ( 
.A1(n_7595),
.A2(n_6516),
.B(n_6499),
.Y(n_8761)
);

OAI21x1_ASAP7_75t_L g8762 ( 
.A1(n_7778),
.A2(n_6577),
.B(n_6575),
.Y(n_8762)
);

INVx1_ASAP7_75t_L g8763 ( 
.A(n_7241),
.Y(n_8763)
);

AOI21xp5_ASAP7_75t_L g8764 ( 
.A1(n_7914),
.A2(n_6230),
.B(n_6335),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_L g8765 ( 
.A(n_7145),
.B(n_6125),
.Y(n_8765)
);

BUFx12f_ASAP7_75t_L g8766 ( 
.A(n_6999),
.Y(n_8766)
);

BUFx6f_ASAP7_75t_L g8767 ( 
.A(n_6926),
.Y(n_8767)
);

OAI21x1_ASAP7_75t_L g8768 ( 
.A1(n_7778),
.A2(n_6577),
.B(n_6575),
.Y(n_8768)
);

O2A1O1Ixp33_ASAP7_75t_L g8769 ( 
.A1(n_7679),
.A2(n_6258),
.B(n_6325),
.C(n_6110),
.Y(n_8769)
);

INVx2_ASAP7_75t_L g8770 ( 
.A(n_7152),
.Y(n_8770)
);

NAND2xp5_ASAP7_75t_SL g8771 ( 
.A(n_7932),
.B(n_7978),
.Y(n_8771)
);

OAI21x1_ASAP7_75t_L g8772 ( 
.A1(n_7237),
.A2(n_6577),
.B(n_6575),
.Y(n_8772)
);

INVx6_ASAP7_75t_L g8773 ( 
.A(n_7568),
.Y(n_8773)
);

OAI21x1_ASAP7_75t_L g8774 ( 
.A1(n_7256),
.A2(n_6578),
.B(n_6577),
.Y(n_8774)
);

NAND2xp5_ASAP7_75t_L g8775 ( 
.A(n_7145),
.B(n_6125),
.Y(n_8775)
);

OAI21x1_ASAP7_75t_L g8776 ( 
.A1(n_7256),
.A2(n_6693),
.B(n_6578),
.Y(n_8776)
);

AOI22xp33_ASAP7_75t_L g8777 ( 
.A1(n_7726),
.A2(n_5955),
.B1(n_6170),
.B2(n_6105),
.Y(n_8777)
);

NAND3xp33_ASAP7_75t_L g8778 ( 
.A(n_7813),
.B(n_7774),
.C(n_7726),
.Y(n_8778)
);

O2A1O1Ixp33_ASAP7_75t_L g8779 ( 
.A1(n_8031),
.A2(n_6473),
.B(n_6529),
.C(n_6325),
.Y(n_8779)
);

INVx4_ASAP7_75t_L g8780 ( 
.A(n_7138),
.Y(n_8780)
);

AOI22xp5_ASAP7_75t_L g8781 ( 
.A1(n_7099),
.A2(n_6581),
.B1(n_6576),
.B2(n_5955),
.Y(n_8781)
);

INVx2_ASAP7_75t_L g8782 ( 
.A(n_7155),
.Y(n_8782)
);

AND2x4_ASAP7_75t_L g8783 ( 
.A(n_7464),
.B(n_6216),
.Y(n_8783)
);

BUFx12f_ASAP7_75t_L g8784 ( 
.A(n_7093),
.Y(n_8784)
);

NAND2x1p5_ASAP7_75t_L g8785 ( 
.A(n_7636),
.B(n_6416),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_7241),
.Y(n_8786)
);

OAI22xp5_ASAP7_75t_L g8787 ( 
.A1(n_7987),
.A2(n_6189),
.B1(n_6155),
.B2(n_6922),
.Y(n_8787)
);

INVx2_ASAP7_75t_L g8788 ( 
.A(n_7155),
.Y(n_8788)
);

OAI21x1_ASAP7_75t_L g8789 ( 
.A1(n_7268),
.A2(n_7334),
.B(n_7269),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_7241),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_7242),
.Y(n_8791)
);

O2A1O1Ixp33_ASAP7_75t_SL g8792 ( 
.A1(n_7917),
.A2(n_6472),
.B(n_6484),
.C(n_6458),
.Y(n_8792)
);

INVx4_ASAP7_75t_L g8793 ( 
.A(n_7138),
.Y(n_8793)
);

INVx2_ASAP7_75t_L g8794 ( 
.A(n_7155),
.Y(n_8794)
);

BUFx2_ASAP7_75t_L g8795 ( 
.A(n_7930),
.Y(n_8795)
);

OAI21x1_ASAP7_75t_SL g8796 ( 
.A1(n_7087),
.A2(n_6860),
.B(n_6818),
.Y(n_8796)
);

OA21x2_ASAP7_75t_L g8797 ( 
.A1(n_7334),
.A2(n_6329),
.B(n_6317),
.Y(n_8797)
);

AOI22xp33_ASAP7_75t_L g8798 ( 
.A1(n_7170),
.A2(n_6105),
.B1(n_6191),
.B2(n_6170),
.Y(n_8798)
);

AO21x2_ASAP7_75t_L g8799 ( 
.A1(n_6984),
.A2(n_5416),
.B(n_5406),
.Y(n_8799)
);

O2A1O1Ixp33_ASAP7_75t_L g8800 ( 
.A1(n_8031),
.A2(n_6529),
.B(n_6540),
.C(n_6473),
.Y(n_8800)
);

AOI221xp5_ASAP7_75t_L g8801 ( 
.A1(n_7630),
.A2(n_6359),
.B1(n_6362),
.B2(n_6336),
.C(n_6329),
.Y(n_8801)
);

BUFx2_ASAP7_75t_L g8802 ( 
.A(n_7930),
.Y(n_8802)
);

OR2x6_ASAP7_75t_L g8803 ( 
.A(n_8118),
.B(n_6332),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_7242),
.Y(n_8804)
);

INVx2_ASAP7_75t_SL g8805 ( 
.A(n_7464),
.Y(n_8805)
);

NOR2xp33_ASAP7_75t_L g8806 ( 
.A(n_7574),
.B(n_5932),
.Y(n_8806)
);

OAI21x1_ASAP7_75t_L g8807 ( 
.A1(n_7334),
.A2(n_7354),
.B(n_7347),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_7242),
.Y(n_8808)
);

INVx1_ASAP7_75t_L g8809 ( 
.A(n_7243),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_7243),
.Y(n_8810)
);

INVx1_ASAP7_75t_L g8811 ( 
.A(n_7243),
.Y(n_8811)
);

OAI21xp5_ASAP7_75t_L g8812 ( 
.A1(n_7420),
.A2(n_7613),
.B(n_7630),
.Y(n_8812)
);

AO21x2_ASAP7_75t_L g8813 ( 
.A1(n_6984),
.A2(n_5416),
.B(n_5406),
.Y(n_8813)
);

BUFx3_ASAP7_75t_L g8814 ( 
.A(n_7177),
.Y(n_8814)
);

NOR2xp33_ASAP7_75t_L g8815 ( 
.A(n_7100),
.B(n_6063),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_7246),
.Y(n_8816)
);

OAI22xp5_ASAP7_75t_L g8817 ( 
.A1(n_7480),
.A2(n_6922),
.B1(n_6818),
.B2(n_6581),
.Y(n_8817)
);

NOR2x1_ASAP7_75t_SL g8818 ( 
.A(n_7336),
.B(n_6017),
.Y(n_8818)
);

INVx3_ASAP7_75t_L g8819 ( 
.A(n_7797),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_L g8820 ( 
.A(n_7006),
.B(n_6156),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_7246),
.Y(n_8821)
);

OR2x2_ASAP7_75t_L g8822 ( 
.A(n_7475),
.B(n_6156),
.Y(n_8822)
);

OA21x2_ASAP7_75t_L g8823 ( 
.A1(n_7347),
.A2(n_6359),
.B(n_6336),
.Y(n_8823)
);

OAI22xp5_ASAP7_75t_L g8824 ( 
.A1(n_7480),
.A2(n_6009),
.B1(n_6144),
.B2(n_6095),
.Y(n_8824)
);

INVx2_ASAP7_75t_L g8825 ( 
.A(n_7155),
.Y(n_8825)
);

INVxp67_ASAP7_75t_SL g8826 ( 
.A(n_7677),
.Y(n_8826)
);

AOI22xp5_ASAP7_75t_L g8827 ( 
.A1(n_7099),
.A2(n_6614),
.B1(n_4604),
.B2(n_6810),
.Y(n_8827)
);

AOI21x1_ASAP7_75t_L g8828 ( 
.A1(n_7913),
.A2(n_5756),
.B(n_5744),
.Y(n_8828)
);

AOI22xp5_ASAP7_75t_L g8829 ( 
.A1(n_7713),
.A2(n_6565),
.B1(n_6514),
.B2(n_6523),
.Y(n_8829)
);

AND2x2_ASAP7_75t_L g8830 ( 
.A(n_6958),
.B(n_8074),
.Y(n_8830)
);

AOI22x1_ASAP7_75t_L g8831 ( 
.A1(n_8031),
.A2(n_6398),
.B1(n_6453),
.B2(n_6300),
.Y(n_8831)
);

O2A1O1Ixp33_ASAP7_75t_L g8832 ( 
.A1(n_7011),
.A2(n_6540),
.B(n_6671),
.C(n_6662),
.Y(n_8832)
);

A2O1A1Ixp33_ASAP7_75t_SL g8833 ( 
.A1(n_7595),
.A2(n_6706),
.B(n_6790),
.C(n_6704),
.Y(n_8833)
);

CKINVDCx5p33_ASAP7_75t_R g8834 ( 
.A(n_7729),
.Y(n_8834)
);

BUFx6f_ASAP7_75t_L g8835 ( 
.A(n_6926),
.Y(n_8835)
);

BUFx3_ASAP7_75t_L g8836 ( 
.A(n_7177),
.Y(n_8836)
);

BUFx6f_ASAP7_75t_L g8837 ( 
.A(n_6926),
.Y(n_8837)
);

OAI221xp5_ASAP7_75t_L g8838 ( 
.A1(n_7250),
.A2(n_7261),
.B1(n_7175),
.B2(n_7170),
.C(n_7318),
.Y(n_8838)
);

OAI21x1_ASAP7_75t_L g8839 ( 
.A1(n_7408),
.A2(n_7455),
.B(n_7415),
.Y(n_8839)
);

INVx1_ASAP7_75t_L g8840 ( 
.A(n_7246),
.Y(n_8840)
);

AOI21xp5_ASAP7_75t_L g8841 ( 
.A1(n_7914),
.A2(n_6361),
.B(n_6335),
.Y(n_8841)
);

INVx2_ASAP7_75t_L g8842 ( 
.A(n_7159),
.Y(n_8842)
);

AND2x2_ASAP7_75t_L g8843 ( 
.A(n_6958),
.B(n_6297),
.Y(n_8843)
);

INVx8_ASAP7_75t_L g8844 ( 
.A(n_7138),
.Y(n_8844)
);

BUFx8_ASAP7_75t_SL g8845 ( 
.A(n_7045),
.Y(n_8845)
);

OAI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_7849),
.A2(n_7175),
.B1(n_7822),
.B2(n_7802),
.Y(n_8846)
);

AOI21xp5_ASAP7_75t_L g8847 ( 
.A1(n_8047),
.A2(n_6361),
.B(n_6335),
.Y(n_8847)
);

BUFx3_ASAP7_75t_L g8848 ( 
.A(n_7177),
.Y(n_8848)
);

AOI21xp5_ASAP7_75t_L g8849 ( 
.A1(n_8047),
.A2(n_7964),
.B(n_7912),
.Y(n_8849)
);

OAI21xp5_ASAP7_75t_L g8850 ( 
.A1(n_7420),
.A2(n_6809),
.B(n_6800),
.Y(n_8850)
);

INVx4_ASAP7_75t_L g8851 ( 
.A(n_7166),
.Y(n_8851)
);

INVx1_ASAP7_75t_L g8852 ( 
.A(n_7290),
.Y(n_8852)
);

BUFx2_ASAP7_75t_L g8853 ( 
.A(n_6958),
.Y(n_8853)
);

HB1xp67_ASAP7_75t_L g8854 ( 
.A(n_7506),
.Y(n_8854)
);

NAND2xp5_ASAP7_75t_L g8855 ( 
.A(n_7006),
.B(n_6167),
.Y(n_8855)
);

OA21x2_ASAP7_75t_L g8856 ( 
.A1(n_7415),
.A2(n_6372),
.B(n_6362),
.Y(n_8856)
);

INVx2_ASAP7_75t_L g8857 ( 
.A(n_7159),
.Y(n_8857)
);

OAI21xp5_ASAP7_75t_L g8858 ( 
.A1(n_7613),
.A2(n_7872),
.B(n_7850),
.Y(n_8858)
);

A2O1A1Ixp33_ASAP7_75t_L g8859 ( 
.A1(n_7044),
.A2(n_6017),
.B(n_6251),
.C(n_6243),
.Y(n_8859)
);

OAI221xp5_ASAP7_75t_L g8860 ( 
.A1(n_7250),
.A2(n_5752),
.B1(n_5904),
.B2(n_5906),
.C(n_5899),
.Y(n_8860)
);

OR2x2_ASAP7_75t_L g8861 ( 
.A(n_7475),
.B(n_6167),
.Y(n_8861)
);

AOI22xp33_ASAP7_75t_SL g8862 ( 
.A1(n_7932),
.A2(n_6319),
.B1(n_6308),
.B2(n_6243),
.Y(n_8862)
);

INVx2_ASAP7_75t_L g8863 ( 
.A(n_7159),
.Y(n_8863)
);

NAND2xp5_ASAP7_75t_L g8864 ( 
.A(n_7006),
.B(n_7986),
.Y(n_8864)
);

O2A1O1Ixp33_ASAP7_75t_L g8865 ( 
.A1(n_7011),
.A2(n_6671),
.B(n_6662),
.C(n_6836),
.Y(n_8865)
);

BUFx3_ASAP7_75t_L g8866 ( 
.A(n_7177),
.Y(n_8866)
);

BUFx2_ASAP7_75t_L g8867 ( 
.A(n_6958),
.Y(n_8867)
);

INVx3_ASAP7_75t_L g8868 ( 
.A(n_7797),
.Y(n_8868)
);

AOI22xp33_ASAP7_75t_SL g8869 ( 
.A1(n_7978),
.A2(n_8050),
.B1(n_7328),
.B2(n_7171),
.Y(n_8869)
);

INVx3_ASAP7_75t_L g8870 ( 
.A(n_7797),
.Y(n_8870)
);

BUFx3_ASAP7_75t_L g8871 ( 
.A(n_7819),
.Y(n_8871)
);

OAI21xp5_ASAP7_75t_L g8872 ( 
.A1(n_7850),
.A2(n_6838),
.B(n_6836),
.Y(n_8872)
);

A2O1A1Ixp33_ASAP7_75t_L g8873 ( 
.A1(n_7137),
.A2(n_6017),
.B(n_6251),
.C(n_6243),
.Y(n_8873)
);

INVx2_ASAP7_75t_L g8874 ( 
.A(n_7159),
.Y(n_8874)
);

AND2x2_ASAP7_75t_L g8875 ( 
.A(n_6958),
.B(n_6297),
.Y(n_8875)
);

OR2x6_ASAP7_75t_L g8876 ( 
.A(n_8118),
.B(n_6332),
.Y(n_8876)
);

INVx2_ASAP7_75t_SL g8877 ( 
.A(n_7464),
.Y(n_8877)
);

CKINVDCx20_ASAP7_75t_R g8878 ( 
.A(n_7527),
.Y(n_8878)
);

BUFx8_ASAP7_75t_L g8879 ( 
.A(n_7166),
.Y(n_8879)
);

OAI21xp5_ASAP7_75t_L g8880 ( 
.A1(n_7872),
.A2(n_6846),
.B(n_6838),
.Y(n_8880)
);

INVx1_ASAP7_75t_SL g8881 ( 
.A(n_7001),
.Y(n_8881)
);

INVx1_ASAP7_75t_L g8882 ( 
.A(n_7290),
.Y(n_8882)
);

AOI21xp33_ASAP7_75t_SL g8883 ( 
.A1(n_7443),
.A2(n_6572),
.B(n_6476),
.Y(n_8883)
);

AND2x4_ASAP7_75t_L g8884 ( 
.A(n_7516),
.B(n_6216),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_7290),
.Y(n_8885)
);

AO31x2_ASAP7_75t_L g8886 ( 
.A1(n_7986),
.A2(n_8100),
.A3(n_8065),
.B(n_7328),
.Y(n_8886)
);

INVx1_ASAP7_75t_L g8887 ( 
.A(n_7297),
.Y(n_8887)
);

AO21x1_ASAP7_75t_L g8888 ( 
.A1(n_7774),
.A2(n_6377),
.B(n_6372),
.Y(n_8888)
);

NAND3xp33_ASAP7_75t_L g8889 ( 
.A(n_7597),
.B(n_6856),
.C(n_6846),
.Y(n_8889)
);

AND2x2_ASAP7_75t_L g8890 ( 
.A(n_8074),
.B(n_6297),
.Y(n_8890)
);

AND2x2_ASAP7_75t_L g8891 ( 
.A(n_8074),
.B(n_8089),
.Y(n_8891)
);

AOI21x1_ASAP7_75t_L g8892 ( 
.A1(n_7913),
.A2(n_5756),
.B(n_5744),
.Y(n_8892)
);

NAND2x1p5_ASAP7_75t_L g8893 ( 
.A(n_7636),
.B(n_6416),
.Y(n_8893)
);

INVx2_ASAP7_75t_L g8894 ( 
.A(n_7178),
.Y(n_8894)
);

INVx2_ASAP7_75t_SL g8895 ( 
.A(n_7516),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_7297),
.Y(n_8896)
);

AND2x4_ASAP7_75t_L g8897 ( 
.A(n_7516),
.B(n_6216),
.Y(n_8897)
);

INVx1_ASAP7_75t_L g8898 ( 
.A(n_7297),
.Y(n_8898)
);

INVx1_ASAP7_75t_L g8899 ( 
.A(n_7310),
.Y(n_8899)
);

NOR2xp67_ASAP7_75t_L g8900 ( 
.A(n_7154),
.B(n_6105),
.Y(n_8900)
);

OAI21xp5_ASAP7_75t_L g8901 ( 
.A1(n_7505),
.A2(n_6856),
.B(n_5842),
.Y(n_8901)
);

INVx2_ASAP7_75t_L g8902 ( 
.A(n_7178),
.Y(n_8902)
);

AOI21xp5_ASAP7_75t_L g8903 ( 
.A1(n_7912),
.A2(n_6361),
.B(n_6335),
.Y(n_8903)
);

INVx4_ASAP7_75t_L g8904 ( 
.A(n_7166),
.Y(n_8904)
);

AO21x2_ASAP7_75t_L g8905 ( 
.A1(n_6984),
.A2(n_5429),
.B(n_5422),
.Y(n_8905)
);

BUFx2_ASAP7_75t_L g8906 ( 
.A(n_7964),
.Y(n_8906)
);

OAI21xp5_ASAP7_75t_L g8907 ( 
.A1(n_7505),
.A2(n_5849),
.B(n_5835),
.Y(n_8907)
);

NAND2xp5_ASAP7_75t_L g8908 ( 
.A(n_7986),
.B(n_6180),
.Y(n_8908)
);

O2A1O1Ixp33_ASAP7_75t_L g8909 ( 
.A1(n_7603),
.A2(n_5771),
.B(n_5815),
.C(n_5749),
.Y(n_8909)
);

INVx2_ASAP7_75t_SL g8910 ( 
.A(n_7516),
.Y(n_8910)
);

OAI21x1_ASAP7_75t_L g8911 ( 
.A1(n_7474),
.A2(n_7487),
.B(n_7484),
.Y(n_8911)
);

INVxp67_ASAP7_75t_SL g8912 ( 
.A(n_7683),
.Y(n_8912)
);

OAI22xp5_ASAP7_75t_L g8913 ( 
.A1(n_7849),
.A2(n_6095),
.B1(n_6144),
.B2(n_6009),
.Y(n_8913)
);

AO21x2_ASAP7_75t_L g8914 ( 
.A1(n_8096),
.A2(n_5429),
.B(n_5422),
.Y(n_8914)
);

INVx1_ASAP7_75t_L g8915 ( 
.A(n_7310),
.Y(n_8915)
);

AO21x2_ASAP7_75t_L g8916 ( 
.A1(n_8096),
.A2(n_5429),
.B(n_5422),
.Y(n_8916)
);

AO21x1_ASAP7_75t_L g8917 ( 
.A1(n_7407),
.A2(n_6391),
.B(n_6377),
.Y(n_8917)
);

OAI22xp5_ASAP7_75t_L g8918 ( 
.A1(n_7802),
.A2(n_6095),
.B1(n_6144),
.B2(n_6009),
.Y(n_8918)
);

INVx2_ASAP7_75t_L g8919 ( 
.A(n_7178),
.Y(n_8919)
);

INVx1_ASAP7_75t_SL g8920 ( 
.A(n_7023),
.Y(n_8920)
);

AND2x4_ASAP7_75t_L g8921 ( 
.A(n_7526),
.B(n_6216),
.Y(n_8921)
);

AND2x4_ASAP7_75t_L g8922 ( 
.A(n_7526),
.B(n_6216),
.Y(n_8922)
);

CKINVDCx5p33_ASAP7_75t_R g8923 ( 
.A(n_7868),
.Y(n_8923)
);

NOR2xp33_ASAP7_75t_SL g8924 ( 
.A(n_7413),
.B(n_6020),
.Y(n_8924)
);

BUFx12f_ASAP7_75t_L g8925 ( 
.A(n_6951),
.Y(n_8925)
);

OAI21xp5_ASAP7_75t_L g8926 ( 
.A1(n_7505),
.A2(n_5867),
.B(n_5864),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_7310),
.Y(n_8927)
);

INVx1_ASAP7_75t_L g8928 ( 
.A(n_7321),
.Y(n_8928)
);

OA21x2_ASAP7_75t_L g8929 ( 
.A1(n_7484),
.A2(n_6399),
.B(n_6391),
.Y(n_8929)
);

OAI22xp5_ASAP7_75t_L g8930 ( 
.A1(n_7802),
.A2(n_6164),
.B1(n_6242),
.B2(n_6196),
.Y(n_8930)
);

NAND2xp5_ASAP7_75t_L g8931 ( 
.A(n_7037),
.B(n_7026),
.Y(n_8931)
);

AO21x2_ASAP7_75t_L g8932 ( 
.A1(n_8096),
.A2(n_7719),
.B(n_7895),
.Y(n_8932)
);

AO31x2_ASAP7_75t_L g8933 ( 
.A1(n_8100),
.A2(n_6414),
.A3(n_6415),
.B(n_6399),
.Y(n_8933)
);

AOI22xp33_ASAP7_75t_SL g8934 ( 
.A1(n_7978),
.A2(n_6319),
.B1(n_6308),
.B2(n_6268),
.Y(n_8934)
);

AOI22xp5_ASAP7_75t_L g8935 ( 
.A1(n_7713),
.A2(n_6565),
.B1(n_6514),
.B2(n_6523),
.Y(n_8935)
);

AOI22xp33_ASAP7_75t_L g8936 ( 
.A1(n_7261),
.A2(n_6170),
.B1(n_6191),
.B2(n_6105),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_7321),
.Y(n_8937)
);

HB1xp67_ASAP7_75t_L g8938 ( 
.A(n_7506),
.Y(n_8938)
);

OAI222xp33_ASAP7_75t_L g8939 ( 
.A1(n_8013),
.A2(n_6332),
.B1(n_6020),
.B2(n_6361),
.C1(n_6393),
.C2(n_6335),
.Y(n_8939)
);

OAI21x1_ASAP7_75t_L g8940 ( 
.A1(n_7498),
.A2(n_7510),
.B(n_7503),
.Y(n_8940)
);

INVx1_ASAP7_75t_L g8941 ( 
.A(n_7321),
.Y(n_8941)
);

OAI21xp5_ASAP7_75t_L g8942 ( 
.A1(n_7597),
.A2(n_5867),
.B(n_5864),
.Y(n_8942)
);

BUFx6f_ASAP7_75t_L g8943 ( 
.A(n_6926),
.Y(n_8943)
);

AOI21xp5_ASAP7_75t_L g8944 ( 
.A1(n_8022),
.A2(n_6361),
.B(n_6335),
.Y(n_8944)
);

OA21x2_ASAP7_75t_L g8945 ( 
.A1(n_7498),
.A2(n_7510),
.B(n_7503),
.Y(n_8945)
);

INVx2_ASAP7_75t_L g8946 ( 
.A(n_7178),
.Y(n_8946)
);

CKINVDCx8_ASAP7_75t_R g8947 ( 
.A(n_6951),
.Y(n_8947)
);

OAI21x1_ASAP7_75t_L g8948 ( 
.A1(n_7498),
.A2(n_7510),
.B(n_7503),
.Y(n_8948)
);

INVx2_ASAP7_75t_SL g8949 ( 
.A(n_7526),
.Y(n_8949)
);

INVx1_ASAP7_75t_L g8950 ( 
.A(n_7322),
.Y(n_8950)
);

BUFx6f_ASAP7_75t_L g8951 ( 
.A(n_6926),
.Y(n_8951)
);

AND2x2_ASAP7_75t_L g8952 ( 
.A(n_8074),
.B(n_6299),
.Y(n_8952)
);

INVx1_ASAP7_75t_L g8953 ( 
.A(n_7322),
.Y(n_8953)
);

AND2x6_ASAP7_75t_L g8954 ( 
.A(n_7795),
.B(n_6002),
.Y(n_8954)
);

INVx5_ASAP7_75t_L g8955 ( 
.A(n_7819),
.Y(n_8955)
);

XNOR2xp5_ASAP7_75t_L g8956 ( 
.A(n_7527),
.B(n_5896),
.Y(n_8956)
);

AOI22xp33_ASAP7_75t_L g8957 ( 
.A1(n_7603),
.A2(n_7760),
.B1(n_7318),
.B2(n_7319),
.Y(n_8957)
);

INVx1_ASAP7_75t_L g8958 ( 
.A(n_7322),
.Y(n_8958)
);

NOR2xp33_ASAP7_75t_L g8959 ( 
.A(n_7100),
.B(n_6849),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_7333),
.Y(n_8960)
);

INVx2_ASAP7_75t_L g8961 ( 
.A(n_7186),
.Y(n_8961)
);

OR2x6_ASAP7_75t_L g8962 ( 
.A(n_8118),
.B(n_6332),
.Y(n_8962)
);

INVx2_ASAP7_75t_L g8963 ( 
.A(n_7186),
.Y(n_8963)
);

OAI22xp5_ASAP7_75t_SL g8964 ( 
.A1(n_7289),
.A2(n_6128),
.B1(n_6653),
.B2(n_6227),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_7333),
.Y(n_8965)
);

AO31x2_ASAP7_75t_L g8966 ( 
.A1(n_8100),
.A2(n_6415),
.A3(n_6418),
.B(n_6414),
.Y(n_8966)
);

AOI21x1_ASAP7_75t_L g8967 ( 
.A1(n_7913),
.A2(n_6433),
.B(n_6182),
.Y(n_8967)
);

CKINVDCx6p67_ASAP7_75t_R g8968 ( 
.A(n_7166),
.Y(n_8968)
);

BUFx6f_ASAP7_75t_L g8969 ( 
.A(n_6926),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_7333),
.Y(n_8970)
);

NAND3xp33_ASAP7_75t_L g8971 ( 
.A(n_7597),
.B(n_6182),
.C(n_6180),
.Y(n_8971)
);

AND2x2_ASAP7_75t_L g8972 ( 
.A(n_8089),
.B(n_6299),
.Y(n_8972)
);

INVx2_ASAP7_75t_L g8973 ( 
.A(n_7186),
.Y(n_8973)
);

OAI22xp5_ASAP7_75t_L g8974 ( 
.A1(n_7822),
.A2(n_6196),
.B1(n_6242),
.B2(n_6164),
.Y(n_8974)
);

AND2x4_ASAP7_75t_L g8975 ( 
.A(n_7526),
.B(n_6226),
.Y(n_8975)
);

INVx2_ASAP7_75t_L g8976 ( 
.A(n_7186),
.Y(n_8976)
);

AND2x4_ASAP7_75t_L g8977 ( 
.A(n_7579),
.B(n_6226),
.Y(n_8977)
);

BUFx2_ASAP7_75t_L g8978 ( 
.A(n_7160),
.Y(n_8978)
);

AND2x2_ASAP7_75t_L g8979 ( 
.A(n_8089),
.B(n_6299),
.Y(n_8979)
);

OAI21xp5_ASAP7_75t_L g8980 ( 
.A1(n_7864),
.A2(n_5771),
.B(n_5749),
.Y(n_8980)
);

AOI22xp33_ASAP7_75t_L g8981 ( 
.A1(n_7760),
.A2(n_6191),
.B1(n_6227),
.B2(n_6170),
.Y(n_8981)
);

NAND2x1p5_ASAP7_75t_L g8982 ( 
.A(n_7636),
.B(n_6435),
.Y(n_8982)
);

INVx3_ASAP7_75t_L g8983 ( 
.A(n_7797),
.Y(n_8983)
);

OA21x2_ASAP7_75t_L g8984 ( 
.A1(n_7633),
.A2(n_6441),
.B(n_6418),
.Y(n_8984)
);

AO21x2_ASAP7_75t_L g8985 ( 
.A1(n_7895),
.A2(n_5429),
.B(n_5422),
.Y(n_8985)
);

AO21x2_ASAP7_75t_L g8986 ( 
.A1(n_7895),
.A2(n_5441),
.B(n_5432),
.Y(n_8986)
);

NAND3xp33_ASAP7_75t_L g8987 ( 
.A(n_7864),
.B(n_6198),
.C(n_6185),
.Y(n_8987)
);

OA21x2_ASAP7_75t_L g8988 ( 
.A1(n_7635),
.A2(n_6447),
.B(n_6441),
.Y(n_8988)
);

INVx1_ASAP7_75t_L g8989 ( 
.A(n_7338),
.Y(n_8989)
);

INVx2_ASAP7_75t_L g8990 ( 
.A(n_7190),
.Y(n_8990)
);

AO21x2_ASAP7_75t_L g8991 ( 
.A1(n_8020),
.A2(n_5441),
.B(n_5432),
.Y(n_8991)
);

BUFx2_ASAP7_75t_L g8992 ( 
.A(n_7160),
.Y(n_8992)
);

AOI21xp33_ASAP7_75t_L g8993 ( 
.A1(n_7785),
.A2(n_6448),
.B(n_6447),
.Y(n_8993)
);

A2O1A1Ixp33_ASAP7_75t_L g8994 ( 
.A1(n_7137),
.A2(n_6268),
.B(n_6285),
.C(n_6251),
.Y(n_8994)
);

OAI21x1_ASAP7_75t_SL g8995 ( 
.A1(n_7109),
.A2(n_6151),
.B(n_6075),
.Y(n_8995)
);

AOI222xp33_ASAP7_75t_L g8996 ( 
.A1(n_7070),
.A2(n_5899),
.B1(n_5904),
.B2(n_5906),
.C1(n_6681),
.C2(n_6664),
.Y(n_8996)
);

AND2x6_ASAP7_75t_L g8997 ( 
.A(n_7795),
.B(n_6002),
.Y(n_8997)
);

OAI21xp5_ASAP7_75t_L g8998 ( 
.A1(n_7864),
.A2(n_5905),
.B(n_5815),
.Y(n_8998)
);

INVx3_ASAP7_75t_L g8999 ( 
.A(n_7797),
.Y(n_8999)
);

AOI22xp5_ASAP7_75t_L g9000 ( 
.A1(n_8085),
.A2(n_6483),
.B1(n_5998),
.B2(n_6030),
.Y(n_9000)
);

NAND2x1p5_ASAP7_75t_L g9001 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9001)
);

OAI21xp5_ASAP7_75t_L g9002 ( 
.A1(n_7768),
.A2(n_5905),
.B(n_6185),
.Y(n_9002)
);

O2A1O1Ixp33_ASAP7_75t_SL g9003 ( 
.A1(n_7929),
.A2(n_6486),
.B(n_6490),
.C(n_6802),
.Y(n_9003)
);

BUFx10_ASAP7_75t_L g9004 ( 
.A(n_7485),
.Y(n_9004)
);

AO21x2_ASAP7_75t_L g9005 ( 
.A1(n_8020),
.A2(n_5441),
.B(n_5432),
.Y(n_9005)
);

NAND3xp33_ASAP7_75t_L g9006 ( 
.A(n_7169),
.B(n_6199),
.C(n_6198),
.Y(n_9006)
);

INVx1_ASAP7_75t_L g9007 ( 
.A(n_7338),
.Y(n_9007)
);

OAI21xp5_ASAP7_75t_L g9008 ( 
.A1(n_7768),
.A2(n_6199),
.B(n_6448),
.Y(n_9008)
);

INVx3_ASAP7_75t_L g9009 ( 
.A(n_7797),
.Y(n_9009)
);

INVx1_ASAP7_75t_SL g9010 ( 
.A(n_7023),
.Y(n_9010)
);

INVx3_ASAP7_75t_L g9011 ( 
.A(n_7809),
.Y(n_9011)
);

BUFx2_ASAP7_75t_L g9012 ( 
.A(n_7160),
.Y(n_9012)
);

OAI22xp5_ASAP7_75t_L g9013 ( 
.A1(n_7822),
.A2(n_6164),
.B1(n_6242),
.B2(n_6196),
.Y(n_9013)
);

INVx2_ASAP7_75t_L g9014 ( 
.A(n_7190),
.Y(n_9014)
);

AO21x2_ASAP7_75t_L g9015 ( 
.A1(n_8020),
.A2(n_5441),
.B(n_5432),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_7338),
.Y(n_9016)
);

OAI21xp5_ASAP7_75t_L g9017 ( 
.A1(n_7768),
.A2(n_6460),
.B(n_6451),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_7357),
.Y(n_9018)
);

NAND2xp5_ASAP7_75t_L g9019 ( 
.A(n_7037),
.B(n_6849),
.Y(n_9019)
);

INVx2_ASAP7_75t_SL g9020 ( 
.A(n_7579),
.Y(n_9020)
);

CKINVDCx5p33_ASAP7_75t_R g9021 ( 
.A(n_7868),
.Y(n_9021)
);

OR2x2_ASAP7_75t_L g9022 ( 
.A(n_7390),
.B(n_6850),
.Y(n_9022)
);

OAI21xp5_ASAP7_75t_L g9023 ( 
.A1(n_7770),
.A2(n_6460),
.B(n_6451),
.Y(n_9023)
);

NOR3xp33_ASAP7_75t_L g9024 ( 
.A(n_7808),
.B(n_5827),
.C(n_5819),
.Y(n_9024)
);

AOI22xp33_ASAP7_75t_L g9025 ( 
.A1(n_7319),
.A2(n_6191),
.B1(n_6227),
.B2(n_6170),
.Y(n_9025)
);

OAI21x1_ASAP7_75t_L g9026 ( 
.A1(n_7641),
.A2(n_6903),
.B(n_6858),
.Y(n_9026)
);

NAND2xp5_ASAP7_75t_L g9027 ( 
.A(n_7037),
.B(n_6850),
.Y(n_9027)
);

INVx1_ASAP7_75t_L g9028 ( 
.A(n_7357),
.Y(n_9028)
);

INVx2_ASAP7_75t_L g9029 ( 
.A(n_7190),
.Y(n_9029)
);

OAI21xp5_ASAP7_75t_L g9030 ( 
.A1(n_7770),
.A2(n_6462),
.B(n_6461),
.Y(n_9030)
);

BUFx6f_ASAP7_75t_L g9031 ( 
.A(n_6949),
.Y(n_9031)
);

NAND2x1p5_ASAP7_75t_L g9032 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_7357),
.Y(n_9033)
);

INVx1_ASAP7_75t_SL g9034 ( 
.A(n_7054),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_SL g9035 ( 
.A(n_8050),
.B(n_6226),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_L g9036 ( 
.A(n_7026),
.B(n_6461),
.Y(n_9036)
);

OAI22xp5_ASAP7_75t_L g9037 ( 
.A1(n_8084),
.A2(n_6314),
.B1(n_6324),
.B2(n_6254),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_7359),
.Y(n_9038)
);

OAI21xp5_ASAP7_75t_L g9039 ( 
.A1(n_7770),
.A2(n_6463),
.B(n_6462),
.Y(n_9039)
);

INVx8_ASAP7_75t_L g9040 ( 
.A(n_7214),
.Y(n_9040)
);

OAI22xp5_ASAP7_75t_SL g9041 ( 
.A1(n_7289),
.A2(n_6653),
.B1(n_6128),
.B2(n_6191),
.Y(n_9041)
);

NAND2xp5_ASAP7_75t_L g9042 ( 
.A(n_7026),
.B(n_7030),
.Y(n_9042)
);

CKINVDCx5p33_ASAP7_75t_R g9043 ( 
.A(n_6956),
.Y(n_9043)
);

HB1xp67_ASAP7_75t_L g9044 ( 
.A(n_7507),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_7359),
.Y(n_9045)
);

OAI21x1_ASAP7_75t_L g9046 ( 
.A1(n_7672),
.A2(n_6903),
.B(n_6858),
.Y(n_9046)
);

OAI21x1_ASAP7_75t_L g9047 ( 
.A1(n_7672),
.A2(n_6903),
.B(n_6759),
.Y(n_9047)
);

OA21x2_ASAP7_75t_L g9048 ( 
.A1(n_7672),
.A2(n_6470),
.B(n_6463),
.Y(n_9048)
);

CKINVDCx5p33_ASAP7_75t_R g9049 ( 
.A(n_6956),
.Y(n_9049)
);

OAI21x1_ASAP7_75t_L g9050 ( 
.A1(n_7673),
.A2(n_6759),
.B(n_6719),
.Y(n_9050)
);

INVx1_ASAP7_75t_L g9051 ( 
.A(n_7359),
.Y(n_9051)
);

NAND2xp5_ASAP7_75t_L g9052 ( 
.A(n_7030),
.B(n_6470),
.Y(n_9052)
);

OAI21x1_ASAP7_75t_L g9053 ( 
.A1(n_7673),
.A2(n_6760),
.B(n_6719),
.Y(n_9053)
);

BUFx6f_ASAP7_75t_L g9054 ( 
.A(n_6949),
.Y(n_9054)
);

BUFx3_ASAP7_75t_L g9055 ( 
.A(n_7819),
.Y(n_9055)
);

AND2x2_ASAP7_75t_SL g9056 ( 
.A(n_7171),
.B(n_6226),
.Y(n_9056)
);

OAI22xp33_ASAP7_75t_L g9057 ( 
.A1(n_8084),
.A2(n_6268),
.B1(n_6285),
.B2(n_6251),
.Y(n_9057)
);

AO31x2_ASAP7_75t_L g9058 ( 
.A1(n_8065),
.A2(n_6496),
.A3(n_6499),
.B(n_6495),
.Y(n_9058)
);

AOI222xp33_ASAP7_75t_L g9059 ( 
.A1(n_7070),
.A2(n_8043),
.B1(n_7902),
.B2(n_7390),
.C1(n_8013),
.C2(n_7991),
.Y(n_9059)
);

INVx4_ASAP7_75t_L g9060 ( 
.A(n_7214),
.Y(n_9060)
);

NAND2xp5_ASAP7_75t_L g9061 ( 
.A(n_7030),
.B(n_6495),
.Y(n_9061)
);

OAI21x1_ASAP7_75t_L g9062 ( 
.A1(n_7673),
.A2(n_7193),
.B(n_7191),
.Y(n_9062)
);

OAI21x1_ASAP7_75t_L g9063 ( 
.A1(n_7191),
.A2(n_6786),
.B(n_6760),
.Y(n_9063)
);

NAND2x1p5_ASAP7_75t_L g9064 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9064)
);

INVx3_ASAP7_75t_L g9065 ( 
.A(n_7809),
.Y(n_9065)
);

OAI21x1_ASAP7_75t_L g9066 ( 
.A1(n_7191),
.A2(n_6841),
.B(n_6786),
.Y(n_9066)
);

OAI21x1_ASAP7_75t_L g9067 ( 
.A1(n_7193),
.A2(n_6865),
.B(n_6841),
.Y(n_9067)
);

OAI21x1_ASAP7_75t_L g9068 ( 
.A1(n_7193),
.A2(n_6885),
.B(n_6865),
.Y(n_9068)
);

OAI21xp5_ASAP7_75t_L g9069 ( 
.A1(n_7786),
.A2(n_6516),
.B(n_6496),
.Y(n_9069)
);

OA21x2_ASAP7_75t_L g9070 ( 
.A1(n_7885),
.A2(n_6521),
.B(n_6519),
.Y(n_9070)
);

CKINVDCx11_ASAP7_75t_R g9071 ( 
.A(n_7054),
.Y(n_9071)
);

AO31x2_ASAP7_75t_L g9072 ( 
.A1(n_8065),
.A2(n_6521),
.A3(n_6537),
.B(n_6519),
.Y(n_9072)
);

OAI22xp33_ASAP7_75t_L g9073 ( 
.A1(n_8084),
.A2(n_6285),
.B1(n_6268),
.B2(n_6308),
.Y(n_9073)
);

OAI21x1_ASAP7_75t_L g9074 ( 
.A1(n_7721),
.A2(n_6885),
.B(n_6483),
.Y(n_9074)
);

NOR2xp33_ASAP7_75t_L g9075 ( 
.A(n_7253),
.B(n_6917),
.Y(n_9075)
);

OAI22xp5_ASAP7_75t_L g9076 ( 
.A1(n_8092),
.A2(n_6314),
.B1(n_6324),
.B2(n_6254),
.Y(n_9076)
);

OAI21x1_ASAP7_75t_L g9077 ( 
.A1(n_7721),
.A2(n_7738),
.B(n_7885),
.Y(n_9077)
);

INVx1_ASAP7_75t_L g9078 ( 
.A(n_7365),
.Y(n_9078)
);

AO31x2_ASAP7_75t_L g9079 ( 
.A1(n_7328),
.A2(n_6538),
.A3(n_6541),
.B(n_6537),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_7365),
.Y(n_9080)
);

OAI22xp5_ASAP7_75t_L g9081 ( 
.A1(n_8092),
.A2(n_6314),
.B1(n_6324),
.B2(n_6254),
.Y(n_9081)
);

NOR2xp33_ASAP7_75t_L g9082 ( 
.A(n_7253),
.B(n_6538),
.Y(n_9082)
);

INVx1_ASAP7_75t_L g9083 ( 
.A(n_7365),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_7386),
.Y(n_9084)
);

INVx2_ASAP7_75t_SL g9085 ( 
.A(n_7579),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_7386),
.Y(n_9086)
);

OA21x2_ASAP7_75t_L g9087 ( 
.A1(n_7885),
.A2(n_6552),
.B(n_6541),
.Y(n_9087)
);

AND2x2_ASAP7_75t_L g9088 ( 
.A(n_8089),
.B(n_6321),
.Y(n_9088)
);

AND2x4_ASAP7_75t_L g9089 ( 
.A(n_7579),
.B(n_6226),
.Y(n_9089)
);

AOI21xp5_ASAP7_75t_SL g9090 ( 
.A1(n_7763),
.A2(n_6490),
.B(n_6486),
.Y(n_9090)
);

NAND2xp5_ASAP7_75t_L g9091 ( 
.A(n_7094),
.B(n_6552),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_7386),
.Y(n_9092)
);

AOI21x1_ASAP7_75t_L g9093 ( 
.A1(n_7925),
.A2(n_6917),
.B(n_6595),
.Y(n_9093)
);

INVx1_ASAP7_75t_L g9094 ( 
.A(n_7399),
.Y(n_9094)
);

OAI21x1_ASAP7_75t_L g9095 ( 
.A1(n_7721),
.A2(n_6595),
.B(n_6567),
.Y(n_9095)
);

INVx2_ASAP7_75t_L g9096 ( 
.A(n_7190),
.Y(n_9096)
);

AND2x2_ASAP7_75t_L g9097 ( 
.A(n_8099),
.B(n_6321),
.Y(n_9097)
);

OAI22xp33_ASAP7_75t_L g9098 ( 
.A1(n_8092),
.A2(n_6285),
.B1(n_6319),
.B2(n_6308),
.Y(n_9098)
);

OAI21x1_ASAP7_75t_L g9099 ( 
.A1(n_7738),
.A2(n_7896),
.B(n_7893),
.Y(n_9099)
);

OAI21xp5_ASAP7_75t_L g9100 ( 
.A1(n_7786),
.A2(n_6617),
.B(n_6567),
.Y(n_9100)
);

INVx1_ASAP7_75t_L g9101 ( 
.A(n_7399),
.Y(n_9101)
);

OAI21x1_ASAP7_75t_L g9102 ( 
.A1(n_7738),
.A2(n_6625),
.B(n_6617),
.Y(n_9102)
);

NAND2x1p5_ASAP7_75t_L g9103 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9103)
);

OR2x2_ASAP7_75t_L g9104 ( 
.A(n_7094),
.B(n_6333),
.Y(n_9104)
);

OAI21x1_ASAP7_75t_L g9105 ( 
.A1(n_7893),
.A2(n_6631),
.B(n_6625),
.Y(n_9105)
);

INVx2_ASAP7_75t_L g9106 ( 
.A(n_7198),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_7399),
.Y(n_9107)
);

OAI21x1_ASAP7_75t_L g9108 ( 
.A1(n_7893),
.A2(n_6650),
.B(n_6631),
.Y(n_9108)
);

AOI21xp5_ASAP7_75t_L g9109 ( 
.A1(n_8022),
.A2(n_6393),
.B(n_6361),
.Y(n_9109)
);

BUFx2_ASAP7_75t_R g9110 ( 
.A(n_7350),
.Y(n_9110)
);

CKINVDCx6p67_ASAP7_75t_R g9111 ( 
.A(n_7214),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_7406),
.Y(n_9112)
);

OAI21x1_ASAP7_75t_L g9113 ( 
.A1(n_7896),
.A2(n_6655),
.B(n_6650),
.Y(n_9113)
);

INVx1_ASAP7_75t_L g9114 ( 
.A(n_7406),
.Y(n_9114)
);

BUFx2_ASAP7_75t_L g9115 ( 
.A(n_7162),
.Y(n_9115)
);

INVx2_ASAP7_75t_L g9116 ( 
.A(n_7198),
.Y(n_9116)
);

NAND3xp33_ASAP7_75t_L g9117 ( 
.A(n_7169),
.B(n_6673),
.C(n_6655),
.Y(n_9117)
);

NOR2xp33_ASAP7_75t_L g9118 ( 
.A(n_7902),
.B(n_6673),
.Y(n_9118)
);

INVx1_ASAP7_75t_L g9119 ( 
.A(n_7406),
.Y(n_9119)
);

OAI21x1_ASAP7_75t_L g9120 ( 
.A1(n_7896),
.A2(n_6690),
.B(n_6687),
.Y(n_9120)
);

A2O1A1Ixp33_ASAP7_75t_L g9121 ( 
.A1(n_7137),
.A2(n_6170),
.B(n_6227),
.C(n_6191),
.Y(n_9121)
);

INVx1_ASAP7_75t_L g9122 ( 
.A(n_7430),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_7198),
.Y(n_9123)
);

OAI21x1_ASAP7_75t_L g9124 ( 
.A1(n_7573),
.A2(n_6690),
.B(n_6687),
.Y(n_9124)
);

OA21x2_ASAP7_75t_L g9125 ( 
.A1(n_8029),
.A2(n_6703),
.B(n_6697),
.Y(n_9125)
);

NAND2x1p5_ASAP7_75t_L g9126 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9126)
);

AOI22xp33_ASAP7_75t_L g9127 ( 
.A1(n_7426),
.A2(n_6191),
.B1(n_6227),
.B2(n_6170),
.Y(n_9127)
);

OAI21x1_ASAP7_75t_L g9128 ( 
.A1(n_7573),
.A2(n_6703),
.B(n_6697),
.Y(n_9128)
);

INVx1_ASAP7_75t_L g9129 ( 
.A(n_7430),
.Y(n_9129)
);

OAI21x1_ASAP7_75t_L g9130 ( 
.A1(n_7573),
.A2(n_6727),
.B(n_6716),
.Y(n_9130)
);

AO21x2_ASAP7_75t_L g9131 ( 
.A1(n_7427),
.A2(n_5662),
.B(n_5659),
.Y(n_9131)
);

A2O1A1Ixp33_ASAP7_75t_L g9132 ( 
.A1(n_6925),
.A2(n_6191),
.B(n_6272),
.C(n_6227),
.Y(n_9132)
);

OAI21x1_ASAP7_75t_L g9133 ( 
.A1(n_7708),
.A2(n_6727),
.B(n_6716),
.Y(n_9133)
);

OAI22xp5_ASAP7_75t_L g9134 ( 
.A1(n_7090),
.A2(n_6333),
.B1(n_6345),
.B2(n_6339),
.Y(n_9134)
);

AO21x2_ASAP7_75t_L g9135 ( 
.A1(n_7427),
.A2(n_5662),
.B(n_5659),
.Y(n_9135)
);

AO31x2_ASAP7_75t_L g9136 ( 
.A1(n_7972),
.A2(n_6751),
.A3(n_6776),
.B(n_6740),
.Y(n_9136)
);

INVx2_ASAP7_75t_SL g9137 ( 
.A(n_7682),
.Y(n_9137)
);

NAND2x1p5_ASAP7_75t_L g9138 ( 
.A(n_7066),
.B(n_6435),
.Y(n_9138)
);

OAI21xp5_ASAP7_75t_L g9139 ( 
.A1(n_7786),
.A2(n_6751),
.B(n_6740),
.Y(n_9139)
);

NAND2xp5_ASAP7_75t_L g9140 ( 
.A(n_7094),
.B(n_6776),
.Y(n_9140)
);

BUFx4f_ASAP7_75t_L g9141 ( 
.A(n_7580),
.Y(n_9141)
);

CKINVDCx11_ASAP7_75t_R g9142 ( 
.A(n_7139),
.Y(n_9142)
);

HB1xp67_ASAP7_75t_L g9143 ( 
.A(n_7507),
.Y(n_9143)
);

INVx4_ASAP7_75t_SL g9144 ( 
.A(n_7393),
.Y(n_9144)
);

INVx2_ASAP7_75t_L g9145 ( 
.A(n_7198),
.Y(n_9145)
);

OR2x6_ASAP7_75t_L g9146 ( 
.A(n_8118),
.B(n_6361),
.Y(n_9146)
);

NAND2x1p5_ASAP7_75t_L g9147 ( 
.A(n_7144),
.B(n_6435),
.Y(n_9147)
);

CKINVDCx5p33_ASAP7_75t_R g9148 ( 
.A(n_7666),
.Y(n_9148)
);

OAI21x1_ASAP7_75t_SL g9149 ( 
.A1(n_7109),
.A2(n_6253),
.B(n_6172),
.Y(n_9149)
);

OAI21x1_ASAP7_75t_L g9150 ( 
.A1(n_7708),
.A2(n_6792),
.B(n_6784),
.Y(n_9150)
);

INVx2_ASAP7_75t_L g9151 ( 
.A(n_7201),
.Y(n_9151)
);

OAI21x1_ASAP7_75t_L g9152 ( 
.A1(n_7708),
.A2(n_6792),
.B(n_6784),
.Y(n_9152)
);

INVx1_ASAP7_75t_L g9153 ( 
.A(n_7430),
.Y(n_9153)
);

NAND2xp5_ASAP7_75t_L g9154 ( 
.A(n_7407),
.B(n_6797),
.Y(n_9154)
);

INVx2_ASAP7_75t_L g9155 ( 
.A(n_7201),
.Y(n_9155)
);

OAI21x1_ASAP7_75t_L g9156 ( 
.A1(n_7723),
.A2(n_6799),
.B(n_6797),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_7436),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_7436),
.Y(n_9158)
);

NOR3xp33_ASAP7_75t_L g9159 ( 
.A(n_7808),
.B(n_5827),
.C(n_5819),
.Y(n_9159)
);

HB1xp67_ASAP7_75t_L g9160 ( 
.A(n_7511),
.Y(n_9160)
);

OAI21x1_ASAP7_75t_L g9161 ( 
.A1(n_7723),
.A2(n_6811),
.B(n_6799),
.Y(n_9161)
);

OAI21x1_ASAP7_75t_L g9162 ( 
.A1(n_7723),
.A2(n_6817),
.B(n_6811),
.Y(n_9162)
);

INVx5_ASAP7_75t_L g9163 ( 
.A(n_7819),
.Y(n_9163)
);

NAND2xp5_ASAP7_75t_L g9164 ( 
.A(n_7407),
.B(n_6817),
.Y(n_9164)
);

AND2x4_ASAP7_75t_L g9165 ( 
.A(n_7682),
.B(n_7706),
.Y(n_9165)
);

AOI21xp5_ASAP7_75t_L g9166 ( 
.A1(n_6925),
.A2(n_7667),
.B(n_7655),
.Y(n_9166)
);

NAND3xp33_ASAP7_75t_L g9167 ( 
.A(n_7551),
.B(n_6828),
.C(n_6823),
.Y(n_9167)
);

INVx2_ASAP7_75t_L g9168 ( 
.A(n_7201),
.Y(n_9168)
);

INVx2_ASAP7_75t_SL g9169 ( 
.A(n_7682),
.Y(n_9169)
);

OAI21x1_ASAP7_75t_L g9170 ( 
.A1(n_7608),
.A2(n_6828),
.B(n_6823),
.Y(n_9170)
);

A2O1A1Ixp33_ASAP7_75t_L g9171 ( 
.A1(n_7089),
.A2(n_7780),
.B(n_7307),
.C(n_7991),
.Y(n_9171)
);

OAI21x1_ASAP7_75t_L g9172 ( 
.A1(n_7608),
.A2(n_6835),
.B(n_6832),
.Y(n_9172)
);

HB1xp67_ASAP7_75t_L g9173 ( 
.A(n_7511),
.Y(n_9173)
);

BUFx8_ASAP7_75t_L g9174 ( 
.A(n_7214),
.Y(n_9174)
);

OAI21x1_ASAP7_75t_L g9175 ( 
.A1(n_8029),
.A2(n_6835),
.B(n_6832),
.Y(n_9175)
);

OAI21x1_ASAP7_75t_L g9176 ( 
.A1(n_8029),
.A2(n_6861),
.B(n_6853),
.Y(n_9176)
);

AND2x2_ASAP7_75t_L g9177 ( 
.A(n_8099),
.B(n_8103),
.Y(n_9177)
);

INVx2_ASAP7_75t_L g9178 ( 
.A(n_7201),
.Y(n_9178)
);

OAI22xp5_ASAP7_75t_L g9179 ( 
.A1(n_7090),
.A2(n_6333),
.B1(n_6345),
.B2(n_6339),
.Y(n_9179)
);

AND2x2_ASAP7_75t_SL g9180 ( 
.A(n_7171),
.B(n_6002),
.Y(n_9180)
);

INVx1_ASAP7_75t_L g9181 ( 
.A(n_7436),
.Y(n_9181)
);

CKINVDCx5p33_ASAP7_75t_R g9182 ( 
.A(n_7666),
.Y(n_9182)
);

AOI22xp33_ASAP7_75t_L g9183 ( 
.A1(n_7426),
.A2(n_6272),
.B1(n_6227),
.B2(n_6393),
.Y(n_9183)
);

XNOR2xp5_ASAP7_75t_L g9184 ( 
.A(n_7531),
.B(n_5896),
.Y(n_9184)
);

AOI22xp33_ASAP7_75t_L g9185 ( 
.A1(n_7508),
.A2(n_6272),
.B1(n_6227),
.B2(n_6393),
.Y(n_9185)
);

BUFx3_ASAP7_75t_L g9186 ( 
.A(n_7819),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_L g9187 ( 
.A(n_7660),
.B(n_7675),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_7453),
.Y(n_9188)
);

INVx1_ASAP7_75t_L g9189 ( 
.A(n_7453),
.Y(n_9189)
);

BUFx2_ASAP7_75t_L g9190 ( 
.A(n_7162),
.Y(n_9190)
);

AND2x6_ASAP7_75t_L g9191 ( 
.A(n_7795),
.B(n_6002),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_7453),
.Y(n_9192)
);

BUFx2_ASAP7_75t_SL g9193 ( 
.A(n_7157),
.Y(n_9193)
);

AOI21xp5_ASAP7_75t_L g9194 ( 
.A1(n_7655),
.A2(n_6393),
.B(n_6587),
.Y(n_9194)
);

OAI21xp5_ASAP7_75t_L g9195 ( 
.A1(n_7439),
.A2(n_6861),
.B(n_6853),
.Y(n_9195)
);

BUFx6f_ASAP7_75t_L g9196 ( 
.A(n_6949),
.Y(n_9196)
);

BUFx6f_ASAP7_75t_L g9197 ( 
.A(n_6949),
.Y(n_9197)
);

AND2x2_ASAP7_75t_L g9198 ( 
.A(n_8099),
.B(n_6321),
.Y(n_9198)
);

AO21x2_ASAP7_75t_L g9199 ( 
.A1(n_7427),
.A2(n_5753),
.B(n_5730),
.Y(n_9199)
);

INVx2_ASAP7_75t_L g9200 ( 
.A(n_7220),
.Y(n_9200)
);

AOI22xp33_ASAP7_75t_L g9201 ( 
.A1(n_7508),
.A2(n_7664),
.B1(n_8085),
.B2(n_7204),
.Y(n_9201)
);

AOI21x1_ASAP7_75t_L g9202 ( 
.A1(n_7925),
.A2(n_7966),
.B(n_7935),
.Y(n_9202)
);

INVx1_ASAP7_75t_L g9203 ( 
.A(n_7454),
.Y(n_9203)
);

INVx1_ASAP7_75t_SL g9204 ( 
.A(n_7139),
.Y(n_9204)
);

AO31x2_ASAP7_75t_L g9205 ( 
.A1(n_7972),
.A2(n_6873),
.A3(n_6879),
.B(n_6869),
.Y(n_9205)
);

OAI21x1_ASAP7_75t_L g9206 ( 
.A1(n_8041),
.A2(n_6873),
.B(n_6869),
.Y(n_9206)
);

INVx3_ASAP7_75t_L g9207 ( 
.A(n_7809),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_7220),
.Y(n_9208)
);

OAI21x1_ASAP7_75t_L g9209 ( 
.A1(n_8041),
.A2(n_6884),
.B(n_6879),
.Y(n_9209)
);

A2O1A1Ixp33_ASAP7_75t_L g9210 ( 
.A1(n_7089),
.A2(n_6272),
.B(n_6319),
.C(n_6308),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_7454),
.Y(n_9211)
);

INVx2_ASAP7_75t_L g9212 ( 
.A(n_7220),
.Y(n_9212)
);

NAND2xp5_ASAP7_75t_L g9213 ( 
.A(n_7660),
.B(n_7675),
.Y(n_9213)
);

INVx3_ASAP7_75t_L g9214 ( 
.A(n_7809),
.Y(n_9214)
);

AOI21xp5_ASAP7_75t_L g9215 ( 
.A1(n_7655),
.A2(n_6393),
.B(n_6587),
.Y(n_9215)
);

OAI22xp5_ASAP7_75t_L g9216 ( 
.A1(n_7185),
.A2(n_6339),
.B1(n_6367),
.B2(n_6345),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_7454),
.Y(n_9217)
);

BUFx6f_ASAP7_75t_L g9218 ( 
.A(n_6949),
.Y(n_9218)
);

OAI21xp5_ASAP7_75t_L g9219 ( 
.A1(n_7439),
.A2(n_7780),
.B(n_7070),
.Y(n_9219)
);

AOI22xp33_ASAP7_75t_L g9220 ( 
.A1(n_7664),
.A2(n_8085),
.B1(n_7204),
.B2(n_7360),
.Y(n_9220)
);

OAI21x1_ASAP7_75t_L g9221 ( 
.A1(n_8041),
.A2(n_6892),
.B(n_6884),
.Y(n_9221)
);

AO21x2_ASAP7_75t_L g9222 ( 
.A1(n_7149),
.A2(n_5753),
.B(n_5730),
.Y(n_9222)
);

INVx3_ASAP7_75t_L g9223 ( 
.A(n_7809),
.Y(n_9223)
);

OAI21x1_ASAP7_75t_L g9224 ( 
.A1(n_6938),
.A2(n_6892),
.B(n_5861),
.Y(n_9224)
);

OAI22xp5_ASAP7_75t_L g9225 ( 
.A1(n_7185),
.A2(n_7360),
.B1(n_8050),
.B2(n_7522),
.Y(n_9225)
);

OAI21x1_ASAP7_75t_L g9226 ( 
.A1(n_6938),
.A2(n_5861),
.B(n_6344),
.Y(n_9226)
);

INVx1_ASAP7_75t_L g9227 ( 
.A(n_7457),
.Y(n_9227)
);

AO31x2_ASAP7_75t_L g9228 ( 
.A1(n_7972),
.A2(n_6091),
.A3(n_6098),
.B(n_6090),
.Y(n_9228)
);

A2O1A1Ixp33_ASAP7_75t_L g9229 ( 
.A1(n_7307),
.A2(n_6272),
.B(n_6319),
.C(n_6308),
.Y(n_9229)
);

BUFx3_ASAP7_75t_L g9230 ( 
.A(n_7819),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_7220),
.Y(n_9231)
);

OAI21x1_ASAP7_75t_L g9232 ( 
.A1(n_6938),
.A2(n_6347),
.B(n_6344),
.Y(n_9232)
);

OAI21x1_ASAP7_75t_L g9233 ( 
.A1(n_6939),
.A2(n_6347),
.B(n_6344),
.Y(n_9233)
);

OAI21x1_ASAP7_75t_L g9234 ( 
.A1(n_6939),
.A2(n_6353),
.B(n_6347),
.Y(n_9234)
);

O2A1O1Ixp33_ASAP7_75t_L g9235 ( 
.A1(n_7373),
.A2(n_5364),
.B(n_5365),
.C(n_5359),
.Y(n_9235)
);

OAI21x1_ASAP7_75t_L g9236 ( 
.A1(n_6939),
.A2(n_6353),
.B(n_6347),
.Y(n_9236)
);

INVx3_ASAP7_75t_L g9237 ( 
.A(n_7809),
.Y(n_9237)
);

AND2x4_ASAP7_75t_L g9238 ( 
.A(n_7682),
.B(n_6272),
.Y(n_9238)
);

NAND2xp5_ASAP7_75t_L g9239 ( 
.A(n_7660),
.B(n_6664),
.Y(n_9239)
);

AND2x4_ASAP7_75t_L g9240 ( 
.A(n_7706),
.B(n_6272),
.Y(n_9240)
);

INVx2_ASAP7_75t_L g9241 ( 
.A(n_6929),
.Y(n_9241)
);

CKINVDCx5p33_ASAP7_75t_R g9242 ( 
.A(n_7671),
.Y(n_9242)
);

INVx2_ASAP7_75t_L g9243 ( 
.A(n_6929),
.Y(n_9243)
);

AO21x2_ASAP7_75t_L g9244 ( 
.A1(n_7149),
.A2(n_5753),
.B(n_5730),
.Y(n_9244)
);

CKINVDCx8_ASAP7_75t_R g9245 ( 
.A(n_7103),
.Y(n_9245)
);

OAI21x1_ASAP7_75t_L g9246 ( 
.A1(n_7928),
.A2(n_7989),
.B(n_8077),
.Y(n_9246)
);

HB1xp67_ASAP7_75t_L g9247 ( 
.A(n_7586),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_7457),
.Y(n_9248)
);

OAI21x1_ASAP7_75t_L g9249 ( 
.A1(n_7928),
.A2(n_6375),
.B(n_6353),
.Y(n_9249)
);

A2O1A1Ixp33_ASAP7_75t_L g9250 ( 
.A1(n_7492),
.A2(n_6272),
.B(n_6319),
.C(n_6308),
.Y(n_9250)
);

INVx2_ASAP7_75t_SL g9251 ( 
.A(n_7706),
.Y(n_9251)
);

CKINVDCx9p33_ASAP7_75t_R g9252 ( 
.A(n_7669),
.Y(n_9252)
);

AO21x2_ASAP7_75t_L g9253 ( 
.A1(n_7149),
.A2(n_5760),
.B(n_5757),
.Y(n_9253)
);

INVx1_ASAP7_75t_L g9254 ( 
.A(n_7457),
.Y(n_9254)
);

NAND2xp5_ASAP7_75t_L g9255 ( 
.A(n_7675),
.B(n_6681),
.Y(n_9255)
);

OA21x2_ASAP7_75t_L g9256 ( 
.A1(n_7845),
.A2(n_6375),
.B(n_6353),
.Y(n_9256)
);

OAI21x1_ASAP7_75t_L g9257 ( 
.A1(n_7928),
.A2(n_6376),
.B(n_6375),
.Y(n_9257)
);

OAI21xp33_ASAP7_75t_L g9258 ( 
.A1(n_7522),
.A2(n_5844),
.B(n_6091),
.Y(n_9258)
);

OAI21x1_ASAP7_75t_L g9259 ( 
.A1(n_7989),
.A2(n_6376),
.B(n_6375),
.Y(n_9259)
);

AO21x2_ASAP7_75t_L g9260 ( 
.A1(n_7184),
.A2(n_5760),
.B(n_5757),
.Y(n_9260)
);

OAI21x1_ASAP7_75t_L g9261 ( 
.A1(n_7989),
.A2(n_6381),
.B(n_6376),
.Y(n_9261)
);

CKINVDCx5p33_ASAP7_75t_R g9262 ( 
.A(n_7671),
.Y(n_9262)
);

AND2x2_ASAP7_75t_L g9263 ( 
.A(n_8099),
.B(n_6351),
.Y(n_9263)
);

OA21x2_ASAP7_75t_L g9264 ( 
.A1(n_7845),
.A2(n_6396),
.B(n_6381),
.Y(n_9264)
);

OR2x2_ASAP7_75t_L g9265 ( 
.A(n_7518),
.B(n_7544),
.Y(n_9265)
);

BUFx2_ASAP7_75t_L g9266 ( 
.A(n_7162),
.Y(n_9266)
);

AOI22xp5_ASAP7_75t_L g9267 ( 
.A1(n_7702),
.A2(n_5998),
.B1(n_6030),
.B2(n_6007),
.Y(n_9267)
);

INVx1_ASAP7_75t_L g9268 ( 
.A(n_7461),
.Y(n_9268)
);

INVx1_ASAP7_75t_L g9269 ( 
.A(n_7461),
.Y(n_9269)
);

OAI21xp5_ASAP7_75t_L g9270 ( 
.A1(n_7883),
.A2(n_5793),
.B(n_5765),
.Y(n_9270)
);

AOI22xp33_ASAP7_75t_L g9271 ( 
.A1(n_7702),
.A2(n_6393),
.B1(n_6319),
.B2(n_6058),
.Y(n_9271)
);

INVx1_ASAP7_75t_L g9272 ( 
.A(n_7461),
.Y(n_9272)
);

AOI21xp33_ASAP7_75t_L g9273 ( 
.A1(n_7785),
.A2(n_5368),
.B(n_5367),
.Y(n_9273)
);

OAI21xp5_ASAP7_75t_L g9274 ( 
.A1(n_7883),
.A2(n_5793),
.B(n_5765),
.Y(n_9274)
);

OR2x6_ASAP7_75t_L g9275 ( 
.A(n_7351),
.B(n_6002),
.Y(n_9275)
);

INVx1_ASAP7_75t_SL g9276 ( 
.A(n_7235),
.Y(n_9276)
);

INVx4_ASAP7_75t_L g9277 ( 
.A(n_7282),
.Y(n_9277)
);

CKINVDCx20_ASAP7_75t_R g9278 ( 
.A(n_7531),
.Y(n_9278)
);

INVxp67_ASAP7_75t_L g9279 ( 
.A(n_7683),
.Y(n_9279)
);

INVx3_ASAP7_75t_L g9280 ( 
.A(n_7809),
.Y(n_9280)
);

OAI22xp33_ASAP7_75t_L g9281 ( 
.A1(n_7879),
.A2(n_6058),
.B1(n_6223),
.B2(n_6147),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_7466),
.Y(n_9282)
);

NAND2xp5_ASAP7_75t_SL g9283 ( 
.A(n_7580),
.B(n_6857),
.Y(n_9283)
);

AOI21xp5_ASAP7_75t_L g9284 ( 
.A1(n_7667),
.A2(n_6589),
.B(n_6822),
.Y(n_9284)
);

CKINVDCx20_ASAP7_75t_R g9285 ( 
.A(n_7609),
.Y(n_9285)
);

INVx3_ASAP7_75t_L g9286 ( 
.A(n_7809),
.Y(n_9286)
);

OAI21xp5_ASAP7_75t_L g9287 ( 
.A1(n_7926),
.A2(n_6397),
.B(n_6367),
.Y(n_9287)
);

AOI22xp5_ASAP7_75t_L g9288 ( 
.A1(n_7167),
.A2(n_7185),
.B1(n_8106),
.B2(n_8046),
.Y(n_9288)
);

INVx1_ASAP7_75t_L g9289 ( 
.A(n_7466),
.Y(n_9289)
);

NAND2xp33_ASAP7_75t_R g9290 ( 
.A(n_7753),
.B(n_6367),
.Y(n_9290)
);

INVx1_ASAP7_75t_SL g9291 ( 
.A(n_7235),
.Y(n_9291)
);

AO31x2_ASAP7_75t_L g9292 ( 
.A1(n_7763),
.A2(n_6113),
.A3(n_6119),
.B(n_6098),
.Y(n_9292)
);

AOI22xp33_ASAP7_75t_L g9293 ( 
.A1(n_7000),
.A2(n_6058),
.B1(n_6223),
.B2(n_6147),
.Y(n_9293)
);

AND2x4_ASAP7_75t_L g9294 ( 
.A(n_7706),
.B(n_6352),
.Y(n_9294)
);

OA21x2_ASAP7_75t_L g9295 ( 
.A1(n_7845),
.A2(n_6714),
.B(n_6682),
.Y(n_9295)
);

HB1xp67_ASAP7_75t_L g9296 ( 
.A(n_7586),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_7466),
.Y(n_9297)
);

BUFx3_ASAP7_75t_L g9298 ( 
.A(n_7819),
.Y(n_9298)
);

OAI22xp33_ASAP7_75t_L g9299 ( 
.A1(n_7879),
.A2(n_6058),
.B1(n_6223),
.B2(n_6147),
.Y(n_9299)
);

HB1xp67_ASAP7_75t_L g9300 ( 
.A(n_7592),
.Y(n_9300)
);

INVxp67_ASAP7_75t_SL g9301 ( 
.A(n_7683),
.Y(n_9301)
);

INVx1_ASAP7_75t_L g9302 ( 
.A(n_7467),
.Y(n_9302)
);

INVx1_ASAP7_75t_SL g9303 ( 
.A(n_7275),
.Y(n_9303)
);

AND2x2_ASAP7_75t_L g9304 ( 
.A(n_8103),
.B(n_6351),
.Y(n_9304)
);

OAI22xp5_ASAP7_75t_L g9305 ( 
.A1(n_7944),
.A2(n_6420),
.B1(n_6421),
.B2(n_6397),
.Y(n_9305)
);

A2O1A1Ixp33_ASAP7_75t_L g9306 ( 
.A1(n_7492),
.A2(n_6436),
.B(n_6826),
.C(n_6802),
.Y(n_9306)
);

OAI222xp33_ASAP7_75t_L g9307 ( 
.A1(n_7154),
.A2(n_6626),
.B1(n_6583),
.B2(n_5933),
.C1(n_5378),
.C2(n_5386),
.Y(n_9307)
);

INVx2_ASAP7_75t_L g9308 ( 
.A(n_6929),
.Y(n_9308)
);

INVx1_ASAP7_75t_L g9309 ( 
.A(n_7467),
.Y(n_9309)
);

NAND3xp33_ASAP7_75t_L g9310 ( 
.A(n_7551),
.B(n_5872),
.C(n_5868),
.Y(n_9310)
);

INVx2_ASAP7_75t_L g9311 ( 
.A(n_6929),
.Y(n_9311)
);

AO31x2_ASAP7_75t_L g9312 ( 
.A1(n_7685),
.A2(n_6124),
.A3(n_6131),
.B(n_6113),
.Y(n_9312)
);

INVx2_ASAP7_75t_SL g9313 ( 
.A(n_7732),
.Y(n_9313)
);

INVx1_ASAP7_75t_L g9314 ( 
.A(n_7467),
.Y(n_9314)
);

BUFx6f_ASAP7_75t_L g9315 ( 
.A(n_6949),
.Y(n_9315)
);

OA21x2_ASAP7_75t_L g9316 ( 
.A1(n_8073),
.A2(n_5783),
.B(n_5780),
.Y(n_9316)
);

HB1xp67_ASAP7_75t_L g9317 ( 
.A(n_7592),
.Y(n_9317)
);

BUFx2_ASAP7_75t_L g9318 ( 
.A(n_7174),
.Y(n_9318)
);

AO21x2_ASAP7_75t_L g9319 ( 
.A1(n_7184),
.A2(n_5783),
.B(n_5780),
.Y(n_9319)
);

NAND2xp5_ASAP7_75t_L g9320 ( 
.A(n_6948),
.B(n_6840),
.Y(n_9320)
);

OR2x2_ASAP7_75t_L g9321 ( 
.A(n_7518),
.B(n_6397),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_7469),
.Y(n_9322)
);

INVx2_ASAP7_75t_L g9323 ( 
.A(n_6931),
.Y(n_9323)
);

CKINVDCx20_ASAP7_75t_R g9324 ( 
.A(n_7609),
.Y(n_9324)
);

BUFx3_ASAP7_75t_L g9325 ( 
.A(n_7819),
.Y(n_9325)
);

AND2x4_ASAP7_75t_L g9326 ( 
.A(n_7732),
.B(n_6352),
.Y(n_9326)
);

AOI21xp5_ASAP7_75t_L g9327 ( 
.A1(n_7667),
.A2(n_6589),
.B(n_6822),
.Y(n_9327)
);

OR2x2_ASAP7_75t_L g9328 ( 
.A(n_7518),
.B(n_6420),
.Y(n_9328)
);

BUFx2_ASAP7_75t_L g9329 ( 
.A(n_7174),
.Y(n_9329)
);

INVx6_ASAP7_75t_L g9330 ( 
.A(n_7568),
.Y(n_9330)
);

NAND2x1p5_ASAP7_75t_L g9331 ( 
.A(n_7144),
.B(n_6436),
.Y(n_9331)
);

NAND3xp33_ASAP7_75t_L g9332 ( 
.A(n_7551),
.B(n_7926),
.C(n_7460),
.Y(n_9332)
);

OAI21xp5_ASAP7_75t_L g9333 ( 
.A1(n_7629),
.A2(n_8120),
.B(n_7807),
.Y(n_9333)
);

BUFx2_ASAP7_75t_L g9334 ( 
.A(n_7174),
.Y(n_9334)
);

BUFx6f_ASAP7_75t_L g9335 ( 
.A(n_6949),
.Y(n_9335)
);

BUFx6f_ASAP7_75t_L g9336 ( 
.A(n_6949),
.Y(n_9336)
);

NAND2x1p5_ASAP7_75t_L g9337 ( 
.A(n_7144),
.B(n_6436),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_7469),
.Y(n_9338)
);

NOR2xp33_ASAP7_75t_L g9339 ( 
.A(n_7874),
.B(n_6479),
.Y(n_9339)
);

AOI22xp33_ASAP7_75t_L g9340 ( 
.A1(n_7000),
.A2(n_6058),
.B1(n_6223),
.B2(n_6147),
.Y(n_9340)
);

OAI21x1_ASAP7_75t_SL g9341 ( 
.A1(n_7109),
.A2(n_6075),
.B(n_6151),
.Y(n_9341)
);

BUFx2_ASAP7_75t_L g9342 ( 
.A(n_7192),
.Y(n_9342)
);

AO31x2_ASAP7_75t_L g9343 ( 
.A1(n_7685),
.A2(n_6124),
.A3(n_6131),
.B(n_6119),
.Y(n_9343)
);

BUFx3_ASAP7_75t_L g9344 ( 
.A(n_7821),
.Y(n_9344)
);

OAI21xp5_ASAP7_75t_L g9345 ( 
.A1(n_7629),
.A2(n_6421),
.B(n_6420),
.Y(n_9345)
);

NOR2xp33_ASAP7_75t_L g9346 ( 
.A(n_7874),
.B(n_6479),
.Y(n_9346)
);

OR2x2_ASAP7_75t_L g9347 ( 
.A(n_7544),
.B(n_6421),
.Y(n_9347)
);

NOR2xp67_ASAP7_75t_L g9348 ( 
.A(n_7154),
.B(n_6533),
.Y(n_9348)
);

NAND2xp5_ASAP7_75t_L g9349 ( 
.A(n_6948),
.B(n_6840),
.Y(n_9349)
);

INVx2_ASAP7_75t_SL g9350 ( 
.A(n_7732),
.Y(n_9350)
);

INVx2_ASAP7_75t_L g9351 ( 
.A(n_6931),
.Y(n_9351)
);

NOR2xp33_ASAP7_75t_L g9352 ( 
.A(n_7944),
.B(n_6479),
.Y(n_9352)
);

OAI21xp5_ASAP7_75t_L g9353 ( 
.A1(n_8120),
.A2(n_6429),
.B(n_6425),
.Y(n_9353)
);

NOR2xp67_ASAP7_75t_L g9354 ( 
.A(n_7182),
.B(n_6533),
.Y(n_9354)
);

AOI21xp5_ASAP7_75t_L g9355 ( 
.A1(n_7680),
.A2(n_6151),
.B(n_6075),
.Y(n_9355)
);

AOI22x1_ASAP7_75t_L g9356 ( 
.A1(n_7493),
.A2(n_6584),
.B1(n_6741),
.B2(n_6574),
.Y(n_9356)
);

AO21x2_ASAP7_75t_L g9357 ( 
.A1(n_7184),
.A2(n_5795),
.B(n_5794),
.Y(n_9357)
);

AND2x6_ASAP7_75t_L g9358 ( 
.A(n_7795),
.B(n_4518),
.Y(n_9358)
);

INVx2_ASAP7_75t_L g9359 ( 
.A(n_6931),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_7469),
.Y(n_9360)
);

BUFx2_ASAP7_75t_SL g9361 ( 
.A(n_7157),
.Y(n_9361)
);

OA21x2_ASAP7_75t_L g9362 ( 
.A1(n_8073),
.A2(n_5814),
.B(n_5798),
.Y(n_9362)
);

OAI21xp5_ASAP7_75t_L g9363 ( 
.A1(n_7807),
.A2(n_6429),
.B(n_6425),
.Y(n_9363)
);

HB1xp67_ASAP7_75t_L g9364 ( 
.A(n_7640),
.Y(n_9364)
);

INVx1_ASAP7_75t_L g9365 ( 
.A(n_7471),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_6931),
.Y(n_9366)
);

OR2x2_ASAP7_75t_L g9367 ( 
.A(n_7544),
.B(n_6425),
.Y(n_9367)
);

OAI21xp5_ASAP7_75t_L g9368 ( 
.A1(n_7742),
.A2(n_6440),
.B(n_6429),
.Y(n_9368)
);

OR2x2_ASAP7_75t_L g9369 ( 
.A(n_7544),
.B(n_6440),
.Y(n_9369)
);

CKINVDCx5p33_ASAP7_75t_R g9370 ( 
.A(n_7746),
.Y(n_9370)
);

NAND2xp5_ASAP7_75t_L g9371 ( 
.A(n_6948),
.B(n_6132),
.Y(n_9371)
);

NAND2xp5_ASAP7_75t_L g9372 ( 
.A(n_6961),
.B(n_6132),
.Y(n_9372)
);

AO21x2_ASAP7_75t_L g9373 ( 
.A1(n_7069),
.A2(n_5820),
.B(n_5818),
.Y(n_9373)
);

NAND2xp5_ASAP7_75t_L g9374 ( 
.A(n_6961),
.B(n_6135),
.Y(n_9374)
);

AOI22xp33_ASAP7_75t_L g9375 ( 
.A1(n_7451),
.A2(n_6147),
.B1(n_6263),
.B2(n_6223),
.Y(n_9375)
);

INVx2_ASAP7_75t_L g9376 ( 
.A(n_6944),
.Y(n_9376)
);

INVx5_ASAP7_75t_SL g9377 ( 
.A(n_7840),
.Y(n_9377)
);

AOI21xp5_ASAP7_75t_L g9378 ( 
.A1(n_7680),
.A2(n_7373),
.B(n_7106),
.Y(n_9378)
);

INVx1_ASAP7_75t_L g9379 ( 
.A(n_7471),
.Y(n_9379)
);

OAI22xp5_ASAP7_75t_L g9380 ( 
.A1(n_7959),
.A2(n_6440),
.B1(n_5844),
.B2(n_5896),
.Y(n_9380)
);

INVx1_ASAP7_75t_L g9381 ( 
.A(n_7471),
.Y(n_9381)
);

AND2x4_ASAP7_75t_L g9382 ( 
.A(n_7732),
.B(n_6352),
.Y(n_9382)
);

OA21x2_ASAP7_75t_L g9383 ( 
.A1(n_8073),
.A2(n_5825),
.B(n_5820),
.Y(n_9383)
);

O2A1O1Ixp33_ASAP7_75t_SL g9384 ( 
.A1(n_7929),
.A2(n_6848),
.B(n_6826),
.C(n_6184),
.Y(n_9384)
);

INVx2_ASAP7_75t_L g9385 ( 
.A(n_6944),
.Y(n_9385)
);

NAND2xp5_ASAP7_75t_L g9386 ( 
.A(n_6961),
.B(n_6963),
.Y(n_9386)
);

INVx4_ASAP7_75t_SL g9387 ( 
.A(n_7393),
.Y(n_9387)
);

INVx1_ASAP7_75t_L g9388 ( 
.A(n_7473),
.Y(n_9388)
);

INVx2_ASAP7_75t_L g9389 ( 
.A(n_6944),
.Y(n_9389)
);

AO32x2_ASAP7_75t_L g9390 ( 
.A1(n_7182),
.A2(n_6898),
.A3(n_6902),
.B1(n_6816),
.B2(n_6762),
.Y(n_9390)
);

INVx1_ASAP7_75t_L g9391 ( 
.A(n_7473),
.Y(n_9391)
);

NAND2xp5_ASAP7_75t_L g9392 ( 
.A(n_6963),
.B(n_6135),
.Y(n_9392)
);

HB1xp67_ASAP7_75t_L g9393 ( 
.A(n_7640),
.Y(n_9393)
);

NAND2xp5_ASAP7_75t_L g9394 ( 
.A(n_6963),
.B(n_6137),
.Y(n_9394)
);

CKINVDCx14_ASAP7_75t_R g9395 ( 
.A(n_7491),
.Y(n_9395)
);

NOR2xp33_ASAP7_75t_L g9396 ( 
.A(n_7959),
.B(n_6479),
.Y(n_9396)
);

AOI22xp33_ASAP7_75t_L g9397 ( 
.A1(n_7451),
.A2(n_6263),
.B1(n_6337),
.B2(n_6323),
.Y(n_9397)
);

AO21x2_ASAP7_75t_L g9398 ( 
.A1(n_7069),
.A2(n_5379),
.B(n_5378),
.Y(n_9398)
);

AND2x4_ASAP7_75t_L g9399 ( 
.A(n_7759),
.B(n_6352),
.Y(n_9399)
);

AOI21xp5_ASAP7_75t_L g9400 ( 
.A1(n_7069),
.A2(n_6184),
.B(n_6172),
.Y(n_9400)
);

A2O1A1Ixp33_ASAP7_75t_L g9401 ( 
.A1(n_7530),
.A2(n_6436),
.B(n_6848),
.C(n_5729),
.Y(n_9401)
);

OA21x2_ASAP7_75t_L g9402 ( 
.A1(n_8102),
.A2(n_5966),
.B(n_5956),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_7473),
.Y(n_9403)
);

BUFx6f_ASAP7_75t_L g9404 ( 
.A(n_6949),
.Y(n_9404)
);

OAI21xp5_ASAP7_75t_L g9405 ( 
.A1(n_7742),
.A2(n_5872),
.B(n_5868),
.Y(n_9405)
);

BUFx2_ASAP7_75t_L g9406 ( 
.A(n_7192),
.Y(n_9406)
);

NAND2xp5_ASAP7_75t_L g9407 ( 
.A(n_6969),
.B(n_7106),
.Y(n_9407)
);

NAND2xp5_ASAP7_75t_L g9408 ( 
.A(n_6969),
.B(n_6137),
.Y(n_9408)
);

NAND2xp5_ASAP7_75t_L g9409 ( 
.A(n_6969),
.B(n_6138),
.Y(n_9409)
);

AOI21xp5_ASAP7_75t_SL g9410 ( 
.A1(n_7662),
.A2(n_6184),
.B(n_6172),
.Y(n_9410)
);

NOR2xp33_ASAP7_75t_SL g9411 ( 
.A(n_7413),
.B(n_6263),
.Y(n_9411)
);

INVx1_ASAP7_75t_L g9412 ( 
.A(n_7476),
.Y(n_9412)
);

AO21x2_ASAP7_75t_L g9413 ( 
.A1(n_7106),
.A2(n_5386),
.B(n_5379),
.Y(n_9413)
);

CKINVDCx6p67_ASAP7_75t_R g9414 ( 
.A(n_7282),
.Y(n_9414)
);

AOI22xp33_ASAP7_75t_L g9415 ( 
.A1(n_7460),
.A2(n_6263),
.B1(n_6337),
.B2(n_6323),
.Y(n_9415)
);

OAI21xp5_ASAP7_75t_L g9416 ( 
.A1(n_7784),
.A2(n_5143),
.B(n_5138),
.Y(n_9416)
);

AO21x2_ASAP7_75t_L g9417 ( 
.A1(n_7116),
.A2(n_7865),
.B(n_7847),
.Y(n_9417)
);

OAI21x1_ASAP7_75t_SL g9418 ( 
.A1(n_7362),
.A2(n_7402),
.B(n_7032),
.Y(n_9418)
);

INVx2_ASAP7_75t_L g9419 ( 
.A(n_6944),
.Y(n_9419)
);

INVx2_ASAP7_75t_L g9420 ( 
.A(n_6950),
.Y(n_9420)
);

OAI21x1_ASAP7_75t_L g9421 ( 
.A1(n_7804),
.A2(n_7843),
.B(n_7876),
.Y(n_9421)
);

INVx2_ASAP7_75t_L g9422 ( 
.A(n_6950),
.Y(n_9422)
);

AO32x2_ASAP7_75t_L g9423 ( 
.A1(n_7182),
.A2(n_6898),
.A3(n_6902),
.B1(n_6816),
.B2(n_6762),
.Y(n_9423)
);

NAND2xp5_ASAP7_75t_L g9424 ( 
.A(n_7116),
.B(n_6138),
.Y(n_9424)
);

OAI21xp5_ASAP7_75t_L g9425 ( 
.A1(n_7784),
.A2(n_5148),
.B(n_5145),
.Y(n_9425)
);

O2A1O1Ixp33_ASAP7_75t_SL g9426 ( 
.A1(n_7776),
.A2(n_6213),
.B(n_6214),
.C(n_6188),
.Y(n_9426)
);

INVx8_ASAP7_75t_L g9427 ( 
.A(n_7282),
.Y(n_9427)
);

AOI21xp5_ASAP7_75t_L g9428 ( 
.A1(n_7116),
.A2(n_6213),
.B(n_6188),
.Y(n_9428)
);

NOR2xp33_ASAP7_75t_SL g9429 ( 
.A(n_7674),
.B(n_6263),
.Y(n_9429)
);

AND2x2_ASAP7_75t_L g9430 ( 
.A(n_8103),
.B(n_6351),
.Y(n_9430)
);

AOI21xp33_ASAP7_75t_L g9431 ( 
.A1(n_7847),
.A2(n_7878),
.B(n_7865),
.Y(n_9431)
);

AOI221x1_ASAP7_75t_L g9432 ( 
.A1(n_7808),
.A2(n_5399),
.B1(n_5395),
.B2(n_5176),
.C(n_5179),
.Y(n_9432)
);

OAI22xp5_ASAP7_75t_L g9433 ( 
.A1(n_7580),
.A2(n_5844),
.B1(n_6893),
.B2(n_6369),
.Y(n_9433)
);

NOR2xp33_ASAP7_75t_L g9434 ( 
.A(n_8011),
.B(n_6479),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_7476),
.Y(n_9435)
);

CKINVDCx11_ASAP7_75t_R g9436 ( 
.A(n_7275),
.Y(n_9436)
);

OR2x2_ASAP7_75t_L g9437 ( 
.A(n_7705),
.B(n_6142),
.Y(n_9437)
);

NAND2xp5_ASAP7_75t_L g9438 ( 
.A(n_7847),
.B(n_7865),
.Y(n_9438)
);

INVx5_ASAP7_75t_L g9439 ( 
.A(n_7821),
.Y(n_9439)
);

BUFx10_ASAP7_75t_L g9440 ( 
.A(n_7493),
.Y(n_9440)
);

INVx1_ASAP7_75t_L g9441 ( 
.A(n_7476),
.Y(n_9441)
);

OAI22xp5_ASAP7_75t_L g9442 ( 
.A1(n_7580),
.A2(n_7825),
.B1(n_7218),
.B2(n_8011),
.Y(n_9442)
);

OR2x2_ASAP7_75t_L g9443 ( 
.A(n_7705),
.B(n_6142),
.Y(n_9443)
);

INVx3_ASAP7_75t_L g9444 ( 
.A(n_7809),
.Y(n_9444)
);

INVx3_ASAP7_75t_L g9445 ( 
.A(n_7809),
.Y(n_9445)
);

AND2x4_ASAP7_75t_L g9446 ( 
.A(n_7759),
.B(n_6352),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_7481),
.Y(n_9447)
);

NAND2x1p5_ASAP7_75t_L g9448 ( 
.A(n_7144),
.B(n_6436),
.Y(n_9448)
);

AOI21xp5_ASAP7_75t_L g9449 ( 
.A1(n_7878),
.A2(n_6213),
.B(n_6188),
.Y(n_9449)
);

OAI21x1_ASAP7_75t_L g9450 ( 
.A1(n_7843),
.A2(n_8012),
.B(n_7876),
.Y(n_9450)
);

NAND2xp5_ASAP7_75t_L g9451 ( 
.A(n_7878),
.B(n_6168),
.Y(n_9451)
);

INVx2_ASAP7_75t_L g9452 ( 
.A(n_6950),
.Y(n_9452)
);

AOI22xp5_ASAP7_75t_L g9453 ( 
.A1(n_7167),
.A2(n_5998),
.B1(n_6030),
.B2(n_6007),
.Y(n_9453)
);

AOI22xp33_ASAP7_75t_L g9454 ( 
.A1(n_7171),
.A2(n_6323),
.B1(n_6340),
.B2(n_6337),
.Y(n_9454)
);

INVx1_ASAP7_75t_L g9455 ( 
.A(n_7481),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_7481),
.Y(n_9456)
);

INVx3_ASAP7_75t_SL g9457 ( 
.A(n_7103),
.Y(n_9457)
);

OA21x2_ASAP7_75t_L g9458 ( 
.A1(n_8102),
.A2(n_5966),
.B(n_5956),
.Y(n_9458)
);

INVx2_ASAP7_75t_L g9459 ( 
.A(n_6950),
.Y(n_9459)
);

BUFx3_ASAP7_75t_L g9460 ( 
.A(n_7821),
.Y(n_9460)
);

OAI21xp5_ASAP7_75t_L g9461 ( 
.A1(n_7571),
.A2(n_5148),
.B(n_5145),
.Y(n_9461)
);

HB1xp67_ASAP7_75t_L g9462 ( 
.A(n_7663),
.Y(n_9462)
);

INVxp67_ASAP7_75t_SL g9463 ( 
.A(n_7119),
.Y(n_9463)
);

OAI21x1_ASAP7_75t_L g9464 ( 
.A1(n_7843),
.A2(n_8012),
.B(n_7876),
.Y(n_9464)
);

OAI21xp5_ASAP7_75t_L g9465 ( 
.A1(n_7571),
.A2(n_5159),
.B(n_5152),
.Y(n_9465)
);

CKINVDCx16_ASAP7_75t_R g9466 ( 
.A(n_7491),
.Y(n_9466)
);

NAND2xp5_ASAP7_75t_L g9467 ( 
.A(n_7815),
.B(n_6168),
.Y(n_9467)
);

OAI21x1_ASAP7_75t_L g9468 ( 
.A1(n_7843),
.A2(n_8012),
.B(n_7876),
.Y(n_9468)
);

INVx1_ASAP7_75t_L g9469 ( 
.A(n_7497),
.Y(n_9469)
);

OAI22xp5_ASAP7_75t_L g9470 ( 
.A1(n_7580),
.A2(n_6893),
.B1(n_6369),
.B2(n_6857),
.Y(n_9470)
);

BUFx4_ASAP7_75t_SL g9471 ( 
.A(n_7670),
.Y(n_9471)
);

NAND2x1p5_ASAP7_75t_L g9472 ( 
.A(n_7144),
.B(n_6436),
.Y(n_9472)
);

OAI21x1_ASAP7_75t_SL g9473 ( 
.A1(n_7362),
.A2(n_6214),
.B(n_6253),
.Y(n_9473)
);

AO31x2_ASAP7_75t_L g9474 ( 
.A1(n_7685),
.A2(n_6173),
.A3(n_6206),
.B(n_6171),
.Y(n_9474)
);

OA21x2_ASAP7_75t_L g9475 ( 
.A1(n_8102),
.A2(n_5966),
.B(n_5956),
.Y(n_9475)
);

INVx2_ASAP7_75t_SL g9476 ( 
.A(n_7759),
.Y(n_9476)
);

AOI22xp33_ASAP7_75t_L g9477 ( 
.A1(n_7171),
.A2(n_6323),
.B1(n_6340),
.B2(n_6337),
.Y(n_9477)
);

OAI221xp5_ASAP7_75t_L g9478 ( 
.A1(n_7611),
.A2(n_7622),
.B1(n_7218),
.B2(n_7124),
.C(n_7147),
.Y(n_9478)
);

OA21x2_ASAP7_75t_L g9479 ( 
.A1(n_6990),
.A2(n_5978),
.B(n_5972),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_7497),
.Y(n_9480)
);

INVx1_ASAP7_75t_L g9481 ( 
.A(n_7497),
.Y(n_9481)
);

OAI221xp5_ASAP7_75t_L g9482 ( 
.A1(n_7611),
.A2(n_5933),
.B1(n_5649),
.B2(n_5159),
.C(n_5168),
.Y(n_9482)
);

OR2x2_ASAP7_75t_L g9483 ( 
.A(n_7705),
.B(n_6171),
.Y(n_9483)
);

INVx2_ASAP7_75t_SL g9484 ( 
.A(n_7759),
.Y(n_9484)
);

INVx6_ASAP7_75t_L g9485 ( 
.A(n_7568),
.Y(n_9485)
);

OAI21x1_ASAP7_75t_L g9486 ( 
.A1(n_6954),
.A2(n_6231),
.B(n_6219),
.Y(n_9486)
);

AND2x4_ASAP7_75t_L g9487 ( 
.A(n_7800),
.B(n_6358),
.Y(n_9487)
);

OAI21x1_ASAP7_75t_L g9488 ( 
.A1(n_6954),
.A2(n_6238),
.B(n_6231),
.Y(n_9488)
);

AOI21xp5_ASAP7_75t_L g9489 ( 
.A1(n_7358),
.A2(n_6253),
.B(n_6214),
.Y(n_9489)
);

OAI21x1_ASAP7_75t_SL g9490 ( 
.A1(n_7362),
.A2(n_6310),
.B(n_6338),
.Y(n_9490)
);

OAI21xp5_ASAP7_75t_L g9491 ( 
.A1(n_7717),
.A2(n_5165),
.B(n_5152),
.Y(n_9491)
);

INVx1_ASAP7_75t_L g9492 ( 
.A(n_7499),
.Y(n_9492)
);

INVx2_ASAP7_75t_L g9493 ( 
.A(n_6952),
.Y(n_9493)
);

AOI21xp5_ASAP7_75t_L g9494 ( 
.A1(n_7358),
.A2(n_6310),
.B(n_5763),
.Y(n_9494)
);

AND2x4_ASAP7_75t_L g9495 ( 
.A(n_7800),
.B(n_6358),
.Y(n_9495)
);

BUFx3_ASAP7_75t_L g9496 ( 
.A(n_7821),
.Y(n_9496)
);

AOI22xp33_ASAP7_75t_L g9497 ( 
.A1(n_7835),
.A2(n_6323),
.B1(n_6340),
.B2(n_6337),
.Y(n_9497)
);

BUFx3_ASAP7_75t_L g9498 ( 
.A(n_7821),
.Y(n_9498)
);

INVx2_ASAP7_75t_L g9499 ( 
.A(n_6952),
.Y(n_9499)
);

INVx4_ASAP7_75t_L g9500 ( 
.A(n_7282),
.Y(n_9500)
);

AOI22xp33_ASAP7_75t_SL g9501 ( 
.A1(n_7197),
.A2(n_6436),
.B1(n_6030),
.B2(n_6007),
.Y(n_9501)
);

INVx1_ASAP7_75t_L g9502 ( 
.A(n_7499),
.Y(n_9502)
);

AO21x2_ASAP7_75t_L g9503 ( 
.A1(n_7717),
.A2(n_5978),
.B(n_5972),
.Y(n_9503)
);

AOI22xp33_ASAP7_75t_L g9504 ( 
.A1(n_7835),
.A2(n_6340),
.B1(n_6405),
.B2(n_6371),
.Y(n_9504)
);

OAI21xp5_ASAP7_75t_L g9505 ( 
.A1(n_7717),
.A2(n_5168),
.B(n_5165),
.Y(n_9505)
);

INVx2_ASAP7_75t_L g9506 ( 
.A(n_6952),
.Y(n_9506)
);

BUFx6f_ASAP7_75t_L g9507 ( 
.A(n_6949),
.Y(n_9507)
);

OAI21x1_ASAP7_75t_L g9508 ( 
.A1(n_6954),
.A2(n_7027),
.B(n_6972),
.Y(n_9508)
);

AND2x6_ASAP7_75t_L g9509 ( 
.A(n_7795),
.B(n_7736),
.Y(n_9509)
);

AND2x4_ASAP7_75t_L g9510 ( 
.A(n_7800),
.B(n_6358),
.Y(n_9510)
);

BUFx2_ASAP7_75t_SL g9511 ( 
.A(n_7341),
.Y(n_9511)
);

OAI21x1_ASAP7_75t_L g9512 ( 
.A1(n_6954),
.A2(n_7027),
.B(n_6972),
.Y(n_9512)
);

OR2x2_ASAP7_75t_L g9513 ( 
.A(n_7705),
.B(n_6173),
.Y(n_9513)
);

AO21x2_ASAP7_75t_L g9514 ( 
.A1(n_7621),
.A2(n_5978),
.B(n_5972),
.Y(n_9514)
);

AOI221x1_ASAP7_75t_L g9515 ( 
.A1(n_7288),
.A2(n_5395),
.B1(n_5176),
.B2(n_5179),
.C(n_5169),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_7499),
.Y(n_9516)
);

BUFx3_ASAP7_75t_L g9517 ( 
.A(n_7821),
.Y(n_9517)
);

OAI22xp33_ASAP7_75t_L g9518 ( 
.A1(n_7879),
.A2(n_6340),
.B1(n_6405),
.B2(n_6371),
.Y(n_9518)
);

INVx2_ASAP7_75t_SL g9519 ( 
.A(n_7800),
.Y(n_9519)
);

CKINVDCx5p33_ASAP7_75t_R g9520 ( 
.A(n_7746),
.Y(n_9520)
);

OA21x2_ASAP7_75t_L g9521 ( 
.A1(n_6990),
.A2(n_5996),
.B(n_5992),
.Y(n_9521)
);

HB1xp67_ASAP7_75t_L g9522 ( 
.A(n_7663),
.Y(n_9522)
);

OR2x2_ASAP7_75t_L g9523 ( 
.A(n_7197),
.B(n_6177),
.Y(n_9523)
);

OA21x2_ASAP7_75t_L g9524 ( 
.A1(n_7206),
.A2(n_5996),
.B(n_5992),
.Y(n_9524)
);

A2O1A1Ixp33_ASAP7_75t_L g9525 ( 
.A1(n_7530),
.A2(n_6436),
.B(n_5759),
.C(n_5767),
.Y(n_9525)
);

OAI21x1_ASAP7_75t_L g9526 ( 
.A1(n_6954),
.A2(n_6238),
.B(n_6231),
.Y(n_9526)
);

NOR2xp33_ASAP7_75t_SL g9527 ( 
.A(n_7674),
.B(n_6371),
.Y(n_9527)
);

OAI21x1_ASAP7_75t_L g9528 ( 
.A1(n_6972),
.A2(n_6264),
.B(n_6238),
.Y(n_9528)
);

NOR2xp33_ASAP7_75t_L g9529 ( 
.A(n_7884),
.B(n_6369),
.Y(n_9529)
);

OR2x2_ASAP7_75t_L g9530 ( 
.A(n_7197),
.B(n_7288),
.Y(n_9530)
);

AND2x4_ASAP7_75t_L g9531 ( 
.A(n_7805),
.B(n_6358),
.Y(n_9531)
);

INVx2_ASAP7_75t_L g9532 ( 
.A(n_6952),
.Y(n_9532)
);

OAI21x1_ASAP7_75t_L g9533 ( 
.A1(n_6972),
.A2(n_6264),
.B(n_6238),
.Y(n_9533)
);

AOI22xp33_ASAP7_75t_SL g9534 ( 
.A1(n_7197),
.A2(n_6030),
.B1(n_6007),
.B2(n_5729),
.Y(n_9534)
);

AO31x2_ASAP7_75t_L g9535 ( 
.A1(n_7602),
.A2(n_6210),
.A3(n_6222),
.B(n_6177),
.Y(n_9535)
);

BUFx8_ASAP7_75t_L g9536 ( 
.A(n_7283),
.Y(n_9536)
);

OAI21x1_ASAP7_75t_SL g9537 ( 
.A1(n_7402),
.A2(n_6310),
.B(n_6338),
.Y(n_9537)
);

AND2x2_ASAP7_75t_L g9538 ( 
.A(n_8103),
.B(n_6518),
.Y(n_9538)
);

AND2x2_ASAP7_75t_L g9539 ( 
.A(n_8114),
.B(n_6518),
.Y(n_9539)
);

NOR2xp33_ASAP7_75t_L g9540 ( 
.A(n_7884),
.B(n_6238),
.Y(n_9540)
);

OAI21x1_ASAP7_75t_L g9541 ( 
.A1(n_6972),
.A2(n_6282),
.B(n_6264),
.Y(n_9541)
);

OAI21x1_ASAP7_75t_L g9542 ( 
.A1(n_7027),
.A2(n_6282),
.B(n_6264),
.Y(n_9542)
);

AO21x2_ASAP7_75t_L g9543 ( 
.A1(n_7621),
.A2(n_5996),
.B(n_5992),
.Y(n_9543)
);

AOI21xp5_ASAP7_75t_L g9544 ( 
.A1(n_7358),
.A2(n_7438),
.B(n_7435),
.Y(n_9544)
);

OA21x2_ASAP7_75t_L g9545 ( 
.A1(n_7206),
.A2(n_6021),
.B(n_6004),
.Y(n_9545)
);

OAI21x1_ASAP7_75t_L g9546 ( 
.A1(n_7027),
.A2(n_6282),
.B(n_6264),
.Y(n_9546)
);

OAI21x1_ASAP7_75t_L g9547 ( 
.A1(n_7027),
.A2(n_6291),
.B(n_6282),
.Y(n_9547)
);

NOR2xp33_ASAP7_75t_L g9548 ( 
.A(n_7884),
.B(n_6282),
.Y(n_9548)
);

INVx1_ASAP7_75t_L g9549 ( 
.A(n_7504),
.Y(n_9549)
);

OAI21xp5_ASAP7_75t_L g9550 ( 
.A1(n_7662),
.A2(n_5173),
.B(n_5172),
.Y(n_9550)
);

OAI21x1_ASAP7_75t_L g9551 ( 
.A1(n_7055),
.A2(n_6307),
.B(n_6291),
.Y(n_9551)
);

OAI21x1_ASAP7_75t_L g9552 ( 
.A1(n_7055),
.A2(n_6307),
.B(n_6291),
.Y(n_9552)
);

AOI21xp33_ASAP7_75t_L g9553 ( 
.A1(n_7288),
.A2(n_5140),
.B(n_5162),
.Y(n_9553)
);

INVx1_ASAP7_75t_L g9554 ( 
.A(n_7504),
.Y(n_9554)
);

HB1xp67_ASAP7_75t_L g9555 ( 
.A(n_7711),
.Y(n_9555)
);

INVx1_ASAP7_75t_SL g9556 ( 
.A(n_7670),
.Y(n_9556)
);

OAI21x1_ASAP7_75t_L g9557 ( 
.A1(n_7055),
.A2(n_6307),
.B(n_6291),
.Y(n_9557)
);

OAI21x1_ASAP7_75t_L g9558 ( 
.A1(n_7055),
.A2(n_7274),
.B(n_8019),
.Y(n_9558)
);

OAI21x1_ASAP7_75t_L g9559 ( 
.A1(n_7055),
.A2(n_6307),
.B(n_6291),
.Y(n_9559)
);

AO21x2_ASAP7_75t_L g9560 ( 
.A1(n_7891),
.A2(n_6021),
.B(n_6004),
.Y(n_9560)
);

OAI22xp5_ASAP7_75t_L g9561 ( 
.A1(n_7825),
.A2(n_6893),
.B1(n_6857),
.B2(n_6128),
.Y(n_9561)
);

OAI22xp33_ASAP7_75t_L g9562 ( 
.A1(n_7462),
.A2(n_6371),
.B1(n_6411),
.B2(n_6405),
.Y(n_9562)
);

OAI21xp5_ASAP7_75t_L g9563 ( 
.A1(n_8007),
.A2(n_5173),
.B(n_5172),
.Y(n_9563)
);

NAND2xp5_ASAP7_75t_L g9564 ( 
.A(n_7815),
.B(n_6206),
.Y(n_9564)
);

AND2x2_ASAP7_75t_L g9565 ( 
.A(n_8114),
.B(n_8123),
.Y(n_9565)
);

O2A1O1Ixp33_ASAP7_75t_L g9566 ( 
.A1(n_8075),
.A2(n_5706),
.B(n_5179),
.C(n_5169),
.Y(n_9566)
);

AND2x2_ASAP7_75t_L g9567 ( 
.A(n_8114),
.B(n_8123),
.Y(n_9567)
);

INVx2_ASAP7_75t_L g9568 ( 
.A(n_6988),
.Y(n_9568)
);

AND2x2_ASAP7_75t_L g9569 ( 
.A(n_8114),
.B(n_6518),
.Y(n_9569)
);

AOI21xp5_ASAP7_75t_L g9570 ( 
.A1(n_7435),
.A2(n_5763),
.B(n_6837),
.Y(n_9570)
);

INVx1_ASAP7_75t_L g9571 ( 
.A(n_7504),
.Y(n_9571)
);

OAI21x1_ASAP7_75t_L g9572 ( 
.A1(n_7274),
.A2(n_6326),
.B(n_6307),
.Y(n_9572)
);

OAI21x1_ASAP7_75t_L g9573 ( 
.A1(n_7274),
.A2(n_6328),
.B(n_6326),
.Y(n_9573)
);

NAND2xp5_ASAP7_75t_L g9574 ( 
.A(n_7815),
.B(n_6210),
.Y(n_9574)
);

AOI22xp33_ASAP7_75t_L g9575 ( 
.A1(n_7622),
.A2(n_6371),
.B1(n_6411),
.B2(n_6405),
.Y(n_9575)
);

AO31x2_ASAP7_75t_L g9576 ( 
.A1(n_7602),
.A2(n_6229),
.A3(n_6261),
.B(n_6233),
.Y(n_9576)
);

NAND2xp5_ASAP7_75t_L g9577 ( 
.A(n_7820),
.B(n_6222),
.Y(n_9577)
);

OA21x2_ASAP7_75t_L g9578 ( 
.A1(n_7295),
.A2(n_7377),
.B(n_7353),
.Y(n_9578)
);

AO31x2_ASAP7_75t_L g9579 ( 
.A1(n_7602),
.A2(n_6233),
.A3(n_6261),
.B(n_6229),
.Y(n_9579)
);

AND2x2_ASAP7_75t_L g9580 ( 
.A(n_8123),
.B(n_6518),
.Y(n_9580)
);

INVx1_ASAP7_75t_L g9581 ( 
.A(n_8135),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_8135),
.Y(n_9582)
);

INVx1_ASAP7_75t_L g9583 ( 
.A(n_8215),
.Y(n_9583)
);

BUFx2_ASAP7_75t_L g9584 ( 
.A(n_8177),
.Y(n_9584)
);

AOI22xp33_ASAP7_75t_L g9585 ( 
.A1(n_8271),
.A2(n_7712),
.B1(n_7710),
.B2(n_7650),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_8215),
.Y(n_9586)
);

INVx3_ASAP7_75t_L g9587 ( 
.A(n_8177),
.Y(n_9587)
);

INVx1_ASAP7_75t_SL g9588 ( 
.A(n_9071),
.Y(n_9588)
);

AOI21x1_ASAP7_75t_L g9589 ( 
.A1(n_8161),
.A2(n_7935),
.B(n_7925),
.Y(n_9589)
);

AO21x2_ASAP7_75t_L g9590 ( 
.A1(n_8358),
.A2(n_7456),
.B(n_7447),
.Y(n_9590)
);

INVx2_ASAP7_75t_SL g9591 ( 
.A(n_8166),
.Y(n_9591)
);

BUFx3_ASAP7_75t_L g9592 ( 
.A(n_8159),
.Y(n_9592)
);

INVx1_ASAP7_75t_L g9593 ( 
.A(n_8225),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_9479),
.Y(n_9594)
);

INVx2_ASAP7_75t_L g9595 ( 
.A(n_9479),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_8225),
.Y(n_9596)
);

AND2x2_ASAP7_75t_L g9597 ( 
.A(n_8177),
.B(n_7805),
.Y(n_9597)
);

BUFx2_ASAP7_75t_L g9598 ( 
.A(n_8177),
.Y(n_9598)
);

OR2x2_ASAP7_75t_L g9599 ( 
.A(n_8166),
.B(n_7367),
.Y(n_9599)
);

INVx1_ASAP7_75t_L g9600 ( 
.A(n_8228),
.Y(n_9600)
);

OAI222xp33_ASAP7_75t_L g9601 ( 
.A1(n_8304),
.A2(n_7517),
.B1(n_7462),
.B2(n_7646),
.C1(n_7082),
.C2(n_6923),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_9479),
.Y(n_9602)
);

INVx1_ASAP7_75t_L g9603 ( 
.A(n_8228),
.Y(n_9603)
);

INVx2_ASAP7_75t_L g9604 ( 
.A(n_9479),
.Y(n_9604)
);

OR2x6_ASAP7_75t_L g9605 ( 
.A(n_8199),
.B(n_6945),
.Y(n_9605)
);

AOI21x1_ASAP7_75t_L g9606 ( 
.A1(n_8161),
.A2(n_7966),
.B(n_7935),
.Y(n_9606)
);

HB1xp67_ASAP7_75t_L g9607 ( 
.A(n_8166),
.Y(n_9607)
);

CKINVDCx8_ASAP7_75t_R g9608 ( 
.A(n_8141),
.Y(n_9608)
);

INVx1_ASAP7_75t_L g9609 ( 
.A(n_8293),
.Y(n_9609)
);

INVx1_ASAP7_75t_L g9610 ( 
.A(n_8293),
.Y(n_9610)
);

INVx1_ASAP7_75t_L g9611 ( 
.A(n_8315),
.Y(n_9611)
);

INVx1_ASAP7_75t_L g9612 ( 
.A(n_8315),
.Y(n_9612)
);

AOI22xp33_ASAP7_75t_SL g9613 ( 
.A1(n_8853),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9613)
);

INVx1_ASAP7_75t_L g9614 ( 
.A(n_8321),
.Y(n_9614)
);

AOI22xp33_ASAP7_75t_L g9615 ( 
.A1(n_8271),
.A2(n_7712),
.B1(n_7710),
.B2(n_7650),
.Y(n_9615)
);

INVx3_ASAP7_75t_L g9616 ( 
.A(n_8191),
.Y(n_9616)
);

AOI21xp5_ASAP7_75t_L g9617 ( 
.A1(n_8195),
.A2(n_8075),
.B(n_7121),
.Y(n_9617)
);

HB1xp67_ASAP7_75t_L g9618 ( 
.A(n_9170),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_8321),
.Y(n_9619)
);

BUFx3_ASAP7_75t_L g9620 ( 
.A(n_8159),
.Y(n_9620)
);

CKINVDCx20_ASAP7_75t_R g9621 ( 
.A(n_8452),
.Y(n_9621)
);

INVx1_ASAP7_75t_L g9622 ( 
.A(n_8362),
.Y(n_9622)
);

INVx1_ASAP7_75t_L g9623 ( 
.A(n_8362),
.Y(n_9623)
);

INVx1_ASAP7_75t_L g9624 ( 
.A(n_8363),
.Y(n_9624)
);

AO21x1_ASAP7_75t_L g9625 ( 
.A1(n_8536),
.A2(n_7438),
.B(n_7363),
.Y(n_9625)
);

INVx4_ASAP7_75t_L g9626 ( 
.A(n_8159),
.Y(n_9626)
);

INVx2_ASAP7_75t_L g9627 ( 
.A(n_9479),
.Y(n_9627)
);

INVx1_ASAP7_75t_L g9628 ( 
.A(n_8363),
.Y(n_9628)
);

INVx2_ASAP7_75t_L g9629 ( 
.A(n_9479),
.Y(n_9629)
);

OAI21x1_ASAP7_75t_L g9630 ( 
.A1(n_8461),
.A2(n_6940),
.B(n_6924),
.Y(n_9630)
);

INVx2_ASAP7_75t_SL g9631 ( 
.A(n_8191),
.Y(n_9631)
);

INVxp67_ASAP7_75t_SL g9632 ( 
.A(n_8137),
.Y(n_9632)
);

INVx1_ASAP7_75t_L g9633 ( 
.A(n_8501),
.Y(n_9633)
);

HB1xp67_ASAP7_75t_L g9634 ( 
.A(n_9170),
.Y(n_9634)
);

INVx2_ASAP7_75t_L g9635 ( 
.A(n_9521),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_8501),
.Y(n_9636)
);

CKINVDCx5p33_ASAP7_75t_R g9637 ( 
.A(n_8747),
.Y(n_9637)
);

AOI22xp33_ASAP7_75t_L g9638 ( 
.A1(n_8222),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9638)
);

OAI21x1_ASAP7_75t_L g9639 ( 
.A1(n_8461),
.A2(n_6940),
.B(n_6924),
.Y(n_9639)
);

INVx1_ASAP7_75t_L g9640 ( 
.A(n_8516),
.Y(n_9640)
);

INVx1_ASAP7_75t_SL g9641 ( 
.A(n_9071),
.Y(n_9641)
);

INVx2_ASAP7_75t_L g9642 ( 
.A(n_9521),
.Y(n_9642)
);

BUFx2_ASAP7_75t_L g9643 ( 
.A(n_8191),
.Y(n_9643)
);

BUFx2_ASAP7_75t_L g9644 ( 
.A(n_8191),
.Y(n_9644)
);

INVx1_ASAP7_75t_SL g9645 ( 
.A(n_9142),
.Y(n_9645)
);

OA21x2_ASAP7_75t_L g9646 ( 
.A1(n_8243),
.A2(n_7353),
.B(n_7295),
.Y(n_9646)
);

INVx1_ASAP7_75t_L g9647 ( 
.A(n_8516),
.Y(n_9647)
);

AOI21xp5_ASAP7_75t_L g9648 ( 
.A1(n_8195),
.A2(n_7121),
.B(n_7969),
.Y(n_9648)
);

OA21x2_ASAP7_75t_L g9649 ( 
.A1(n_8243),
.A2(n_7405),
.B(n_7377),
.Y(n_9649)
);

AOI21x1_ASAP7_75t_L g9650 ( 
.A1(n_8161),
.A2(n_7966),
.B(n_7266),
.Y(n_9650)
);

AND2x2_ASAP7_75t_L g9651 ( 
.A(n_8158),
.B(n_7805),
.Y(n_9651)
);

AOI22xp5_ASAP7_75t_L g9652 ( 
.A1(n_8129),
.A2(n_8106),
.B1(n_8046),
.B2(n_7314),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_9521),
.Y(n_9653)
);

AOI21x1_ASAP7_75t_L g9654 ( 
.A1(n_8285),
.A2(n_8536),
.B(n_8358),
.Y(n_9654)
);

OAI21x1_ASAP7_75t_L g9655 ( 
.A1(n_8461),
.A2(n_7820),
.B(n_6940),
.Y(n_9655)
);

OA21x2_ASAP7_75t_L g9656 ( 
.A1(n_8243),
.A2(n_7405),
.B(n_7820),
.Y(n_9656)
);

BUFx12f_ASAP7_75t_L g9657 ( 
.A(n_8159),
.Y(n_9657)
);

INVxp67_ASAP7_75t_SL g9658 ( 
.A(n_8137),
.Y(n_9658)
);

AOI22xp33_ASAP7_75t_L g9659 ( 
.A1(n_8222),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9659)
);

AOI22xp33_ASAP7_75t_L g9660 ( 
.A1(n_9059),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_8553),
.Y(n_9661)
);

INVx1_ASAP7_75t_L g9662 ( 
.A(n_8553),
.Y(n_9662)
);

INVx2_ASAP7_75t_L g9663 ( 
.A(n_9521),
.Y(n_9663)
);

INVx2_ASAP7_75t_SL g9664 ( 
.A(n_8441),
.Y(n_9664)
);

BUFx12f_ASAP7_75t_L g9665 ( 
.A(n_8160),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8557),
.Y(n_9666)
);

INVx1_ASAP7_75t_L g9667 ( 
.A(n_8557),
.Y(n_9667)
);

BUFx2_ASAP7_75t_L g9668 ( 
.A(n_8158),
.Y(n_9668)
);

BUFx2_ASAP7_75t_L g9669 ( 
.A(n_8158),
.Y(n_9669)
);

INVx3_ASAP7_75t_L g9670 ( 
.A(n_8886),
.Y(n_9670)
);

INVx2_ASAP7_75t_SL g9671 ( 
.A(n_8441),
.Y(n_9671)
);

AND2x2_ASAP7_75t_L g9672 ( 
.A(n_8158),
.B(n_7805),
.Y(n_9672)
);

INVx1_ASAP7_75t_L g9673 ( 
.A(n_8562),
.Y(n_9673)
);

OAI22xp5_ASAP7_75t_L g9674 ( 
.A1(n_8304),
.A2(n_7305),
.B1(n_7825),
.B2(n_7936),
.Y(n_9674)
);

BUFx2_ASAP7_75t_L g9675 ( 
.A(n_8158),
.Y(n_9675)
);

CKINVDCx20_ASAP7_75t_R g9676 ( 
.A(n_8452),
.Y(n_9676)
);

AO21x1_ASAP7_75t_L g9677 ( 
.A1(n_8757),
.A2(n_8475),
.B(n_8148),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_9521),
.Y(n_9678)
);

INVx2_ASAP7_75t_L g9679 ( 
.A(n_9521),
.Y(n_9679)
);

AOI22xp33_ASAP7_75t_L g9680 ( 
.A1(n_9059),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9680)
);

BUFx3_ASAP7_75t_L g9681 ( 
.A(n_8160),
.Y(n_9681)
);

INVx1_ASAP7_75t_L g9682 ( 
.A(n_8562),
.Y(n_9682)
);

AOI22xp33_ASAP7_75t_L g9683 ( 
.A1(n_8565),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9683)
);

INVx1_ASAP7_75t_L g9684 ( 
.A(n_8638),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9524),
.Y(n_9685)
);

INVx1_ASAP7_75t_L g9686 ( 
.A(n_8638),
.Y(n_9686)
);

AND2x4_ASAP7_75t_L g9687 ( 
.A(n_8319),
.B(n_7810),
.Y(n_9687)
);

NAND2xp5_ASAP7_75t_L g9688 ( 
.A(n_8475),
.B(n_7281),
.Y(n_9688)
);

HB1xp67_ASAP7_75t_L g9689 ( 
.A(n_9170),
.Y(n_9689)
);

HB1xp67_ASAP7_75t_L g9690 ( 
.A(n_9172),
.Y(n_9690)
);

AOI22xp33_ASAP7_75t_SL g9691 ( 
.A1(n_8853),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9691)
);

AOI22xp33_ASAP7_75t_L g9692 ( 
.A1(n_8565),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9692)
);

OAI21x1_ASAP7_75t_L g9693 ( 
.A1(n_8219),
.A2(n_6940),
.B(n_6924),
.Y(n_9693)
);

INVx1_ASAP7_75t_SL g9694 ( 
.A(n_9142),
.Y(n_9694)
);

CKINVDCx6p67_ASAP7_75t_R g9695 ( 
.A(n_8160),
.Y(n_9695)
);

CKINVDCx11_ASAP7_75t_R g9696 ( 
.A(n_8200),
.Y(n_9696)
);

CKINVDCx11_ASAP7_75t_R g9697 ( 
.A(n_8200),
.Y(n_9697)
);

INVx1_ASAP7_75t_L g9698 ( 
.A(n_8645),
.Y(n_9698)
);

AOI21xp5_ASAP7_75t_L g9699 ( 
.A1(n_8526),
.A2(n_7121),
.B(n_7969),
.Y(n_9699)
);

INVx2_ASAP7_75t_L g9700 ( 
.A(n_9524),
.Y(n_9700)
);

OAI21x1_ASAP7_75t_L g9701 ( 
.A1(n_8199),
.A2(n_6940),
.B(n_6924),
.Y(n_9701)
);

AND2x4_ASAP7_75t_SL g9702 ( 
.A(n_8441),
.B(n_7840),
.Y(n_9702)
);

INVx3_ASAP7_75t_SL g9703 ( 
.A(n_8141),
.Y(n_9703)
);

INVx2_ASAP7_75t_L g9704 ( 
.A(n_9524),
.Y(n_9704)
);

OR2x2_ASAP7_75t_L g9705 ( 
.A(n_8218),
.B(n_7367),
.Y(n_9705)
);

CKINVDCx20_ASAP7_75t_R g9706 ( 
.A(n_8517),
.Y(n_9706)
);

INVx1_ASAP7_75t_L g9707 ( 
.A(n_8645),
.Y(n_9707)
);

BUFx6f_ASAP7_75t_L g9708 ( 
.A(n_8160),
.Y(n_9708)
);

INVx1_ASAP7_75t_SL g9709 ( 
.A(n_9436),
.Y(n_9709)
);

CKINVDCx5p33_ASAP7_75t_R g9710 ( 
.A(n_8747),
.Y(n_9710)
);

INVx1_ASAP7_75t_L g9711 ( 
.A(n_8646),
.Y(n_9711)
);

INVx2_ASAP7_75t_L g9712 ( 
.A(n_9524),
.Y(n_9712)
);

INVx2_ASAP7_75t_SL g9713 ( 
.A(n_8441),
.Y(n_9713)
);

INVx1_ASAP7_75t_L g9714 ( 
.A(n_8646),
.Y(n_9714)
);

HB1xp67_ASAP7_75t_L g9715 ( 
.A(n_9172),
.Y(n_9715)
);

OAI21x1_ASAP7_75t_L g9716 ( 
.A1(n_8219),
.A2(n_6940),
.B(n_6924),
.Y(n_9716)
);

BUFx3_ASAP7_75t_L g9717 ( 
.A(n_8180),
.Y(n_9717)
);

OAI21xp5_ASAP7_75t_L g9718 ( 
.A1(n_8129),
.A2(n_7308),
.B(n_7281),
.Y(n_9718)
);

BUFx2_ASAP7_75t_L g9719 ( 
.A(n_8170),
.Y(n_9719)
);

AOI22xp33_ASAP7_75t_L g9720 ( 
.A1(n_8133),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9720)
);

NOR2xp33_ASAP7_75t_L g9721 ( 
.A(n_8524),
.B(n_7545),
.Y(n_9721)
);

INVx3_ASAP7_75t_L g9722 ( 
.A(n_8886),
.Y(n_9722)
);

INVx1_ASAP7_75t_L g9723 ( 
.A(n_8808),
.Y(n_9723)
);

INVx2_ASAP7_75t_SL g9724 ( 
.A(n_8441),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_9524),
.Y(n_9725)
);

OA21x2_ASAP7_75t_L g9726 ( 
.A1(n_8224),
.A2(n_7456),
.B(n_7447),
.Y(n_9726)
);

AOI21x1_ASAP7_75t_L g9727 ( 
.A1(n_8285),
.A2(n_7266),
.B(n_7262),
.Y(n_9727)
);

INVx1_ASAP7_75t_L g9728 ( 
.A(n_8808),
.Y(n_9728)
);

INVx1_ASAP7_75t_SL g9729 ( 
.A(n_9436),
.Y(n_9729)
);

AOI22xp33_ASAP7_75t_L g9730 ( 
.A1(n_8133),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9730)
);

INVx2_ASAP7_75t_L g9731 ( 
.A(n_9524),
.Y(n_9731)
);

HB1xp67_ASAP7_75t_L g9732 ( 
.A(n_9172),
.Y(n_9732)
);

AOI22xp33_ASAP7_75t_L g9733 ( 
.A1(n_8325),
.A2(n_7650),
.B1(n_7743),
.B2(n_7736),
.Y(n_9733)
);

HB1xp67_ASAP7_75t_L g9734 ( 
.A(n_8170),
.Y(n_9734)
);

BUFx2_ASAP7_75t_R g9735 ( 
.A(n_8845),
.Y(n_9735)
);

BUFx3_ASAP7_75t_L g9736 ( 
.A(n_8180),
.Y(n_9736)
);

INVx2_ASAP7_75t_L g9737 ( 
.A(n_9545),
.Y(n_9737)
);

INVx1_ASAP7_75t_L g9738 ( 
.A(n_8809),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_8809),
.Y(n_9739)
);

INVx1_ASAP7_75t_L g9740 ( 
.A(n_8810),
.Y(n_9740)
);

INVx1_ASAP7_75t_L g9741 ( 
.A(n_8810),
.Y(n_9741)
);

OAI22xp33_ASAP7_75t_R g9742 ( 
.A1(n_8148),
.A2(n_7316),
.B1(n_7119),
.B2(n_7084),
.Y(n_9742)
);

BUFx4f_ASAP7_75t_SL g9743 ( 
.A(n_8180),
.Y(n_9743)
);

AOI22xp33_ASAP7_75t_SL g9744 ( 
.A1(n_8853),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_8811),
.Y(n_9745)
);

AND2x2_ASAP7_75t_L g9746 ( 
.A(n_8843),
.B(n_7810),
.Y(n_9746)
);

INVx2_ASAP7_75t_SL g9747 ( 
.A(n_9004),
.Y(n_9747)
);

AOI22xp33_ASAP7_75t_L g9748 ( 
.A1(n_8325),
.A2(n_7650),
.B1(n_7756),
.B2(n_7743),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_8811),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_8816),
.Y(n_9750)
);

INVx2_ASAP7_75t_L g9751 ( 
.A(n_9545),
.Y(n_9751)
);

INVx1_ASAP7_75t_L g9752 ( 
.A(n_8816),
.Y(n_9752)
);

INVx1_ASAP7_75t_L g9753 ( 
.A(n_8821),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_8821),
.Y(n_9754)
);

INVx2_ASAP7_75t_L g9755 ( 
.A(n_9545),
.Y(n_9755)
);

INVx1_ASAP7_75t_L g9756 ( 
.A(n_8840),
.Y(n_9756)
);

AND2x2_ASAP7_75t_L g9757 ( 
.A(n_8843),
.B(n_8875),
.Y(n_9757)
);

BUFx2_ASAP7_75t_L g9758 ( 
.A(n_9395),
.Y(n_9758)
);

INVx5_ASAP7_75t_L g9759 ( 
.A(n_8784),
.Y(n_9759)
);

OAI22xp5_ASAP7_75t_L g9760 ( 
.A1(n_8162),
.A2(n_7305),
.B1(n_7825),
.B2(n_7936),
.Y(n_9760)
);

AOI22xp33_ASAP7_75t_SL g9761 ( 
.A1(n_8867),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_8840),
.Y(n_9762)
);

INVx1_ASAP7_75t_L g9763 ( 
.A(n_8852),
.Y(n_9763)
);

BUFx6f_ASAP7_75t_L g9764 ( 
.A(n_8180),
.Y(n_9764)
);

BUFx2_ASAP7_75t_R g9765 ( 
.A(n_8845),
.Y(n_9765)
);

INVx3_ASAP7_75t_L g9766 ( 
.A(n_8886),
.Y(n_9766)
);

CKINVDCx20_ASAP7_75t_R g9767 ( 
.A(n_8517),
.Y(n_9767)
);

INVx2_ASAP7_75t_L g9768 ( 
.A(n_9545),
.Y(n_9768)
);

AND2x4_ASAP7_75t_L g9769 ( 
.A(n_8319),
.B(n_7810),
.Y(n_9769)
);

AOI22xp33_ASAP7_75t_L g9770 ( 
.A1(n_8325),
.A2(n_7650),
.B1(n_7757),
.B2(n_7756),
.Y(n_9770)
);

AOI22xp33_ASAP7_75t_L g9771 ( 
.A1(n_8233),
.A2(n_7650),
.B1(n_7757),
.B2(n_7756),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_8852),
.Y(n_9772)
);

INVx1_ASAP7_75t_L g9773 ( 
.A(n_8882),
.Y(n_9773)
);

BUFx2_ASAP7_75t_SL g9774 ( 
.A(n_8200),
.Y(n_9774)
);

AOI22xp33_ASAP7_75t_L g9775 ( 
.A1(n_8233),
.A2(n_7650),
.B1(n_7757),
.B2(n_7756),
.Y(n_9775)
);

CKINVDCx11_ASAP7_75t_R g9776 ( 
.A(n_8443),
.Y(n_9776)
);

INVx2_ASAP7_75t_L g9777 ( 
.A(n_9545),
.Y(n_9777)
);

NAND2xp5_ASAP7_75t_L g9778 ( 
.A(n_8267),
.B(n_7308),
.Y(n_9778)
);

INVx2_ASAP7_75t_L g9779 ( 
.A(n_9545),
.Y(n_9779)
);

INVx1_ASAP7_75t_L g9780 ( 
.A(n_8882),
.Y(n_9780)
);

OAI22xp5_ASAP7_75t_L g9781 ( 
.A1(n_8162),
.A2(n_7305),
.B1(n_7825),
.B2(n_7936),
.Y(n_9781)
);

BUFx3_ASAP7_75t_L g9782 ( 
.A(n_8587),
.Y(n_9782)
);

INVx5_ASAP7_75t_L g9783 ( 
.A(n_8784),
.Y(n_9783)
);

INVx2_ASAP7_75t_L g9784 ( 
.A(n_8691),
.Y(n_9784)
);

AND2x2_ASAP7_75t_L g9785 ( 
.A(n_8843),
.B(n_7810),
.Y(n_9785)
);

AND2x2_ASAP7_75t_L g9786 ( 
.A(n_8875),
.B(n_7838),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_8885),
.Y(n_9787)
);

INVx2_ASAP7_75t_L g9788 ( 
.A(n_8691),
.Y(n_9788)
);

INVx2_ASAP7_75t_L g9789 ( 
.A(n_8691),
.Y(n_9789)
);

INVx1_ASAP7_75t_L g9790 ( 
.A(n_8885),
.Y(n_9790)
);

INVx1_ASAP7_75t_L g9791 ( 
.A(n_8887),
.Y(n_9791)
);

OAI21xp5_ASAP7_75t_L g9792 ( 
.A1(n_8757),
.A2(n_7428),
.B(n_7411),
.Y(n_9792)
);

INVx1_ASAP7_75t_L g9793 ( 
.A(n_8887),
.Y(n_9793)
);

AOI22xp33_ASAP7_75t_L g9794 ( 
.A1(n_8231),
.A2(n_7650),
.B1(n_7757),
.B2(n_7756),
.Y(n_9794)
);

AOI22xp33_ASAP7_75t_SL g9795 ( 
.A1(n_8867),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_8896),
.Y(n_9796)
);

OAI22xp5_ASAP7_75t_L g9797 ( 
.A1(n_8418),
.A2(n_8637),
.B1(n_8194),
.B2(n_8284),
.Y(n_9797)
);

NAND2x1p5_ASAP7_75t_L g9798 ( 
.A(n_9141),
.B(n_8119),
.Y(n_9798)
);

BUFx8_ASAP7_75t_L g9799 ( 
.A(n_8587),
.Y(n_9799)
);

AOI22xp33_ASAP7_75t_L g9800 ( 
.A1(n_8231),
.A2(n_7757),
.B1(n_7779),
.B2(n_7756),
.Y(n_9800)
);

INVx1_ASAP7_75t_L g9801 ( 
.A(n_8896),
.Y(n_9801)
);

HB1xp67_ASAP7_75t_L g9802 ( 
.A(n_9270),
.Y(n_9802)
);

AOI22xp33_ASAP7_75t_L g9803 ( 
.A1(n_8192),
.A2(n_8198),
.B1(n_8867),
.B2(n_8858),
.Y(n_9803)
);

CKINVDCx20_ASAP7_75t_R g9804 ( 
.A(n_8545),
.Y(n_9804)
);

AO21x2_ASAP7_75t_L g9805 ( 
.A1(n_8358),
.A2(n_8183),
.B(n_8130),
.Y(n_9805)
);

INVx3_ASAP7_75t_L g9806 ( 
.A(n_8886),
.Y(n_9806)
);

OAI21xp5_ASAP7_75t_L g9807 ( 
.A1(n_8316),
.A2(n_7428),
.B(n_7411),
.Y(n_9807)
);

INVx2_ASAP7_75t_L g9808 ( 
.A(n_8691),
.Y(n_9808)
);

OAI22xp5_ASAP7_75t_L g9809 ( 
.A1(n_8418),
.A2(n_8637),
.B1(n_8194),
.B2(n_8284),
.Y(n_9809)
);

OA21x2_ASAP7_75t_L g9810 ( 
.A1(n_8224),
.A2(n_7456),
.B(n_7447),
.Y(n_9810)
);

INVx1_ASAP7_75t_SL g9811 ( 
.A(n_9471),
.Y(n_9811)
);

INVx1_ASAP7_75t_L g9812 ( 
.A(n_8898),
.Y(n_9812)
);

AOI22xp33_ASAP7_75t_L g9813 ( 
.A1(n_8192),
.A2(n_7757),
.B1(n_7779),
.B2(n_7756),
.Y(n_9813)
);

AOI22xp33_ASAP7_75t_L g9814 ( 
.A1(n_8198),
.A2(n_7757),
.B1(n_7779),
.B2(n_7756),
.Y(n_9814)
);

NAND2xp5_ASAP7_75t_L g9815 ( 
.A(n_8267),
.B(n_7440),
.Y(n_9815)
);

INVx1_ASAP7_75t_L g9816 ( 
.A(n_8898),
.Y(n_9816)
);

OAI22xp5_ASAP7_75t_L g9817 ( 
.A1(n_8778),
.A2(n_7305),
.B1(n_7953),
.B2(n_7348),
.Y(n_9817)
);

AO21x1_ASAP7_75t_L g9818 ( 
.A1(n_8718),
.A2(n_7363),
.B(n_7343),
.Y(n_9818)
);

INVx1_ASAP7_75t_L g9819 ( 
.A(n_8899),
.Y(n_9819)
);

INVxp67_ASAP7_75t_L g9820 ( 
.A(n_8410),
.Y(n_9820)
);

BUFx8_ASAP7_75t_SL g9821 ( 
.A(n_8142),
.Y(n_9821)
);

OAI21xp33_ASAP7_75t_SL g9822 ( 
.A1(n_8175),
.A2(n_7846),
.B(n_7838),
.Y(n_9822)
);

BUFx12f_ASAP7_75t_L g9823 ( 
.A(n_8587),
.Y(n_9823)
);

HB1xp67_ASAP7_75t_L g9824 ( 
.A(n_9270),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_8899),
.Y(n_9825)
);

AOI21x1_ASAP7_75t_L g9826 ( 
.A1(n_8771),
.A2(n_8175),
.B(n_8906),
.Y(n_9826)
);

OA21x2_ASAP7_75t_L g9827 ( 
.A1(n_8224),
.A2(n_7009),
.B(n_7007),
.Y(n_9827)
);

BUFx3_ASAP7_75t_L g9828 ( 
.A(n_8587),
.Y(n_9828)
);

INVx2_ASAP7_75t_L g9829 ( 
.A(n_8691),
.Y(n_9829)
);

BUFx4f_ASAP7_75t_SL g9830 ( 
.A(n_8681),
.Y(n_9830)
);

HB1xp67_ASAP7_75t_L g9831 ( 
.A(n_9274),
.Y(n_9831)
);

AND2x2_ASAP7_75t_L g9832 ( 
.A(n_8875),
.B(n_7838),
.Y(n_9832)
);

BUFx3_ASAP7_75t_L g9833 ( 
.A(n_8598),
.Y(n_9833)
);

AO21x1_ASAP7_75t_SL g9834 ( 
.A1(n_8307),
.A2(n_7368),
.B(n_7367),
.Y(n_9834)
);

INVx3_ASAP7_75t_L g9835 ( 
.A(n_8886),
.Y(n_9835)
);

AND2x2_ASAP7_75t_L g9836 ( 
.A(n_8288),
.B(n_7838),
.Y(n_9836)
);

AND2x2_ASAP7_75t_L g9837 ( 
.A(n_8288),
.B(n_7846),
.Y(n_9837)
);

INVx1_ASAP7_75t_L g9838 ( 
.A(n_8915),
.Y(n_9838)
);

INVx3_ASAP7_75t_L g9839 ( 
.A(n_8886),
.Y(n_9839)
);

INVx2_ASAP7_75t_L g9840 ( 
.A(n_8691),
.Y(n_9840)
);

BUFx3_ASAP7_75t_L g9841 ( 
.A(n_8598),
.Y(n_9841)
);

CKINVDCx6p67_ASAP7_75t_R g9842 ( 
.A(n_8524),
.Y(n_9842)
);

INVx3_ASAP7_75t_L g9843 ( 
.A(n_8886),
.Y(n_9843)
);

INVx2_ASAP7_75t_L g9844 ( 
.A(n_8945),
.Y(n_9844)
);

BUFx2_ASAP7_75t_SL g9845 ( 
.A(n_8443),
.Y(n_9845)
);

BUFx3_ASAP7_75t_L g9846 ( 
.A(n_8598),
.Y(n_9846)
);

AOI22xp33_ASAP7_75t_SL g9847 ( 
.A1(n_8209),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9847)
);

AOI22xp33_ASAP7_75t_L g9848 ( 
.A1(n_8858),
.A2(n_7757),
.B1(n_7779),
.B2(n_7756),
.Y(n_9848)
);

CKINVDCx6p67_ASAP7_75t_R g9849 ( 
.A(n_8524),
.Y(n_9849)
);

INVx1_ASAP7_75t_L g9850 ( 
.A(n_8915),
.Y(n_9850)
);

OAI21x1_ASAP7_75t_L g9851 ( 
.A1(n_8219),
.A2(n_6953),
.B(n_6924),
.Y(n_9851)
);

INVx2_ASAP7_75t_SL g9852 ( 
.A(n_9004),
.Y(n_9852)
);

CKINVDCx6p67_ASAP7_75t_R g9853 ( 
.A(n_8524),
.Y(n_9853)
);

AOI21x1_ASAP7_75t_L g9854 ( 
.A1(n_8771),
.A2(n_7266),
.B(n_7262),
.Y(n_9854)
);

NAND2xp5_ASAP7_75t_L g9855 ( 
.A(n_9417),
.B(n_8888),
.Y(n_9855)
);

BUFx6f_ASAP7_75t_L g9856 ( 
.A(n_8784),
.Y(n_9856)
);

INVx3_ASAP7_75t_L g9857 ( 
.A(n_8886),
.Y(n_9857)
);

INVx1_ASAP7_75t_L g9858 ( 
.A(n_8927),
.Y(n_9858)
);

BUFx2_ASAP7_75t_R g9859 ( 
.A(n_8142),
.Y(n_9859)
);

INVx2_ASAP7_75t_SL g9860 ( 
.A(n_9004),
.Y(n_9860)
);

INVx2_ASAP7_75t_L g9861 ( 
.A(n_8945),
.Y(n_9861)
);

AOI21xp5_ASAP7_75t_L g9862 ( 
.A1(n_8526),
.A2(n_7969),
.B(n_7143),
.Y(n_9862)
);

AOI22xp33_ASAP7_75t_SL g9863 ( 
.A1(n_8217),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9863)
);

AOI22xp33_ASAP7_75t_L g9864 ( 
.A1(n_8207),
.A2(n_7757),
.B1(n_7779),
.B2(n_7756),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_8927),
.Y(n_9865)
);

INVx3_ASAP7_75t_L g9866 ( 
.A(n_9099),
.Y(n_9866)
);

INVxp33_ASAP7_75t_L g9867 ( 
.A(n_9356),
.Y(n_9867)
);

INVx1_ASAP7_75t_L g9868 ( 
.A(n_8928),
.Y(n_9868)
);

CKINVDCx20_ASAP7_75t_R g9869 ( 
.A(n_8545),
.Y(n_9869)
);

INVx2_ASAP7_75t_L g9870 ( 
.A(n_8945),
.Y(n_9870)
);

AO21x2_ASAP7_75t_L g9871 ( 
.A1(n_8183),
.A2(n_7009),
.B(n_7007),
.Y(n_9871)
);

INVx3_ASAP7_75t_L g9872 ( 
.A(n_9099),
.Y(n_9872)
);

INVx2_ASAP7_75t_L g9873 ( 
.A(n_8945),
.Y(n_9873)
);

AOI22xp33_ASAP7_75t_L g9874 ( 
.A1(n_8207),
.A2(n_7779),
.B1(n_7757),
.B2(n_7709),
.Y(n_9874)
);

INVx2_ASAP7_75t_L g9875 ( 
.A(n_8945),
.Y(n_9875)
);

AOI21x1_ASAP7_75t_L g9876 ( 
.A1(n_8906),
.A2(n_7309),
.B(n_7262),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_8928),
.Y(n_9877)
);

INVx1_ASAP7_75t_L g9878 ( 
.A(n_8937),
.Y(n_9878)
);

BUFx2_ASAP7_75t_L g9879 ( 
.A(n_9395),
.Y(n_9879)
);

AOI21x1_ASAP7_75t_L g9880 ( 
.A1(n_8906),
.A2(n_7335),
.B(n_7309),
.Y(n_9880)
);

INVx3_ASAP7_75t_L g9881 ( 
.A(n_9099),
.Y(n_9881)
);

OAI22xp5_ASAP7_75t_L g9882 ( 
.A1(n_8778),
.A2(n_8275),
.B1(n_8153),
.B2(n_8286),
.Y(n_9882)
);

AOI22xp33_ASAP7_75t_L g9883 ( 
.A1(n_8190),
.A2(n_7779),
.B1(n_7709),
.B2(n_7707),
.Y(n_9883)
);

AND2x2_ASAP7_75t_L g9884 ( 
.A(n_8288),
.B(n_7846),
.Y(n_9884)
);

INVx1_ASAP7_75t_L g9885 ( 
.A(n_8937),
.Y(n_9885)
);

BUFx3_ASAP7_75t_L g9886 ( 
.A(n_8598),
.Y(n_9886)
);

BUFx3_ASAP7_75t_L g9887 ( 
.A(n_8598),
.Y(n_9887)
);

INVx3_ASAP7_75t_L g9888 ( 
.A(n_8474),
.Y(n_9888)
);

CKINVDCx11_ASAP7_75t_R g9889 ( 
.A(n_8443),
.Y(n_9889)
);

AOI21x1_ASAP7_75t_L g9890 ( 
.A1(n_9378),
.A2(n_7335),
.B(n_7309),
.Y(n_9890)
);

INVx1_ASAP7_75t_SL g9891 ( 
.A(n_9471),
.Y(n_9891)
);

INVx1_ASAP7_75t_L g9892 ( 
.A(n_8941),
.Y(n_9892)
);

HB1xp67_ASAP7_75t_L g9893 ( 
.A(n_9274),
.Y(n_9893)
);

BUFx6f_ASAP7_75t_L g9894 ( 
.A(n_8784),
.Y(n_9894)
);

INVx2_ASAP7_75t_L g9895 ( 
.A(n_8945),
.Y(n_9895)
);

OAI21x1_ASAP7_75t_SL g9896 ( 
.A1(n_8372),
.A2(n_7032),
.B(n_6935),
.Y(n_9896)
);

OAI22xp5_ASAP7_75t_L g9897 ( 
.A1(n_8275),
.A2(n_7305),
.B1(n_7953),
.B2(n_7348),
.Y(n_9897)
);

OAI22xp33_ASAP7_75t_R g9898 ( 
.A1(n_8439),
.A2(n_7316),
.B1(n_7084),
.B2(n_7111),
.Y(n_9898)
);

AO21x1_ASAP7_75t_L g9899 ( 
.A1(n_8718),
.A2(n_7363),
.B(n_7343),
.Y(n_9899)
);

BUFx3_ASAP7_75t_L g9900 ( 
.A(n_8598),
.Y(n_9900)
);

INVx2_ASAP7_75t_L g9901 ( 
.A(n_9256),
.Y(n_9901)
);

INVx1_ASAP7_75t_L g9902 ( 
.A(n_8941),
.Y(n_9902)
);

AOI22xp33_ASAP7_75t_L g9903 ( 
.A1(n_8190),
.A2(n_8957),
.B1(n_8838),
.B2(n_8846),
.Y(n_9903)
);

AND2x2_ASAP7_75t_L g9904 ( 
.A(n_8152),
.B(n_7846),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_8950),
.Y(n_9905)
);

INVx2_ASAP7_75t_L g9906 ( 
.A(n_9256),
.Y(n_9906)
);

INVx1_ASAP7_75t_L g9907 ( 
.A(n_8950),
.Y(n_9907)
);

INVx2_ASAP7_75t_L g9908 ( 
.A(n_9256),
.Y(n_9908)
);

INVx1_ASAP7_75t_SL g9909 ( 
.A(n_8878),
.Y(n_9909)
);

CKINVDCx20_ASAP7_75t_R g9910 ( 
.A(n_8878),
.Y(n_9910)
);

BUFx6f_ASAP7_75t_L g9911 ( 
.A(n_8596),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_8953),
.Y(n_9912)
);

NAND2x1p5_ASAP7_75t_L g9913 ( 
.A(n_9141),
.B(n_8119),
.Y(n_9913)
);

INVx11_ASAP7_75t_L g9914 ( 
.A(n_8681),
.Y(n_9914)
);

HB1xp67_ASAP7_75t_L g9915 ( 
.A(n_9279),
.Y(n_9915)
);

BUFx2_ASAP7_75t_L g9916 ( 
.A(n_8152),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_8953),
.Y(n_9917)
);

BUFx6f_ASAP7_75t_L g9918 ( 
.A(n_8596),
.Y(n_9918)
);

INVx2_ASAP7_75t_L g9919 ( 
.A(n_9256),
.Y(n_9919)
);

INVx2_ASAP7_75t_L g9920 ( 
.A(n_9256),
.Y(n_9920)
);

INVx1_ASAP7_75t_L g9921 ( 
.A(n_8958),
.Y(n_9921)
);

AOI22xp33_ASAP7_75t_SL g9922 ( 
.A1(n_8209),
.A2(n_8263),
.B1(n_8310),
.B2(n_8217),
.Y(n_9922)
);

AOI21x1_ASAP7_75t_L g9923 ( 
.A1(n_9378),
.A2(n_9202),
.B(n_8558),
.Y(n_9923)
);

INVx2_ASAP7_75t_L g9924 ( 
.A(n_9256),
.Y(n_9924)
);

NAND2x1p5_ASAP7_75t_L g9925 ( 
.A(n_9141),
.B(n_8119),
.Y(n_9925)
);

INVx2_ASAP7_75t_SL g9926 ( 
.A(n_9004),
.Y(n_9926)
);

INVx2_ASAP7_75t_L g9927 ( 
.A(n_9264),
.Y(n_9927)
);

AOI22xp33_ASAP7_75t_L g9928 ( 
.A1(n_8957),
.A2(n_7779),
.B1(n_7707),
.B2(n_7147),
.Y(n_9928)
);

INVx1_ASAP7_75t_L g9929 ( 
.A(n_8958),
.Y(n_9929)
);

AOI22xp33_ASAP7_75t_L g9930 ( 
.A1(n_8838),
.A2(n_7779),
.B1(n_7124),
.B2(n_7891),
.Y(n_9930)
);

AOI22xp33_ASAP7_75t_L g9931 ( 
.A1(n_8846),
.A2(n_7779),
.B1(n_7488),
.B2(n_7272),
.Y(n_9931)
);

BUFx8_ASAP7_75t_L g9932 ( 
.A(n_8681),
.Y(n_9932)
);

INVx2_ASAP7_75t_L g9933 ( 
.A(n_9264),
.Y(n_9933)
);

BUFx2_ASAP7_75t_SL g9934 ( 
.A(n_8947),
.Y(n_9934)
);

INVx4_ASAP7_75t_L g9935 ( 
.A(n_8671),
.Y(n_9935)
);

AND2x2_ASAP7_75t_L g9936 ( 
.A(n_8152),
.B(n_7854),
.Y(n_9936)
);

AOI22xp33_ASAP7_75t_L g9937 ( 
.A1(n_8196),
.A2(n_7488),
.B1(n_7272),
.B2(n_7277),
.Y(n_9937)
);

INVx1_ASAP7_75t_L g9938 ( 
.A(n_8960),
.Y(n_9938)
);

NAND2xp5_ASAP7_75t_L g9939 ( 
.A(n_9417),
.B(n_7440),
.Y(n_9939)
);

INVx2_ASAP7_75t_L g9940 ( 
.A(n_9264),
.Y(n_9940)
);

AOI22xp33_ASAP7_75t_SL g9941 ( 
.A1(n_8209),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_9941)
);

INVx1_ASAP7_75t_L g9942 ( 
.A(n_8960),
.Y(n_9942)
);

INVx1_ASAP7_75t_L g9943 ( 
.A(n_8965),
.Y(n_9943)
);

INVx1_ASAP7_75t_L g9944 ( 
.A(n_8965),
.Y(n_9944)
);

BUFx2_ASAP7_75t_SL g9945 ( 
.A(n_8947),
.Y(n_9945)
);

INVx2_ASAP7_75t_L g9946 ( 
.A(n_9264),
.Y(n_9946)
);

BUFx12f_ASAP7_75t_L g9947 ( 
.A(n_8535),
.Y(n_9947)
);

INVx2_ASAP7_75t_L g9948 ( 
.A(n_9264),
.Y(n_9948)
);

INVx3_ASAP7_75t_L g9949 ( 
.A(n_8474),
.Y(n_9949)
);

HB1xp67_ASAP7_75t_L g9950 ( 
.A(n_9279),
.Y(n_9950)
);

INVx2_ASAP7_75t_L g9951 ( 
.A(n_9264),
.Y(n_9951)
);

INVx1_ASAP7_75t_L g9952 ( 
.A(n_9248),
.Y(n_9952)
);

INVx6_ASAP7_75t_L g9953 ( 
.A(n_8879),
.Y(n_9953)
);

INVx6_ASAP7_75t_L g9954 ( 
.A(n_8879),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_9248),
.Y(n_9955)
);

BUFx2_ASAP7_75t_L g9956 ( 
.A(n_8176),
.Y(n_9956)
);

INVx2_ASAP7_75t_L g9957 ( 
.A(n_9295),
.Y(n_9957)
);

OAI21x1_ASAP7_75t_L g9958 ( 
.A1(n_8396),
.A2(n_8210),
.B(n_8527),
.Y(n_9958)
);

INVx2_ASAP7_75t_SL g9959 ( 
.A(n_9004),
.Y(n_9959)
);

INVx3_ASAP7_75t_L g9960 ( 
.A(n_8474),
.Y(n_9960)
);

INVx2_ASAP7_75t_L g9961 ( 
.A(n_9295),
.Y(n_9961)
);

INVx1_ASAP7_75t_L g9962 ( 
.A(n_9254),
.Y(n_9962)
);

INVx2_ASAP7_75t_SL g9963 ( 
.A(n_9440),
.Y(n_9963)
);

INVx1_ASAP7_75t_L g9964 ( 
.A(n_9254),
.Y(n_9964)
);

AND2x2_ASAP7_75t_L g9965 ( 
.A(n_8176),
.B(n_7854),
.Y(n_9965)
);

AOI22xp33_ASAP7_75t_L g9966 ( 
.A1(n_8196),
.A2(n_7277),
.B1(n_7313),
.B2(n_7263),
.Y(n_9966)
);

NAND2xp5_ASAP7_75t_L g9967 ( 
.A(n_9417),
.B(n_7343),
.Y(n_9967)
);

OR2x2_ASAP7_75t_L g9968 ( 
.A(n_8218),
.B(n_7368),
.Y(n_9968)
);

BUFx2_ASAP7_75t_R g9969 ( 
.A(n_8535),
.Y(n_9969)
);

INVx6_ASAP7_75t_L g9970 ( 
.A(n_8879),
.Y(n_9970)
);

INVx2_ASAP7_75t_L g9971 ( 
.A(n_9295),
.Y(n_9971)
);

BUFx3_ASAP7_75t_L g9972 ( 
.A(n_8681),
.Y(n_9972)
);

NAND2xp5_ASAP7_75t_L g9973 ( 
.A(n_9417),
.B(n_7368),
.Y(n_9973)
);

AOI22xp33_ASAP7_75t_L g9974 ( 
.A1(n_8130),
.A2(n_8241),
.B1(n_8153),
.B2(n_9478),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_9338),
.Y(n_9975)
);

INVx2_ASAP7_75t_L g9976 ( 
.A(n_9295),
.Y(n_9976)
);

AND2x2_ASAP7_75t_L g9977 ( 
.A(n_8176),
.B(n_7854),
.Y(n_9977)
);

INVx1_ASAP7_75t_L g9978 ( 
.A(n_9338),
.Y(n_9978)
);

AOI22xp33_ASAP7_75t_L g9979 ( 
.A1(n_8241),
.A2(n_7313),
.B1(n_7263),
.B2(n_6923),
.Y(n_9979)
);

INVx2_ASAP7_75t_L g9980 ( 
.A(n_9295),
.Y(n_9980)
);

INVx1_ASAP7_75t_L g9981 ( 
.A(n_9379),
.Y(n_9981)
);

INVx1_ASAP7_75t_SL g9982 ( 
.A(n_9278),
.Y(n_9982)
);

HB1xp67_ASAP7_75t_L g9983 ( 
.A(n_9312),
.Y(n_9983)
);

AOI22xp33_ASAP7_75t_L g9984 ( 
.A1(n_9478),
.A2(n_6923),
.B1(n_7517),
.B2(n_7462),
.Y(n_9984)
);

AOI22xp33_ASAP7_75t_L g9985 ( 
.A1(n_8181),
.A2(n_7517),
.B1(n_7067),
.B2(n_7064),
.Y(n_9985)
);

NAND2xp5_ASAP7_75t_L g9986 ( 
.A(n_9417),
.B(n_6974),
.Y(n_9986)
);

INVx2_ASAP7_75t_L g9987 ( 
.A(n_9295),
.Y(n_9987)
);

NAND2x1p5_ASAP7_75t_L g9988 ( 
.A(n_9141),
.B(n_8119),
.Y(n_9988)
);

INVx1_ASAP7_75t_L g9989 ( 
.A(n_9379),
.Y(n_9989)
);

BUFx3_ASAP7_75t_L g9990 ( 
.A(n_8759),
.Y(n_9990)
);

OA21x2_ASAP7_75t_L g9991 ( 
.A1(n_8396),
.A2(n_7009),
.B(n_7007),
.Y(n_9991)
);

BUFx8_ASAP7_75t_L g9992 ( 
.A(n_8759),
.Y(n_9992)
);

OAI22xp5_ASAP7_75t_L g9993 ( 
.A1(n_8286),
.A2(n_7953),
.B1(n_7291),
.B2(n_7482),
.Y(n_9993)
);

INVx3_ASAP7_75t_L g9994 ( 
.A(n_8474),
.Y(n_9994)
);

OAI22xp33_ASAP7_75t_L g9995 ( 
.A1(n_9288),
.A2(n_7646),
.B1(n_7135),
.B2(n_7452),
.Y(n_9995)
);

NAND2xp5_ASAP7_75t_L g9996 ( 
.A(n_8888),
.B(n_6974),
.Y(n_9996)
);

BUFx4f_ASAP7_75t_SL g9997 ( 
.A(n_8759),
.Y(n_9997)
);

AO21x1_ASAP7_75t_SL g9998 ( 
.A1(n_8307),
.A2(n_7324),
.B(n_7320),
.Y(n_9998)
);

INVx6_ASAP7_75t_L g9999 ( 
.A(n_8879),
.Y(n_9999)
);

INVx1_ASAP7_75t_L g10000 ( 
.A(n_9381),
.Y(n_10000)
);

OR2x6_ASAP7_75t_L g10001 ( 
.A(n_8251),
.B(n_6945),
.Y(n_10001)
);

CKINVDCx20_ASAP7_75t_R g10002 ( 
.A(n_9278),
.Y(n_10002)
);

AOI22xp33_ASAP7_75t_L g10003 ( 
.A1(n_8181),
.A2(n_7067),
.B1(n_7064),
.B2(n_7108),
.Y(n_10003)
);

NAND2xp5_ASAP7_75t_L g10004 ( 
.A(n_8888),
.B(n_6974),
.Y(n_10004)
);

AOI22xp33_ASAP7_75t_SL g10005 ( 
.A1(n_8217),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_10005)
);

INVx2_ASAP7_75t_L g10006 ( 
.A(n_9316),
.Y(n_10006)
);

INVx1_ASAP7_75t_L g10007 ( 
.A(n_9381),
.Y(n_10007)
);

AOI22xp33_ASAP7_75t_L g10008 ( 
.A1(n_8229),
.A2(n_7113),
.B1(n_7108),
.B2(n_7195),
.Y(n_10008)
);

BUFx3_ASAP7_75t_L g10009 ( 
.A(n_8759),
.Y(n_10009)
);

INVx1_ASAP7_75t_L g10010 ( 
.A(n_9388),
.Y(n_10010)
);

AND2x4_ASAP7_75t_L g10011 ( 
.A(n_8262),
.B(n_7854),
.Y(n_10011)
);

INVx6_ASAP7_75t_L g10012 ( 
.A(n_8879),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_9388),
.Y(n_10013)
);

INVx1_ASAP7_75t_L g10014 ( 
.A(n_9391),
.Y(n_10014)
);

AND2x4_ASAP7_75t_L g10015 ( 
.A(n_8262),
.B(n_7857),
.Y(n_10015)
);

INVx2_ASAP7_75t_L g10016 ( 
.A(n_9316),
.Y(n_10016)
);

AND2x2_ASAP7_75t_L g10017 ( 
.A(n_8830),
.B(n_7857),
.Y(n_10017)
);

INVx4_ASAP7_75t_L g10018 ( 
.A(n_8671),
.Y(n_10018)
);

INVx2_ASAP7_75t_L g10019 ( 
.A(n_9316),
.Y(n_10019)
);

AO21x2_ASAP7_75t_L g10020 ( 
.A1(n_8183),
.A2(n_7314),
.B(n_7489),
.Y(n_10020)
);

INVx2_ASAP7_75t_L g10021 ( 
.A(n_9316),
.Y(n_10021)
);

INVx1_ASAP7_75t_L g10022 ( 
.A(n_9391),
.Y(n_10022)
);

AND2x4_ASAP7_75t_L g10023 ( 
.A(n_8318),
.B(n_7857),
.Y(n_10023)
);

OAI22x1_ASAP7_75t_L g10024 ( 
.A1(n_9332),
.A2(n_7043),
.B1(n_7452),
.B2(n_7203),
.Y(n_10024)
);

INVx2_ASAP7_75t_L g10025 ( 
.A(n_9316),
.Y(n_10025)
);

AOI21x1_ASAP7_75t_L g10026 ( 
.A1(n_9202),
.A2(n_7346),
.B(n_7335),
.Y(n_10026)
);

OAI22xp5_ASAP7_75t_L g10027 ( 
.A1(n_8229),
.A2(n_7291),
.B1(n_7482),
.B2(n_7348),
.Y(n_10027)
);

BUFx8_ASAP7_75t_L g10028 ( 
.A(n_8766),
.Y(n_10028)
);

CKINVDCx11_ASAP7_75t_R g10029 ( 
.A(n_8947),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_9549),
.Y(n_10030)
);

INVx1_ASAP7_75t_L g10031 ( 
.A(n_9549),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_9554),
.Y(n_10032)
);

OAI21xp5_ASAP7_75t_L g10033 ( 
.A1(n_8316),
.A2(n_7858),
.B(n_7792),
.Y(n_10033)
);

OAI22xp5_ASAP7_75t_L g10034 ( 
.A1(n_8415),
.A2(n_7291),
.B1(n_7482),
.B2(n_7348),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_9316),
.Y(n_10035)
);

INVx2_ASAP7_75t_L g10036 ( 
.A(n_9362),
.Y(n_10036)
);

NAND2x1p5_ASAP7_75t_L g10037 ( 
.A(n_9141),
.B(n_8119),
.Y(n_10037)
);

CKINVDCx5p33_ASAP7_75t_R g10038 ( 
.A(n_9148),
.Y(n_10038)
);

CKINVDCx11_ASAP7_75t_R g10039 ( 
.A(n_9245),
.Y(n_10039)
);

AO21x1_ASAP7_75t_L g10040 ( 
.A1(n_9333),
.A2(n_7775),
.B(n_7772),
.Y(n_10040)
);

INVx1_ASAP7_75t_L g10041 ( 
.A(n_9554),
.Y(n_10041)
);

INVx2_ASAP7_75t_SL g10042 ( 
.A(n_9440),
.Y(n_10042)
);

BUFx8_ASAP7_75t_L g10043 ( 
.A(n_8766),
.Y(n_10043)
);

OAI21x1_ASAP7_75t_L g10044 ( 
.A1(n_8396),
.A2(n_6959),
.B(n_6953),
.Y(n_10044)
);

INVx2_ASAP7_75t_L g10045 ( 
.A(n_9362),
.Y(n_10045)
);

HB1xp67_ASAP7_75t_L g10046 ( 
.A(n_9312),
.Y(n_10046)
);

INVx2_ASAP7_75t_SL g10047 ( 
.A(n_9440),
.Y(n_10047)
);

INVx1_ASAP7_75t_L g10048 ( 
.A(n_9437),
.Y(n_10048)
);

INVx3_ASAP7_75t_L g10049 ( 
.A(n_8474),
.Y(n_10049)
);

INVxp67_ASAP7_75t_L g10050 ( 
.A(n_8410),
.Y(n_10050)
);

BUFx12f_ASAP7_75t_L g10051 ( 
.A(n_8651),
.Y(n_10051)
);

INVx3_ASAP7_75t_L g10052 ( 
.A(n_8474),
.Y(n_10052)
);

AOI21x1_ASAP7_75t_L g10053 ( 
.A1(n_9202),
.A2(n_8558),
.B(n_8242),
.Y(n_10053)
);

AND2x4_ASAP7_75t_L g10054 ( 
.A(n_8318),
.B(n_7857),
.Y(n_10054)
);

AOI22xp33_ASAP7_75t_L g10055 ( 
.A1(n_9220),
.A2(n_7113),
.B1(n_7200),
.B2(n_7195),
.Y(n_10055)
);

CKINVDCx5p33_ASAP7_75t_R g10056 ( 
.A(n_9148),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_9437),
.Y(n_10057)
);

AOI22xp33_ASAP7_75t_SL g10058 ( 
.A1(n_8310),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_10058)
);

CKINVDCx12_ASAP7_75t_R g10059 ( 
.A(n_8338),
.Y(n_10059)
);

AOI22xp33_ASAP7_75t_SL g10060 ( 
.A1(n_8310),
.A2(n_7126),
.B1(n_7231),
.B2(n_7172),
.Y(n_10060)
);

BUFx6f_ASAP7_75t_L g10061 ( 
.A(n_8596),
.Y(n_10061)
);

INVx2_ASAP7_75t_L g10062 ( 
.A(n_9362),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_9437),
.Y(n_10063)
);

INVx2_ASAP7_75t_L g10064 ( 
.A(n_9362),
.Y(n_10064)
);

AND2x2_ASAP7_75t_L g10065 ( 
.A(n_8830),
.B(n_7881),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9443),
.Y(n_10066)
);

INVx2_ASAP7_75t_L g10067 ( 
.A(n_9362),
.Y(n_10067)
);

AOI22xp33_ASAP7_75t_L g10068 ( 
.A1(n_9220),
.A2(n_7200),
.B1(n_7052),
.B2(n_6945),
.Y(n_10068)
);

AOI22xp33_ASAP7_75t_L g10069 ( 
.A1(n_9219),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10069)
);

INVx1_ASAP7_75t_L g10070 ( 
.A(n_9443),
.Y(n_10070)
);

AOI22xp33_ASAP7_75t_L g10071 ( 
.A1(n_9219),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10071)
);

CKINVDCx11_ASAP7_75t_R g10072 ( 
.A(n_9245),
.Y(n_10072)
);

INVx2_ASAP7_75t_L g10073 ( 
.A(n_9362),
.Y(n_10073)
);

INVx2_ASAP7_75t_L g10074 ( 
.A(n_9383),
.Y(n_10074)
);

AND2x2_ASAP7_75t_L g10075 ( 
.A(n_8830),
.B(n_7881),
.Y(n_10075)
);

INVx1_ASAP7_75t_L g10076 ( 
.A(n_9443),
.Y(n_10076)
);

INVx2_ASAP7_75t_L g10077 ( 
.A(n_9383),
.Y(n_10077)
);

INVx1_ASAP7_75t_L g10078 ( 
.A(n_9483),
.Y(n_10078)
);

INVx2_ASAP7_75t_L g10079 ( 
.A(n_9383),
.Y(n_10079)
);

CKINVDCx10_ASAP7_75t_R g10080 ( 
.A(n_9466),
.Y(n_10080)
);

BUFx3_ASAP7_75t_L g10081 ( 
.A(n_8766),
.Y(n_10081)
);

BUFx12f_ASAP7_75t_L g10082 ( 
.A(n_8651),
.Y(n_10082)
);

NOR2xp33_ASAP7_75t_L g10083 ( 
.A(n_8619),
.B(n_7545),
.Y(n_10083)
);

INVx1_ASAP7_75t_L g10084 ( 
.A(n_9483),
.Y(n_10084)
);

OR2x2_ASAP7_75t_L g10085 ( 
.A(n_8218),
.B(n_8174),
.Y(n_10085)
);

BUFx3_ASAP7_75t_L g10086 ( 
.A(n_8766),
.Y(n_10086)
);

INVx1_ASAP7_75t_L g10087 ( 
.A(n_9483),
.Y(n_10087)
);

INVx1_ASAP7_75t_L g10088 ( 
.A(n_9513),
.Y(n_10088)
);

AOI22xp33_ASAP7_75t_L g10089 ( 
.A1(n_8251),
.A2(n_9333),
.B1(n_8399),
.B2(n_9201),
.Y(n_10089)
);

AOI22xp5_ASAP7_75t_L g10090 ( 
.A1(n_8416),
.A2(n_7489),
.B1(n_8007),
.B2(n_7082),
.Y(n_10090)
);

INVx1_ASAP7_75t_L g10091 ( 
.A(n_9513),
.Y(n_10091)
);

INVx1_ASAP7_75t_L g10092 ( 
.A(n_9513),
.Y(n_10092)
);

BUFx12f_ASAP7_75t_L g10093 ( 
.A(n_8923),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_8139),
.Y(n_10094)
);

INVx4_ASAP7_75t_L g10095 ( 
.A(n_8619),
.Y(n_10095)
);

INVx2_ASAP7_75t_L g10096 ( 
.A(n_9383),
.Y(n_10096)
);

HB1xp67_ASAP7_75t_L g10097 ( 
.A(n_9312),
.Y(n_10097)
);

INVx1_ASAP7_75t_L g10098 ( 
.A(n_8139),
.Y(n_10098)
);

INVx2_ASAP7_75t_L g10099 ( 
.A(n_9383),
.Y(n_10099)
);

OR2x2_ASAP7_75t_L g10100 ( 
.A(n_8218),
.B(n_7194),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_8139),
.Y(n_10101)
);

BUFx12f_ASAP7_75t_L g10102 ( 
.A(n_8923),
.Y(n_10102)
);

OAI21x1_ASAP7_75t_L g10103 ( 
.A1(n_8210),
.A2(n_6959),
.B(n_6953),
.Y(n_10103)
);

INVx1_ASAP7_75t_L g10104 ( 
.A(n_8147),
.Y(n_10104)
);

AOI22xp33_ASAP7_75t_L g10105 ( 
.A1(n_8399),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10105)
);

AOI22xp33_ASAP7_75t_L g10106 ( 
.A1(n_9201),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10106)
);

INVx2_ASAP7_75t_SL g10107 ( 
.A(n_9440),
.Y(n_10107)
);

CKINVDCx16_ASAP7_75t_R g10108 ( 
.A(n_9466),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_8147),
.Y(n_10109)
);

OA21x2_ASAP7_75t_L g10110 ( 
.A1(n_8210),
.A2(n_8249),
.B(n_8527),
.Y(n_10110)
);

INVx2_ASAP7_75t_L g10111 ( 
.A(n_9383),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_8147),
.Y(n_10112)
);

BUFx2_ASAP7_75t_R g10113 ( 
.A(n_9021),
.Y(n_10113)
);

NAND2xp5_ASAP7_75t_L g10114 ( 
.A(n_9438),
.B(n_7772),
.Y(n_10114)
);

OAI21x1_ASAP7_75t_L g10115 ( 
.A1(n_8527),
.A2(n_6959),
.B(n_6953),
.Y(n_10115)
);

OAI21xp5_ASAP7_75t_L g10116 ( 
.A1(n_8327),
.A2(n_7858),
.B(n_7792),
.Y(n_10116)
);

AOI22xp33_ASAP7_75t_SL g10117 ( 
.A1(n_8263),
.A2(n_8404),
.B1(n_8636),
.B2(n_8635),
.Y(n_10117)
);

INVx2_ASAP7_75t_L g10118 ( 
.A(n_9402),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_8154),
.Y(n_10119)
);

INVx1_ASAP7_75t_L g10120 ( 
.A(n_8154),
.Y(n_10120)
);

OAI21x1_ASAP7_75t_L g10121 ( 
.A1(n_8789),
.A2(n_6959),
.B(n_6953),
.Y(n_10121)
);

INVx2_ASAP7_75t_L g10122 ( 
.A(n_9402),
.Y(n_10122)
);

INVx3_ASAP7_75t_L g10123 ( 
.A(n_9070),
.Y(n_10123)
);

INVx2_ASAP7_75t_L g10124 ( 
.A(n_9402),
.Y(n_10124)
);

AND2x4_ASAP7_75t_L g10125 ( 
.A(n_8372),
.B(n_7881),
.Y(n_10125)
);

AOI22xp33_ASAP7_75t_L g10126 ( 
.A1(n_9332),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10126)
);

INVx1_ASAP7_75t_L g10127 ( 
.A(n_8154),
.Y(n_10127)
);

INVx2_ASAP7_75t_L g10128 ( 
.A(n_9402),
.Y(n_10128)
);

OAI22xp5_ASAP7_75t_L g10129 ( 
.A1(n_8415),
.A2(n_7291),
.B1(n_7482),
.B2(n_7348),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_8169),
.Y(n_10130)
);

AOI22xp33_ASAP7_75t_L g10131 ( 
.A1(n_8263),
.A2(n_7052),
.B1(n_7298),
.B2(n_6945),
.Y(n_10131)
);

INVx2_ASAP7_75t_L g10132 ( 
.A(n_9402),
.Y(n_10132)
);

AOI22xp33_ASAP7_75t_SL g10133 ( 
.A1(n_8404),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10133)
);

AOI22xp33_ASAP7_75t_L g10134 ( 
.A1(n_8404),
.A2(n_7298),
.B1(n_7323),
.B2(n_7052),
.Y(n_10134)
);

HB1xp67_ASAP7_75t_L g10135 ( 
.A(n_9312),
.Y(n_10135)
);

INVx1_ASAP7_75t_L g10136 ( 
.A(n_8169),
.Y(n_10136)
);

BUFx6f_ASAP7_75t_L g10137 ( 
.A(n_8596),
.Y(n_10137)
);

INVx2_ASAP7_75t_L g10138 ( 
.A(n_9402),
.Y(n_10138)
);

OA21x2_ASAP7_75t_L g10139 ( 
.A1(n_8249),
.A2(n_7234),
.B(n_7192),
.Y(n_10139)
);

INVx2_ASAP7_75t_L g10140 ( 
.A(n_9458),
.Y(n_10140)
);

INVx2_ASAP7_75t_L g10141 ( 
.A(n_9458),
.Y(n_10141)
);

CKINVDCx11_ASAP7_75t_R g10142 ( 
.A(n_9245),
.Y(n_10142)
);

AOI21x1_ASAP7_75t_L g10143 ( 
.A1(n_8558),
.A2(n_7346),
.B(n_7403),
.Y(n_10143)
);

OAI21x1_ASAP7_75t_L g10144 ( 
.A1(n_8464),
.A2(n_6959),
.B(n_6953),
.Y(n_10144)
);

AOI22xp33_ASAP7_75t_SL g10145 ( 
.A1(n_8635),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10145)
);

INVx1_ASAP7_75t_L g10146 ( 
.A(n_8169),
.Y(n_10146)
);

BUFx2_ASAP7_75t_L g10147 ( 
.A(n_8218),
.Y(n_10147)
);

AOI22xp33_ASAP7_75t_L g10148 ( 
.A1(n_8635),
.A2(n_8636),
.B1(n_8795),
.B2(n_8749),
.Y(n_10148)
);

AOI22xp33_ASAP7_75t_SL g10149 ( 
.A1(n_8636),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10149)
);

AND2x2_ASAP7_75t_L g10150 ( 
.A(n_8525),
.B(n_7881),
.Y(n_10150)
);

CKINVDCx20_ASAP7_75t_R g10151 ( 
.A(n_9285),
.Y(n_10151)
);

BUFx6f_ASAP7_75t_L g10152 ( 
.A(n_8605),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_8184),
.Y(n_10153)
);

NAND2xp5_ASAP7_75t_L g10154 ( 
.A(n_9438),
.B(n_7772),
.Y(n_10154)
);

NOR2xp33_ASAP7_75t_L g10155 ( 
.A(n_8619),
.B(n_7370),
.Y(n_10155)
);

INVx1_ASAP7_75t_L g10156 ( 
.A(n_8184),
.Y(n_10156)
);

BUFx2_ASAP7_75t_L g10157 ( 
.A(n_8218),
.Y(n_10157)
);

OAI22xp33_ASAP7_75t_L g10158 ( 
.A1(n_9288),
.A2(n_7646),
.B1(n_7135),
.B2(n_7452),
.Y(n_10158)
);

OAI21x1_ASAP7_75t_SL g10159 ( 
.A1(n_8372),
.A2(n_7032),
.B(n_6935),
.Y(n_10159)
);

OAI21x1_ASAP7_75t_L g10160 ( 
.A1(n_8464),
.A2(n_6967),
.B(n_6959),
.Y(n_10160)
);

NAND2x1p5_ASAP7_75t_L g10161 ( 
.A(n_8507),
.B(n_7509),
.Y(n_10161)
);

AOI22xp33_ASAP7_75t_SL g10162 ( 
.A1(n_8795),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10162)
);

INVx2_ASAP7_75t_L g10163 ( 
.A(n_9458),
.Y(n_10163)
);

OR2x6_ASAP7_75t_L g10164 ( 
.A(n_8447),
.B(n_8408),
.Y(n_10164)
);

HB1xp67_ASAP7_75t_L g10165 ( 
.A(n_9312),
.Y(n_10165)
);

INVx1_ASAP7_75t_L g10166 ( 
.A(n_8184),
.Y(n_10166)
);

AOI22xp33_ASAP7_75t_L g10167 ( 
.A1(n_8749),
.A2(n_7298),
.B1(n_7323),
.B2(n_7052),
.Y(n_10167)
);

BUFx2_ASAP7_75t_R g10168 ( 
.A(n_9021),
.Y(n_10168)
);

INVx3_ASAP7_75t_L g10169 ( 
.A(n_9070),
.Y(n_10169)
);

INVx2_ASAP7_75t_L g10170 ( 
.A(n_9458),
.Y(n_10170)
);

BUFx2_ASAP7_75t_L g10171 ( 
.A(n_8218),
.Y(n_10171)
);

INVx1_ASAP7_75t_L g10172 ( 
.A(n_8193),
.Y(n_10172)
);

AOI21x1_ASAP7_75t_L g10173 ( 
.A1(n_8188),
.A2(n_7346),
.B(n_7403),
.Y(n_10173)
);

NAND2x1p5_ASAP7_75t_L g10174 ( 
.A(n_8507),
.B(n_7509),
.Y(n_10174)
);

CKINVDCx20_ASAP7_75t_R g10175 ( 
.A(n_9285),
.Y(n_10175)
);

INVx1_ASAP7_75t_L g10176 ( 
.A(n_8193),
.Y(n_10176)
);

INVx1_ASAP7_75t_L g10177 ( 
.A(n_8193),
.Y(n_10177)
);

AND2x2_ASAP7_75t_L g10178 ( 
.A(n_8525),
.B(n_7887),
.Y(n_10178)
);

AOI22xp33_ASAP7_75t_SL g10179 ( 
.A1(n_8749),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10179)
);

AND2x2_ASAP7_75t_L g10180 ( 
.A(n_8525),
.B(n_8538),
.Y(n_10180)
);

AOI22xp33_ASAP7_75t_L g10181 ( 
.A1(n_8795),
.A2(n_7323),
.B1(n_7298),
.B2(n_6927),
.Y(n_10181)
);

INVx2_ASAP7_75t_L g10182 ( 
.A(n_9458),
.Y(n_10182)
);

AND2x2_ASAP7_75t_L g10183 ( 
.A(n_8538),
.B(n_7887),
.Y(n_10183)
);

AOI22xp33_ASAP7_75t_SL g10184 ( 
.A1(n_8802),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_L g10185 ( 
.A(n_9187),
.B(n_7775),
.Y(n_10185)
);

INVx3_ASAP7_75t_L g10186 ( 
.A(n_9070),
.Y(n_10186)
);

OAI21xp33_ASAP7_75t_L g10187 ( 
.A1(n_8439),
.A2(n_8287),
.B(n_8329),
.Y(n_10187)
);

INVx1_ASAP7_75t_L g10188 ( 
.A(n_8201),
.Y(n_10188)
);

INVx3_ASAP7_75t_L g10189 ( 
.A(n_9070),
.Y(n_10189)
);

AND2x2_ASAP7_75t_L g10190 ( 
.A(n_8538),
.B(n_7887),
.Y(n_10190)
);

CKINVDCx20_ASAP7_75t_R g10191 ( 
.A(n_9324),
.Y(n_10191)
);

INVx1_ASAP7_75t_L g10192 ( 
.A(n_8201),
.Y(n_10192)
);

INVx2_ASAP7_75t_L g10193 ( 
.A(n_9458),
.Y(n_10193)
);

NAND2xp5_ASAP7_75t_L g10194 ( 
.A(n_9187),
.B(n_7775),
.Y(n_10194)
);

INVx1_ASAP7_75t_SL g10195 ( 
.A(n_9324),
.Y(n_10195)
);

HB1xp67_ASAP7_75t_L g10196 ( 
.A(n_9312),
.Y(n_10196)
);

HB1xp67_ASAP7_75t_L g10197 ( 
.A(n_9312),
.Y(n_10197)
);

INVx3_ASAP7_75t_L g10198 ( 
.A(n_9070),
.Y(n_10198)
);

INVx1_ASAP7_75t_L g10199 ( 
.A(n_8201),
.Y(n_10199)
);

INVx1_ASAP7_75t_L g10200 ( 
.A(n_8235),
.Y(n_10200)
);

INVx2_ASAP7_75t_L g10201 ( 
.A(n_9475),
.Y(n_10201)
);

OAI21xp5_ASAP7_75t_L g10202 ( 
.A1(n_8327),
.A2(n_7973),
.B(n_7897),
.Y(n_10202)
);

INVx2_ASAP7_75t_L g10203 ( 
.A(n_9475),
.Y(n_10203)
);

AOI22xp5_ASAP7_75t_L g10204 ( 
.A1(n_8416),
.A2(n_7082),
.B1(n_8039),
.B2(n_7203),
.Y(n_10204)
);

INVx3_ASAP7_75t_L g10205 ( 
.A(n_9070),
.Y(n_10205)
);

AO21x1_ASAP7_75t_L g10206 ( 
.A1(n_8864),
.A2(n_7794),
.B(n_7789),
.Y(n_10206)
);

OAI22xp5_ASAP7_75t_L g10207 ( 
.A1(n_8467),
.A2(n_7291),
.B1(n_7482),
.B2(n_7897),
.Y(n_10207)
);

NAND2x1p5_ASAP7_75t_L g10208 ( 
.A(n_8276),
.B(n_7509),
.Y(n_10208)
);

AND2x2_ASAP7_75t_L g10209 ( 
.A(n_8559),
.B(n_7887),
.Y(n_10209)
);

NOR2xp67_ASAP7_75t_L g10210 ( 
.A(n_8454),
.B(n_7919),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_9475),
.Y(n_10211)
);

INVx2_ASAP7_75t_L g10212 ( 
.A(n_9475),
.Y(n_10212)
);

AND2x2_ASAP7_75t_L g10213 ( 
.A(n_8559),
.B(n_7919),
.Y(n_10213)
);

NAND2xp5_ASAP7_75t_L g10214 ( 
.A(n_9213),
.B(n_7789),
.Y(n_10214)
);

BUFx2_ASAP7_75t_L g10215 ( 
.A(n_8218),
.Y(n_10215)
);

BUFx6f_ASAP7_75t_L g10216 ( 
.A(n_8605),
.Y(n_10216)
);

AOI21x1_ASAP7_75t_L g10217 ( 
.A1(n_8188),
.A2(n_8242),
.B(n_8802),
.Y(n_10217)
);

INVx1_ASAP7_75t_L g10218 ( 
.A(n_8235),
.Y(n_10218)
);

AND2x2_ASAP7_75t_L g10219 ( 
.A(n_8559),
.B(n_8633),
.Y(n_10219)
);

INVx1_ASAP7_75t_L g10220 ( 
.A(n_8235),
.Y(n_10220)
);

OA21x2_ASAP7_75t_L g10221 ( 
.A1(n_8249),
.A2(n_8682),
.B(n_8255),
.Y(n_10221)
);

BUFx6f_ASAP7_75t_L g10222 ( 
.A(n_8605),
.Y(n_10222)
);

HB1xp67_ASAP7_75t_L g10223 ( 
.A(n_9312),
.Y(n_10223)
);

INVx2_ASAP7_75t_SL g10224 ( 
.A(n_9440),
.Y(n_10224)
);

HB1xp67_ASAP7_75t_L g10225 ( 
.A(n_9343),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_8248),
.Y(n_10226)
);

AOI22xp33_ASAP7_75t_SL g10227 ( 
.A1(n_8802),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10227)
);

INVx2_ASAP7_75t_L g10228 ( 
.A(n_9475),
.Y(n_10228)
);

BUFx12f_ASAP7_75t_L g10229 ( 
.A(n_8925),
.Y(n_10229)
);

CKINVDCx5p33_ASAP7_75t_R g10230 ( 
.A(n_9182),
.Y(n_10230)
);

AOI22xp33_ASAP7_75t_L g10231 ( 
.A1(n_8183),
.A2(n_7323),
.B1(n_6927),
.B2(n_7123),
.Y(n_10231)
);

CKINVDCx6p67_ASAP7_75t_R g10232 ( 
.A(n_8619),
.Y(n_10232)
);

BUFx3_ASAP7_75t_L g10233 ( 
.A(n_8925),
.Y(n_10233)
);

INVx1_ASAP7_75t_L g10234 ( 
.A(n_8248),
.Y(n_10234)
);

INVx2_ASAP7_75t_L g10235 ( 
.A(n_9475),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_8248),
.Y(n_10236)
);

INVx2_ASAP7_75t_L g10237 ( 
.A(n_8291),
.Y(n_10237)
);

INVx1_ASAP7_75t_L g10238 ( 
.A(n_8253),
.Y(n_10238)
);

INVx1_ASAP7_75t_L g10239 ( 
.A(n_8253),
.Y(n_10239)
);

INVx2_ASAP7_75t_L g10240 ( 
.A(n_8291),
.Y(n_10240)
);

INVx1_ASAP7_75t_L g10241 ( 
.A(n_8253),
.Y(n_10241)
);

CKINVDCx20_ASAP7_75t_R g10242 ( 
.A(n_8171),
.Y(n_10242)
);

INVx1_ASAP7_75t_L g10243 ( 
.A(n_8261),
.Y(n_10243)
);

INVx2_ASAP7_75t_L g10244 ( 
.A(n_8291),
.Y(n_10244)
);

INVx1_ASAP7_75t_L g10245 ( 
.A(n_8261),
.Y(n_10245)
);

OAI22xp5_ASAP7_75t_L g10246 ( 
.A1(n_8467),
.A2(n_8424),
.B1(n_8324),
.B2(n_8869),
.Y(n_10246)
);

INVx2_ASAP7_75t_SL g10247 ( 
.A(n_8649),
.Y(n_10247)
);

OAI22xp33_ASAP7_75t_L g10248 ( 
.A1(n_8827),
.A2(n_7135),
.B1(n_7203),
.B2(n_7409),
.Y(n_10248)
);

INVx1_ASAP7_75t_L g10249 ( 
.A(n_8261),
.Y(n_10249)
);

AOI22xp33_ASAP7_75t_L g10250 ( 
.A1(n_8183),
.A2(n_7323),
.B1(n_6927),
.B2(n_7123),
.Y(n_10250)
);

INVx3_ASAP7_75t_L g10251 ( 
.A(n_9087),
.Y(n_10251)
);

AOI22xp33_ASAP7_75t_SL g10252 ( 
.A1(n_9225),
.A2(n_8324),
.B1(n_8268),
.B2(n_8447),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_8265),
.Y(n_10253)
);

OAI22xp5_ASAP7_75t_L g10254 ( 
.A1(n_8424),
.A2(n_7973),
.B1(n_7982),
.B2(n_7952),
.Y(n_10254)
);

BUFx12f_ASAP7_75t_L g10255 ( 
.A(n_8925),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_8265),
.Y(n_10256)
);

INVx2_ASAP7_75t_L g10257 ( 
.A(n_8291),
.Y(n_10257)
);

CKINVDCx6p67_ASAP7_75t_R g10258 ( 
.A(n_8756),
.Y(n_10258)
);

INVx3_ASAP7_75t_L g10259 ( 
.A(n_9087),
.Y(n_10259)
);

AND2x2_ASAP7_75t_L g10260 ( 
.A(n_8633),
.B(n_7919),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_8265),
.Y(n_10261)
);

INVx1_ASAP7_75t_L g10262 ( 
.A(n_8273),
.Y(n_10262)
);

INVx1_ASAP7_75t_SL g10263 ( 
.A(n_9110),
.Y(n_10263)
);

INVx1_ASAP7_75t_L g10264 ( 
.A(n_8273),
.Y(n_10264)
);

AOI22xp33_ASAP7_75t_L g10265 ( 
.A1(n_9225),
.A2(n_7323),
.B1(n_7118),
.B2(n_7148),
.Y(n_10265)
);

INVx1_ASAP7_75t_L g10266 ( 
.A(n_8273),
.Y(n_10266)
);

INVx3_ASAP7_75t_L g10267 ( 
.A(n_9087),
.Y(n_10267)
);

INVx2_ASAP7_75t_L g10268 ( 
.A(n_8291),
.Y(n_10268)
);

CKINVDCx11_ASAP7_75t_R g10269 ( 
.A(n_8756),
.Y(n_10269)
);

BUFx2_ASAP7_75t_L g10270 ( 
.A(n_8462),
.Y(n_10270)
);

INVx3_ASAP7_75t_L g10271 ( 
.A(n_9087),
.Y(n_10271)
);

OR2x2_ASAP7_75t_L g10272 ( 
.A(n_8174),
.B(n_7194),
.Y(n_10272)
);

AOI22xp5_ASAP7_75t_L g10273 ( 
.A1(n_8473),
.A2(n_8039),
.B1(n_7252),
.B2(n_7042),
.Y(n_10273)
);

BUFx2_ASAP7_75t_R g10274 ( 
.A(n_8171),
.Y(n_10274)
);

AOI22xp33_ASAP7_75t_L g10275 ( 
.A1(n_8932),
.A2(n_7323),
.B1(n_7118),
.B2(n_7148),
.Y(n_10275)
);

INVx1_ASAP7_75t_L g10276 ( 
.A(n_8283),
.Y(n_10276)
);

BUFx2_ASAP7_75t_L g10277 ( 
.A(n_8462),
.Y(n_10277)
);

INVx1_ASAP7_75t_SL g10278 ( 
.A(n_9110),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_8283),
.Y(n_10279)
);

NAND2xp5_ASAP7_75t_L g10280 ( 
.A(n_9213),
.B(n_7789),
.Y(n_10280)
);

AOI22xp33_ASAP7_75t_L g10281 ( 
.A1(n_8932),
.A2(n_7323),
.B1(n_7118),
.B2(n_7148),
.Y(n_10281)
);

INVx1_ASAP7_75t_L g10282 ( 
.A(n_8283),
.Y(n_10282)
);

AOI22xp5_ASAP7_75t_L g10283 ( 
.A1(n_8473),
.A2(n_7252),
.B1(n_7042),
.B2(n_7409),
.Y(n_10283)
);

AOI22xp33_ASAP7_75t_SL g10284 ( 
.A1(n_8268),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10284)
);

AO21x1_ASAP7_75t_L g10285 ( 
.A1(n_8864),
.A2(n_7794),
.B(n_7324),
.Y(n_10285)
);

INVx1_ASAP7_75t_L g10286 ( 
.A(n_8298),
.Y(n_10286)
);

INVx2_ASAP7_75t_L g10287 ( 
.A(n_8291),
.Y(n_10287)
);

OR2x6_ASAP7_75t_L g10288 ( 
.A(n_8454),
.B(n_7323),
.Y(n_10288)
);

INVx1_ASAP7_75t_L g10289 ( 
.A(n_8298),
.Y(n_10289)
);

AND2x2_ASAP7_75t_L g10290 ( 
.A(n_8633),
.B(n_7919),
.Y(n_10290)
);

INVx1_ASAP7_75t_L g10291 ( 
.A(n_8298),
.Y(n_10291)
);

OAI22xp5_ASAP7_75t_L g10292 ( 
.A1(n_8869),
.A2(n_8355),
.B1(n_8287),
.B2(n_8503),
.Y(n_10292)
);

BUFx6f_ASAP7_75t_SL g10293 ( 
.A(n_8605),
.Y(n_10293)
);

AOI22xp33_ASAP7_75t_L g10294 ( 
.A1(n_8932),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10294)
);

HB1xp67_ASAP7_75t_L g10295 ( 
.A(n_9343),
.Y(n_10295)
);

INVx1_ASAP7_75t_SL g10296 ( 
.A(n_8709),
.Y(n_10296)
);

INVx2_ASAP7_75t_L g10297 ( 
.A(n_8354),
.Y(n_10297)
);

OA21x2_ASAP7_75t_L g10298 ( 
.A1(n_8682),
.A2(n_7239),
.B(n_7234),
.Y(n_10298)
);

AOI22xp33_ASAP7_75t_L g10299 ( 
.A1(n_8932),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10299)
);

AOI22xp33_ASAP7_75t_L g10300 ( 
.A1(n_8932),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10300)
);

BUFx8_ASAP7_75t_L g10301 ( 
.A(n_8925),
.Y(n_10301)
);

AOI21x1_ASAP7_75t_L g10302 ( 
.A1(n_8335),
.A2(n_7416),
.B(n_7403),
.Y(n_10302)
);

AND2x4_ASAP7_75t_L g10303 ( 
.A(n_8627),
.B(n_7949),
.Y(n_10303)
);

OA21x2_ASAP7_75t_L g10304 ( 
.A1(n_8682),
.A2(n_7239),
.B(n_7234),
.Y(n_10304)
);

INVx2_ASAP7_75t_L g10305 ( 
.A(n_8354),
.Y(n_10305)
);

INVx3_ASAP7_75t_L g10306 ( 
.A(n_9087),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_8303),
.Y(n_10307)
);

INVx2_ASAP7_75t_L g10308 ( 
.A(n_8354),
.Y(n_10308)
);

BUFx3_ASAP7_75t_L g10309 ( 
.A(n_8649),
.Y(n_10309)
);

AOI22xp33_ASAP7_75t_SL g10310 ( 
.A1(n_8628),
.A2(n_7374),
.B1(n_7412),
.B2(n_7404),
.Y(n_10310)
);

INVx2_ASAP7_75t_L g10311 ( 
.A(n_8354),
.Y(n_10311)
);

BUFx3_ASAP7_75t_L g10312 ( 
.A(n_8649),
.Y(n_10312)
);

INVx4_ASAP7_75t_L g10313 ( 
.A(n_8844),
.Y(n_10313)
);

INVx3_ASAP7_75t_L g10314 ( 
.A(n_9087),
.Y(n_10314)
);

INVx1_ASAP7_75t_L g10315 ( 
.A(n_8303),
.Y(n_10315)
);

INVx2_ASAP7_75t_L g10316 ( 
.A(n_8354),
.Y(n_10316)
);

OAI21x1_ASAP7_75t_SL g10317 ( 
.A1(n_8818),
.A2(n_7032),
.B(n_6935),
.Y(n_10317)
);

CKINVDCx11_ASAP7_75t_R g10318 ( 
.A(n_8756),
.Y(n_10318)
);

INVx1_ASAP7_75t_L g10319 ( 
.A(n_8303),
.Y(n_10319)
);

BUFx3_ASAP7_75t_L g10320 ( 
.A(n_8649),
.Y(n_10320)
);

INVx3_ASAP7_75t_SL g10321 ( 
.A(n_8644),
.Y(n_10321)
);

OAI22xp5_ASAP7_75t_L g10322 ( 
.A1(n_8355),
.A2(n_7982),
.B1(n_7952),
.B2(n_7754),
.Y(n_10322)
);

AND2x4_ASAP7_75t_L g10323 ( 
.A(n_8720),
.B(n_7949),
.Y(n_10323)
);

CKINVDCx11_ASAP7_75t_R g10324 ( 
.A(n_8756),
.Y(n_10324)
);

OAI21x1_ASAP7_75t_SL g10325 ( 
.A1(n_8818),
.A2(n_7065),
.B(n_6935),
.Y(n_10325)
);

INVx1_ASAP7_75t_L g10326 ( 
.A(n_8334),
.Y(n_10326)
);

OAI21x1_ASAP7_75t_SL g10327 ( 
.A1(n_8818),
.A2(n_7080),
.B(n_7065),
.Y(n_10327)
);

CKINVDCx20_ASAP7_75t_R g10328 ( 
.A(n_8269),
.Y(n_10328)
);

AO21x1_ASAP7_75t_L g10329 ( 
.A1(n_9431),
.A2(n_8812),
.B(n_8329),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_8334),
.Y(n_10330)
);

AND2x2_ASAP7_75t_L g10331 ( 
.A(n_8678),
.B(n_7949),
.Y(n_10331)
);

AO21x2_ASAP7_75t_L g10332 ( 
.A1(n_8185),
.A2(n_7997),
.B(n_7981),
.Y(n_10332)
);

INVx3_ASAP7_75t_L g10333 ( 
.A(n_8530),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_8334),
.Y(n_10334)
);

INVx2_ASAP7_75t_L g10335 ( 
.A(n_8354),
.Y(n_10335)
);

INVx2_ASAP7_75t_L g10336 ( 
.A(n_8393),
.Y(n_10336)
);

NAND2xp5_ASAP7_75t_L g10337 ( 
.A(n_8801),
.B(n_8761),
.Y(n_10337)
);

INVx2_ASAP7_75t_SL g10338 ( 
.A(n_8649),
.Y(n_10338)
);

INVx2_ASAP7_75t_L g10339 ( 
.A(n_8393),
.Y(n_10339)
);

HB1xp67_ASAP7_75t_L g10340 ( 
.A(n_9343),
.Y(n_10340)
);

BUFx6f_ASAP7_75t_L g10341 ( 
.A(n_8717),
.Y(n_10341)
);

BUFx2_ASAP7_75t_R g10342 ( 
.A(n_8269),
.Y(n_10342)
);

INVx2_ASAP7_75t_L g10343 ( 
.A(n_8393),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_8393),
.Y(n_10344)
);

AOI21x1_ASAP7_75t_L g10345 ( 
.A1(n_8335),
.A2(n_7418),
.B(n_7416),
.Y(n_10345)
);

NOR2x1_ASAP7_75t_R g10346 ( 
.A(n_8630),
.B(n_7283),
.Y(n_10346)
);

CKINVDCx16_ASAP7_75t_R g10347 ( 
.A(n_8350),
.Y(n_10347)
);

AOI22xp33_ASAP7_75t_L g10348 ( 
.A1(n_8503),
.A2(n_8214),
.B1(n_8356),
.B2(n_8337),
.Y(n_10348)
);

INVx1_ASAP7_75t_L g10349 ( 
.A(n_8339),
.Y(n_10349)
);

INVx6_ASAP7_75t_L g10350 ( 
.A(n_8879),
.Y(n_10350)
);

INVx1_ASAP7_75t_L g10351 ( 
.A(n_8339),
.Y(n_10351)
);

INVx1_ASAP7_75t_L g10352 ( 
.A(n_8339),
.Y(n_10352)
);

BUFx2_ASAP7_75t_L g10353 ( 
.A(n_8462),
.Y(n_10353)
);

HB1xp67_ASAP7_75t_L g10354 ( 
.A(n_9343),
.Y(n_10354)
);

INVx2_ASAP7_75t_L g10355 ( 
.A(n_8393),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_8343),
.Y(n_10356)
);

CKINVDCx12_ASAP7_75t_R g10357 ( 
.A(n_8338),
.Y(n_10357)
);

INVx1_ASAP7_75t_L g10358 ( 
.A(n_8343),
.Y(n_10358)
);

INVx2_ASAP7_75t_L g10359 ( 
.A(n_8426),
.Y(n_10359)
);

INVx1_ASAP7_75t_L g10360 ( 
.A(n_8343),
.Y(n_10360)
);

AOI22xp33_ASAP7_75t_L g10361 ( 
.A1(n_8214),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10361)
);

INVx1_ASAP7_75t_L g10362 ( 
.A(n_8351),
.Y(n_10362)
);

OAI22xp33_ASAP7_75t_L g10363 ( 
.A1(n_8827),
.A2(n_7417),
.B1(n_7409),
.B2(n_7990),
.Y(n_10363)
);

INVx1_ASAP7_75t_L g10364 ( 
.A(n_8351),
.Y(n_10364)
);

INVx4_ASAP7_75t_L g10365 ( 
.A(n_8844),
.Y(n_10365)
);

BUFx2_ASAP7_75t_L g10366 ( 
.A(n_8462),
.Y(n_10366)
);

INVx1_ASAP7_75t_L g10367 ( 
.A(n_8351),
.Y(n_10367)
);

AOI22xp33_ASAP7_75t_L g10368 ( 
.A1(n_8214),
.A2(n_8356),
.B1(n_8337),
.B2(n_8692),
.Y(n_10368)
);

OAI22xp5_ASAP7_75t_L g10369 ( 
.A1(n_8423),
.A2(n_7982),
.B1(n_7952),
.B2(n_7754),
.Y(n_10369)
);

OAI22xp5_ASAP7_75t_L g10370 ( 
.A1(n_8423),
.A2(n_7754),
.B1(n_7043),
.B2(n_7247),
.Y(n_10370)
);

BUFx8_ASAP7_75t_L g10371 ( 
.A(n_8717),
.Y(n_10371)
);

CKINVDCx20_ASAP7_75t_R g10372 ( 
.A(n_8361),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_8373),
.Y(n_10373)
);

OAI22xp5_ASAP7_75t_L g10374 ( 
.A1(n_8422),
.A2(n_7043),
.B1(n_7247),
.B2(n_7990),
.Y(n_10374)
);

AOI22xp33_ASAP7_75t_L g10375 ( 
.A1(n_8214),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10375)
);

BUFx2_ASAP7_75t_R g10376 ( 
.A(n_8361),
.Y(n_10376)
);

BUFx6f_ASAP7_75t_L g10377 ( 
.A(n_8717),
.Y(n_10377)
);

AO21x2_ASAP7_75t_L g10378 ( 
.A1(n_8185),
.A2(n_7997),
.B(n_7981),
.Y(n_10378)
);

INVx6_ASAP7_75t_L g10379 ( 
.A(n_9174),
.Y(n_10379)
);

AOI22xp33_ASAP7_75t_SL g10380 ( 
.A1(n_8628),
.A2(n_7404),
.B1(n_7412),
.B2(n_7374),
.Y(n_10380)
);

INVx1_ASAP7_75t_L g10381 ( 
.A(n_8373),
.Y(n_10381)
);

INVx2_ASAP7_75t_L g10382 ( 
.A(n_8426),
.Y(n_10382)
);

INVx1_ASAP7_75t_L g10383 ( 
.A(n_8373),
.Y(n_10383)
);

HB1xp67_ASAP7_75t_L g10384 ( 
.A(n_9343),
.Y(n_10384)
);

AOI22xp33_ASAP7_75t_SL g10385 ( 
.A1(n_8628),
.A2(n_8836),
.B1(n_8848),
.B2(n_8814),
.Y(n_10385)
);

AOI22xp33_ASAP7_75t_L g10386 ( 
.A1(n_8214),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10386)
);

AND2x4_ASAP7_75t_L g10387 ( 
.A(n_8627),
.B(n_7949),
.Y(n_10387)
);

BUFx2_ASAP7_75t_R g10388 ( 
.A(n_8412),
.Y(n_10388)
);

BUFx6f_ASAP7_75t_L g10389 ( 
.A(n_8717),
.Y(n_10389)
);

INVxp67_ASAP7_75t_L g10390 ( 
.A(n_8349),
.Y(n_10390)
);

AND2x2_ASAP7_75t_L g10391 ( 
.A(n_8678),
.B(n_7955),
.Y(n_10391)
);

INVx2_ASAP7_75t_L g10392 ( 
.A(n_8426),
.Y(n_10392)
);

OR2x2_ASAP7_75t_L g10393 ( 
.A(n_8230),
.B(n_7194),
.Y(n_10393)
);

OA21x2_ASAP7_75t_L g10394 ( 
.A1(n_8254),
.A2(n_7239),
.B(n_6993),
.Y(n_10394)
);

BUFx6f_ASAP7_75t_L g10395 ( 
.A(n_8644),
.Y(n_10395)
);

AND2x4_ASAP7_75t_L g10396 ( 
.A(n_8627),
.B(n_7955),
.Y(n_10396)
);

INVx1_ASAP7_75t_L g10397 ( 
.A(n_8375),
.Y(n_10397)
);

INVx4_ASAP7_75t_L g10398 ( 
.A(n_8844),
.Y(n_10398)
);

INVx5_ASAP7_75t_L g10399 ( 
.A(n_9358),
.Y(n_10399)
);

CKINVDCx20_ASAP7_75t_R g10400 ( 
.A(n_8412),
.Y(n_10400)
);

INVx1_ASAP7_75t_L g10401 ( 
.A(n_8375),
.Y(n_10401)
);

OR2x2_ASAP7_75t_L g10402 ( 
.A(n_8230),
.B(n_7208),
.Y(n_10402)
);

INVx2_ASAP7_75t_L g10403 ( 
.A(n_8426),
.Y(n_10403)
);

NAND2xp5_ASAP7_75t_L g10404 ( 
.A(n_8801),
.B(n_7794),
.Y(n_10404)
);

AOI21x1_ASAP7_75t_L g10405 ( 
.A1(n_8584),
.A2(n_7418),
.B(n_7416),
.Y(n_10405)
);

AOI22xp33_ASAP7_75t_L g10406 ( 
.A1(n_8692),
.A2(n_7118),
.B1(n_7148),
.B2(n_7123),
.Y(n_10406)
);

OAI21xp5_ASAP7_75t_L g10407 ( 
.A1(n_8431),
.A2(n_8392),
.B(n_8980),
.Y(n_10407)
);

INVx1_ASAP7_75t_L g10408 ( 
.A(n_8375),
.Y(n_10408)
);

INVx1_ASAP7_75t_SL g10409 ( 
.A(n_8709),
.Y(n_10409)
);

AO22x1_ASAP7_75t_L g10410 ( 
.A1(n_8392),
.A2(n_7445),
.B1(n_7443),
.B2(n_7080),
.Y(n_10410)
);

INVx1_ASAP7_75t_L g10411 ( 
.A(n_8379),
.Y(n_10411)
);

INVx1_ASAP7_75t_L g10412 ( 
.A(n_8379),
.Y(n_10412)
);

INVx2_ASAP7_75t_L g10413 ( 
.A(n_8426),
.Y(n_10413)
);

OR2x2_ASAP7_75t_L g10414 ( 
.A(n_8294),
.B(n_7208),
.Y(n_10414)
);

INVx2_ASAP7_75t_L g10415 ( 
.A(n_8426),
.Y(n_10415)
);

INVx6_ASAP7_75t_L g10416 ( 
.A(n_9174),
.Y(n_10416)
);

INVx2_ASAP7_75t_L g10417 ( 
.A(n_8445),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_8379),
.Y(n_10418)
);

INVx2_ASAP7_75t_L g10419 ( 
.A(n_8445),
.Y(n_10419)
);

INVx2_ASAP7_75t_SL g10420 ( 
.A(n_8844),
.Y(n_10420)
);

INVx2_ASAP7_75t_L g10421 ( 
.A(n_8445),
.Y(n_10421)
);

INVx3_ASAP7_75t_L g10422 ( 
.A(n_8530),
.Y(n_10422)
);

AOI22xp33_ASAP7_75t_SL g10423 ( 
.A1(n_8814),
.A2(n_7404),
.B1(n_7412),
.B2(n_7374),
.Y(n_10423)
);

AND2x4_ASAP7_75t_L g10424 ( 
.A(n_8627),
.B(n_8720),
.Y(n_10424)
);

INVx3_ASAP7_75t_L g10425 ( 
.A(n_8530),
.Y(n_10425)
);

INVx1_ASAP7_75t_SL g10426 ( 
.A(n_8881),
.Y(n_10426)
);

OAI22xp33_ASAP7_75t_L g10427 ( 
.A1(n_8622),
.A2(n_7417),
.B1(n_8009),
.B2(n_7990),
.Y(n_10427)
);

INVx2_ASAP7_75t_L g10428 ( 
.A(n_8445),
.Y(n_10428)
);

NAND2xp5_ASAP7_75t_L g10429 ( 
.A(n_8761),
.B(n_8665),
.Y(n_10429)
);

AOI22xp5_ASAP7_75t_L g10430 ( 
.A1(n_8395),
.A2(n_7042),
.B1(n_7417),
.B2(n_7681),
.Y(n_10430)
);

INVx1_ASAP7_75t_L g10431 ( 
.A(n_8384),
.Y(n_10431)
);

INVx3_ASAP7_75t_L g10432 ( 
.A(n_8530),
.Y(n_10432)
);

INVx2_ASAP7_75t_L g10433 ( 
.A(n_8445),
.Y(n_10433)
);

BUFx12f_ASAP7_75t_L g10434 ( 
.A(n_9174),
.Y(n_10434)
);

HB1xp67_ASAP7_75t_L g10435 ( 
.A(n_9343),
.Y(n_10435)
);

INVx1_ASAP7_75t_L g10436 ( 
.A(n_8384),
.Y(n_10436)
);

INVx1_ASAP7_75t_L g10437 ( 
.A(n_8384),
.Y(n_10437)
);

CKINVDCx11_ASAP7_75t_R g10438 ( 
.A(n_9457),
.Y(n_10438)
);

BUFx2_ASAP7_75t_L g10439 ( 
.A(n_8462),
.Y(n_10439)
);

OAI22xp5_ASAP7_75t_L g10440 ( 
.A1(n_8422),
.A2(n_7247),
.B1(n_8009),
.B2(n_7900),
.Y(n_10440)
);

INVx3_ASAP7_75t_L g10441 ( 
.A(n_8530),
.Y(n_10441)
);

INVx5_ASAP7_75t_L g10442 ( 
.A(n_9358),
.Y(n_10442)
);

INVx1_ASAP7_75t_L g10443 ( 
.A(n_8389),
.Y(n_10443)
);

INVx1_ASAP7_75t_L g10444 ( 
.A(n_8389),
.Y(n_10444)
);

AOI22xp33_ASAP7_75t_L g10445 ( 
.A1(n_9431),
.A2(n_7123),
.B1(n_7211),
.B2(n_7196),
.Y(n_10445)
);

INVx2_ASAP7_75t_L g10446 ( 
.A(n_8445),
.Y(n_10446)
);

NAND2xp5_ASAP7_75t_L g10447 ( 
.A(n_8665),
.B(n_7320),
.Y(n_10447)
);

BUFx8_ASAP7_75t_L g10448 ( 
.A(n_8674),
.Y(n_10448)
);

OR2x6_ASAP7_75t_L g10449 ( 
.A(n_8521),
.B(n_8033),
.Y(n_10449)
);

INVx2_ASAP7_75t_L g10450 ( 
.A(n_8471),
.Y(n_10450)
);

INVx1_ASAP7_75t_L g10451 ( 
.A(n_8389),
.Y(n_10451)
);

INVx1_ASAP7_75t_L g10452 ( 
.A(n_8398),
.Y(n_10452)
);

NOR2x1_ASAP7_75t_R g10453 ( 
.A(n_8630),
.B(n_7283),
.Y(n_10453)
);

AND2x2_ASAP7_75t_L g10454 ( 
.A(n_8678),
.B(n_7955),
.Y(n_10454)
);

BUFx2_ASAP7_75t_L g10455 ( 
.A(n_8462),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_8398),
.Y(n_10456)
);

BUFx6f_ASAP7_75t_L g10457 ( 
.A(n_8644),
.Y(n_10457)
);

BUFx6f_ASAP7_75t_L g10458 ( 
.A(n_8471),
.Y(n_10458)
);

OAI21x1_ASAP7_75t_L g10459 ( 
.A1(n_8464),
.A2(n_7013),
.B(n_6967),
.Y(n_10459)
);

AOI22xp33_ASAP7_75t_SL g10460 ( 
.A1(n_8814),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10460)
);

AOI22xp33_ASAP7_75t_SL g10461 ( 
.A1(n_8814),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10461)
);

INVx2_ASAP7_75t_L g10462 ( 
.A(n_8471),
.Y(n_10462)
);

INVx1_ASAP7_75t_L g10463 ( 
.A(n_8398),
.Y(n_10463)
);

OR2x6_ASAP7_75t_L g10464 ( 
.A(n_8521),
.B(n_8202),
.Y(n_10464)
);

INVx4_ASAP7_75t_L g10465 ( 
.A(n_8844),
.Y(n_10465)
);

INVx1_ASAP7_75t_L g10466 ( 
.A(n_8436),
.Y(n_10466)
);

OAI22xp33_ASAP7_75t_L g10467 ( 
.A1(n_8622),
.A2(n_8009),
.B1(n_7270),
.B2(n_6933),
.Y(n_10467)
);

AOI22xp33_ASAP7_75t_SL g10468 ( 
.A1(n_8836),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10468)
);

AND2x2_ASAP7_75t_L g10469 ( 
.A(n_8891),
.B(n_7955),
.Y(n_10469)
);

HB1xp67_ASAP7_75t_L g10470 ( 
.A(n_9343),
.Y(n_10470)
);

INVx3_ASAP7_75t_L g10471 ( 
.A(n_8530),
.Y(n_10471)
);

INVx2_ASAP7_75t_L g10472 ( 
.A(n_8471),
.Y(n_10472)
);

BUFx2_ASAP7_75t_L g10473 ( 
.A(n_8462),
.Y(n_10473)
);

OAI21x1_ASAP7_75t_L g10474 ( 
.A1(n_8599),
.A2(n_7013),
.B(n_6967),
.Y(n_10474)
);

NAND2x1p5_ASAP7_75t_L g10475 ( 
.A(n_8276),
.B(n_7509),
.Y(n_10475)
);

BUFx3_ASAP7_75t_L g10476 ( 
.A(n_9174),
.Y(n_10476)
);

OAI21xp5_ASAP7_75t_L g10477 ( 
.A1(n_8431),
.A2(n_7993),
.B(n_7951),
.Y(n_10477)
);

INVx1_ASAP7_75t_L g10478 ( 
.A(n_8436),
.Y(n_10478)
);

AOI22xp33_ASAP7_75t_L g10479 ( 
.A1(n_8563),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10479)
);

INVx1_ASAP7_75t_L g10480 ( 
.A(n_8436),
.Y(n_10480)
);

NAND2x1p5_ASAP7_75t_L g10481 ( 
.A(n_8276),
.B(n_7509),
.Y(n_10481)
);

INVx4_ASAP7_75t_L g10482 ( 
.A(n_8844),
.Y(n_10482)
);

INVx1_ASAP7_75t_SL g10483 ( 
.A(n_8881),
.Y(n_10483)
);

INVx2_ASAP7_75t_L g10484 ( 
.A(n_8471),
.Y(n_10484)
);

AOI22xp5_ASAP7_75t_L g10485 ( 
.A1(n_8395),
.A2(n_8511),
.B1(n_8996),
.B2(n_8563),
.Y(n_10485)
);

BUFx12f_ASAP7_75t_L g10486 ( 
.A(n_9174),
.Y(n_10486)
);

BUFx2_ASAP7_75t_SL g10487 ( 
.A(n_8240),
.Y(n_10487)
);

OAI22xp33_ASAP7_75t_L g10488 ( 
.A1(n_8781),
.A2(n_7270),
.B1(n_6933),
.B2(n_6968),
.Y(n_10488)
);

AO21x2_ASAP7_75t_L g10489 ( 
.A1(n_8185),
.A2(n_6934),
.B(n_6932),
.Y(n_10489)
);

INVx1_ASAP7_75t_L g10490 ( 
.A(n_8442),
.Y(n_10490)
);

AOI22xp33_ASAP7_75t_SL g10491 ( 
.A1(n_8836),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10491)
);

AND2x2_ASAP7_75t_L g10492 ( 
.A(n_8891),
.B(n_7984),
.Y(n_10492)
);

CKINVDCx20_ASAP7_75t_R g10493 ( 
.A(n_9182),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_8442),
.Y(n_10494)
);

OAI21x1_ASAP7_75t_L g10495 ( 
.A1(n_8789),
.A2(n_8839),
.B(n_8807),
.Y(n_10495)
);

INVx1_ASAP7_75t_L g10496 ( 
.A(n_8442),
.Y(n_10496)
);

OAI22xp5_ASAP7_75t_L g10497 ( 
.A1(n_8340),
.A2(n_7875),
.B1(n_7942),
.B2(n_7900),
.Y(n_10497)
);

CKINVDCx11_ASAP7_75t_R g10498 ( 
.A(n_9457),
.Y(n_10498)
);

INVx1_ASAP7_75t_L g10499 ( 
.A(n_8446),
.Y(n_10499)
);

CKINVDCx11_ASAP7_75t_R g10500 ( 
.A(n_9457),
.Y(n_10500)
);

BUFx2_ASAP7_75t_SL g10501 ( 
.A(n_8240),
.Y(n_10501)
);

OAI21x1_ASAP7_75t_L g10502 ( 
.A1(n_8789),
.A2(n_7013),
.B(n_6967),
.Y(n_10502)
);

OAI22xp5_ASAP7_75t_L g10503 ( 
.A1(n_8340),
.A2(n_7875),
.B1(n_7942),
.B2(n_7951),
.Y(n_10503)
);

BUFx4f_ASAP7_75t_L g10504 ( 
.A(n_8968),
.Y(n_10504)
);

HB1xp67_ASAP7_75t_L g10505 ( 
.A(n_9343),
.Y(n_10505)
);

INVx4_ASAP7_75t_L g10506 ( 
.A(n_8844),
.Y(n_10506)
);

AND2x2_ASAP7_75t_L g10507 ( 
.A(n_8891),
.B(n_7984),
.Y(n_10507)
);

INVx1_ASAP7_75t_L g10508 ( 
.A(n_8446),
.Y(n_10508)
);

AO21x1_ASAP7_75t_L g10509 ( 
.A1(n_8812),
.A2(n_7324),
.B(n_7320),
.Y(n_10509)
);

CKINVDCx11_ASAP7_75t_R g10510 ( 
.A(n_9457),
.Y(n_10510)
);

AND2x2_ASAP7_75t_L g10511 ( 
.A(n_9177),
.B(n_7984),
.Y(n_10511)
);

OA21x2_ASAP7_75t_L g10512 ( 
.A1(n_8254),
.A2(n_6993),
.B(n_6988),
.Y(n_10512)
);

HB1xp67_ASAP7_75t_L g10513 ( 
.A(n_9474),
.Y(n_10513)
);

BUFx2_ASAP7_75t_R g10514 ( 
.A(n_8484),
.Y(n_10514)
);

HB1xp67_ASAP7_75t_L g10515 ( 
.A(n_9474),
.Y(n_10515)
);

INVx3_ASAP7_75t_L g10516 ( 
.A(n_8537),
.Y(n_10516)
);

BUFx6f_ASAP7_75t_L g10517 ( 
.A(n_8471),
.Y(n_10517)
);

AND2x2_ASAP7_75t_SL g10518 ( 
.A(n_8276),
.B(n_7848),
.Y(n_10518)
);

INVx2_ASAP7_75t_L g10519 ( 
.A(n_8140),
.Y(n_10519)
);

INVx3_ASAP7_75t_L g10520 ( 
.A(n_8537),
.Y(n_10520)
);

INVx2_ASAP7_75t_L g10521 ( 
.A(n_8140),
.Y(n_10521)
);

CKINVDCx11_ASAP7_75t_R g10522 ( 
.A(n_8308),
.Y(n_10522)
);

CKINVDCx11_ASAP7_75t_R g10523 ( 
.A(n_8308),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_8446),
.Y(n_10524)
);

BUFx3_ASAP7_75t_L g10525 ( 
.A(n_9174),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_8465),
.Y(n_10526)
);

AND2x2_ASAP7_75t_L g10527 ( 
.A(n_9177),
.B(n_9565),
.Y(n_10527)
);

INVx1_ASAP7_75t_L g10528 ( 
.A(n_8465),
.Y(n_10528)
);

BUFx2_ASAP7_75t_L g10529 ( 
.A(n_8462),
.Y(n_10529)
);

AOI22xp33_ASAP7_75t_L g10530 ( 
.A1(n_8451),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10530)
);

INVx2_ASAP7_75t_SL g10531 ( 
.A(n_9040),
.Y(n_10531)
);

AOI21xp33_ASAP7_75t_L g10532 ( 
.A1(n_8647),
.A2(n_7860),
.B(n_7812),
.Y(n_10532)
);

OA21x2_ASAP7_75t_L g10533 ( 
.A1(n_8254),
.A2(n_8255),
.B(n_8706),
.Y(n_10533)
);

INVx1_ASAP7_75t_L g10534 ( 
.A(n_8465),
.Y(n_10534)
);

INVx2_ASAP7_75t_L g10535 ( 
.A(n_8140),
.Y(n_10535)
);

INVx2_ASAP7_75t_L g10536 ( 
.A(n_8140),
.Y(n_10536)
);

INVx2_ASAP7_75t_L g10537 ( 
.A(n_8140),
.Y(n_10537)
);

BUFx6f_ASAP7_75t_L g10538 ( 
.A(n_8211),
.Y(n_10538)
);

BUFx6f_ASAP7_75t_L g10539 ( 
.A(n_8211),
.Y(n_10539)
);

AOI22xp33_ASAP7_75t_SL g10540 ( 
.A1(n_8836),
.A2(n_8866),
.B1(n_8848),
.B2(n_8276),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_8477),
.Y(n_10541)
);

BUFx6f_ASAP7_75t_L g10542 ( 
.A(n_8211),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_8477),
.Y(n_10543)
);

OR2x6_ASAP7_75t_L g10544 ( 
.A(n_8202),
.B(n_8033),
.Y(n_10544)
);

OAI21x1_ASAP7_75t_L g10545 ( 
.A1(n_8599),
.A2(n_7013),
.B(n_6967),
.Y(n_10545)
);

CKINVDCx11_ASAP7_75t_R g10546 ( 
.A(n_8407),
.Y(n_10546)
);

AOI22xp33_ASAP7_75t_L g10547 ( 
.A1(n_8451),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10547)
);

INVx1_ASAP7_75t_SL g10548 ( 
.A(n_8920),
.Y(n_10548)
);

OAI22xp33_ASAP7_75t_L g10549 ( 
.A1(n_8781),
.A2(n_7270),
.B1(n_6933),
.B2(n_6968),
.Y(n_10549)
);

INVx1_ASAP7_75t_L g10550 ( 
.A(n_8477),
.Y(n_10550)
);

BUFx3_ASAP7_75t_L g10551 ( 
.A(n_9536),
.Y(n_10551)
);

INVx1_ASAP7_75t_L g10552 ( 
.A(n_8483),
.Y(n_10552)
);

INVx1_ASAP7_75t_SL g10553 ( 
.A(n_8920),
.Y(n_10553)
);

NOR2xp33_ASAP7_75t_L g10554 ( 
.A(n_8722),
.B(n_7370),
.Y(n_10554)
);

NOR2xp33_ASAP7_75t_L g10555 ( 
.A(n_8722),
.B(n_7283),
.Y(n_10555)
);

NAND2x1p5_ASAP7_75t_L g10556 ( 
.A(n_8276),
.B(n_7821),
.Y(n_10556)
);

BUFx2_ASAP7_75t_L g10557 ( 
.A(n_8577),
.Y(n_10557)
);

INVx1_ASAP7_75t_L g10558 ( 
.A(n_8483),
.Y(n_10558)
);

OA21x2_ASAP7_75t_L g10559 ( 
.A1(n_8255),
.A2(n_6993),
.B(n_6988),
.Y(n_10559)
);

INVx1_ASAP7_75t_L g10560 ( 
.A(n_8483),
.Y(n_10560)
);

BUFx4_ASAP7_75t_SL g10561 ( 
.A(n_9043),
.Y(n_10561)
);

INVx2_ASAP7_75t_L g10562 ( 
.A(n_8140),
.Y(n_10562)
);

HB1xp67_ASAP7_75t_L g10563 ( 
.A(n_9474),
.Y(n_10563)
);

INVx2_ASAP7_75t_SL g10564 ( 
.A(n_9040),
.Y(n_10564)
);

INVx1_ASAP7_75t_L g10565 ( 
.A(n_8487),
.Y(n_10565)
);

CKINVDCx11_ASAP7_75t_R g10566 ( 
.A(n_8407),
.Y(n_10566)
);

INVxp67_ASAP7_75t_L g10567 ( 
.A(n_8349),
.Y(n_10567)
);

INVx8_ASAP7_75t_L g10568 ( 
.A(n_9040),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_8487),
.Y(n_10569)
);

CKINVDCx11_ASAP7_75t_R g10570 ( 
.A(n_8664),
.Y(n_10570)
);

INVx1_ASAP7_75t_L g10571 ( 
.A(n_8487),
.Y(n_10571)
);

BUFx3_ASAP7_75t_L g10572 ( 
.A(n_9536),
.Y(n_10572)
);

INVx2_ASAP7_75t_L g10573 ( 
.A(n_8140),
.Y(n_10573)
);

AOI22xp33_ASAP7_75t_L g10574 ( 
.A1(n_8506),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_8489),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_8489),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_8489),
.Y(n_10577)
);

NAND2x1p5_ASAP7_75t_L g10578 ( 
.A(n_8480),
.B(n_7821),
.Y(n_10578)
);

INVx2_ASAP7_75t_L g10579 ( 
.A(n_8140),
.Y(n_10579)
);

AOI21x1_ASAP7_75t_L g10580 ( 
.A1(n_8584),
.A2(n_7432),
.B(n_7418),
.Y(n_10580)
);

INVx2_ASAP7_75t_L g10581 ( 
.A(n_8187),
.Y(n_10581)
);

NAND2x1p5_ASAP7_75t_L g10582 ( 
.A(n_8480),
.B(n_7821),
.Y(n_10582)
);

AND2x4_ASAP7_75t_L g10583 ( 
.A(n_8627),
.B(n_7984),
.Y(n_10583)
);

BUFx6f_ASAP7_75t_L g10584 ( 
.A(n_8211),
.Y(n_10584)
);

INVx2_ASAP7_75t_L g10585 ( 
.A(n_8187),
.Y(n_10585)
);

INVx2_ASAP7_75t_L g10586 ( 
.A(n_8187),
.Y(n_10586)
);

INVx2_ASAP7_75t_L g10587 ( 
.A(n_8187),
.Y(n_10587)
);

OAI21x1_ASAP7_75t_L g10588 ( 
.A1(n_8807),
.A2(n_7013),
.B(n_6967),
.Y(n_10588)
);

INVx1_ASAP7_75t_L g10589 ( 
.A(n_8500),
.Y(n_10589)
);

AND2x2_ASAP7_75t_L g10590 ( 
.A(n_9177),
.B(n_9565),
.Y(n_10590)
);

AND2x4_ASAP7_75t_L g10591 ( 
.A(n_8627),
.B(n_8018),
.Y(n_10591)
);

INVx1_ASAP7_75t_L g10592 ( 
.A(n_8500),
.Y(n_10592)
);

BUFx3_ASAP7_75t_L g10593 ( 
.A(n_9536),
.Y(n_10593)
);

OAI21x1_ASAP7_75t_L g10594 ( 
.A1(n_8807),
.A2(n_7062),
.B(n_7013),
.Y(n_10594)
);

INVx2_ASAP7_75t_L g10595 ( 
.A(n_8187),
.Y(n_10595)
);

INVx2_ASAP7_75t_L g10596 ( 
.A(n_8187),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_8500),
.Y(n_10597)
);

INVx1_ASAP7_75t_L g10598 ( 
.A(n_8533),
.Y(n_10598)
);

AOI22xp33_ASAP7_75t_L g10599 ( 
.A1(n_8506),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10599)
);

INVx1_ASAP7_75t_L g10600 ( 
.A(n_8533),
.Y(n_10600)
);

INVx1_ASAP7_75t_L g10601 ( 
.A(n_8533),
.Y(n_10601)
);

BUFx12f_ASAP7_75t_L g10602 ( 
.A(n_9536),
.Y(n_10602)
);

AOI22xp33_ASAP7_75t_L g10603 ( 
.A1(n_8917),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10603)
);

AOI22xp33_ASAP7_75t_L g10604 ( 
.A1(n_8917),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10604)
);

INVx3_ASAP7_75t_L g10605 ( 
.A(n_8537),
.Y(n_10605)
);

BUFx3_ASAP7_75t_L g10606 ( 
.A(n_9536),
.Y(n_10606)
);

OR2x2_ASAP7_75t_L g10607 ( 
.A(n_8294),
.B(n_7208),
.Y(n_10607)
);

AOI22xp33_ASAP7_75t_L g10608 ( 
.A1(n_8917),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10608)
);

INVx3_ASAP7_75t_L g10609 ( 
.A(n_8537),
.Y(n_10609)
);

AND2x4_ASAP7_75t_L g10610 ( 
.A(n_8627),
.B(n_8018),
.Y(n_10610)
);

BUFx4f_ASAP7_75t_L g10611 ( 
.A(n_8968),
.Y(n_10611)
);

HB1xp67_ASAP7_75t_L g10612 ( 
.A(n_9474),
.Y(n_10612)
);

BUFx12f_ASAP7_75t_L g10613 ( 
.A(n_9536),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_8540),
.Y(n_10614)
);

OR2x6_ASAP7_75t_L g10615 ( 
.A(n_8202),
.B(n_8033),
.Y(n_10615)
);

INVx3_ASAP7_75t_L g10616 ( 
.A(n_8537),
.Y(n_10616)
);

AOI22xp33_ASAP7_75t_SL g10617 ( 
.A1(n_8848),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10617)
);

CKINVDCx5p33_ASAP7_75t_R g10618 ( 
.A(n_9242),
.Y(n_10618)
);

INVx2_ASAP7_75t_SL g10619 ( 
.A(n_9040),
.Y(n_10619)
);

AO21x1_ASAP7_75t_L g10620 ( 
.A1(n_8731),
.A2(n_7329),
.B(n_7325),
.Y(n_10620)
);

AND2x2_ASAP7_75t_L g10621 ( 
.A(n_9565),
.B(n_8018),
.Y(n_10621)
);

NAND2x1p5_ASAP7_75t_L g10622 ( 
.A(n_8480),
.B(n_7821),
.Y(n_10622)
);

AOI22xp33_ASAP7_75t_L g10623 ( 
.A1(n_8996),
.A2(n_7196),
.B1(n_7225),
.B2(n_7211),
.Y(n_10623)
);

INVx2_ASAP7_75t_SL g10624 ( 
.A(n_9040),
.Y(n_10624)
);

INVx3_ASAP7_75t_L g10625 ( 
.A(n_8537),
.Y(n_10625)
);

HB1xp67_ASAP7_75t_L g10626 ( 
.A(n_9474),
.Y(n_10626)
);

INVx3_ASAP7_75t_L g10627 ( 
.A(n_8561),
.Y(n_10627)
);

INVxp67_ASAP7_75t_L g10628 ( 
.A(n_8485),
.Y(n_10628)
);

AO21x1_ASAP7_75t_L g10629 ( 
.A1(n_8731),
.A2(n_7329),
.B(n_7325),
.Y(n_10629)
);

CKINVDCx5p33_ASAP7_75t_R g10630 ( 
.A(n_9242),
.Y(n_10630)
);

AOI22xp33_ASAP7_75t_L g10631 ( 
.A1(n_8413),
.A2(n_7225),
.B1(n_7245),
.B2(n_7230),
.Y(n_10631)
);

AOI21x1_ASAP7_75t_L g10632 ( 
.A1(n_8145),
.A2(n_7477),
.B(n_7432),
.Y(n_10632)
);

NAND2x1p5_ASAP7_75t_L g10633 ( 
.A(n_9508),
.B(n_7834),
.Y(n_10633)
);

OAI21x1_ASAP7_75t_L g10634 ( 
.A1(n_8599),
.A2(n_7068),
.B(n_7062),
.Y(n_10634)
);

INVx1_ASAP7_75t_L g10635 ( 
.A(n_8540),
.Y(n_10635)
);

INVx3_ASAP7_75t_L g10636 ( 
.A(n_8561),
.Y(n_10636)
);

OAI21x1_ASAP7_75t_L g10637 ( 
.A1(n_8849),
.A2(n_7068),
.B(n_7062),
.Y(n_10637)
);

CKINVDCx5p33_ASAP7_75t_R g10638 ( 
.A(n_9262),
.Y(n_10638)
);

AO21x1_ASAP7_75t_SL g10639 ( 
.A1(n_8620),
.A2(n_7329),
.B(n_7325),
.Y(n_10639)
);

OAI22xp33_ASAP7_75t_L g10640 ( 
.A1(n_8643),
.A2(n_6968),
.B1(n_8049),
.B2(n_8023),
.Y(n_10640)
);

BUFx2_ASAP7_75t_R g10641 ( 
.A(n_8484),
.Y(n_10641)
);

BUFx2_ASAP7_75t_L g10642 ( 
.A(n_8577),
.Y(n_10642)
);

CKINVDCx5p33_ASAP7_75t_R g10643 ( 
.A(n_9262),
.Y(n_10643)
);

INVx1_ASAP7_75t_L g10644 ( 
.A(n_8540),
.Y(n_10644)
);

BUFx4f_ASAP7_75t_SL g10645 ( 
.A(n_8664),
.Y(n_10645)
);

INVx2_ASAP7_75t_L g10646 ( 
.A(n_8187),
.Y(n_10646)
);

INVx2_ASAP7_75t_L g10647 ( 
.A(n_8187),
.Y(n_10647)
);

INVx1_ASAP7_75t_L g10648 ( 
.A(n_8574),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_8574),
.Y(n_10649)
);

AOI22xp5_ASAP7_75t_SL g10650 ( 
.A1(n_8529),
.A2(n_7065),
.B1(n_7080),
.B2(n_7445),
.Y(n_10650)
);

AOI22xp33_ASAP7_75t_L g10651 ( 
.A1(n_8413),
.A2(n_8370),
.B1(n_8617),
.B2(n_8486),
.Y(n_10651)
);

INVx2_ASAP7_75t_L g10652 ( 
.A(n_9523),
.Y(n_10652)
);

AOI22xp33_ASAP7_75t_SL g10653 ( 
.A1(n_8848),
.A2(n_7483),
.B1(n_7860),
.B2(n_7812),
.Y(n_10653)
);

HB1xp67_ASAP7_75t_L g10654 ( 
.A(n_9474),
.Y(n_10654)
);

INVx2_ASAP7_75t_L g10655 ( 
.A(n_9523),
.Y(n_10655)
);

INVx1_ASAP7_75t_L g10656 ( 
.A(n_8574),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_8590),
.Y(n_10657)
);

INVx1_ASAP7_75t_SL g10658 ( 
.A(n_9010),
.Y(n_10658)
);

BUFx6f_ASAP7_75t_L g10659 ( 
.A(n_8211),
.Y(n_10659)
);

INVx1_ASAP7_75t_L g10660 ( 
.A(n_8590),
.Y(n_10660)
);

INVx2_ASAP7_75t_L g10661 ( 
.A(n_9523),
.Y(n_10661)
);

AND2x2_ASAP7_75t_L g10662 ( 
.A(n_9567),
.B(n_8018),
.Y(n_10662)
);

BUFx2_ASAP7_75t_L g10663 ( 
.A(n_8577),
.Y(n_10663)
);

OA21x2_ASAP7_75t_L g10664 ( 
.A1(n_8706),
.A2(n_6993),
.B(n_6988),
.Y(n_10664)
);

CKINVDCx16_ASAP7_75t_R g10665 ( 
.A(n_8350),
.Y(n_10665)
);

BUFx6f_ASAP7_75t_L g10666 ( 
.A(n_8211),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_8590),
.Y(n_10667)
);

INVx2_ASAP7_75t_L g10668 ( 
.A(n_9259),
.Y(n_10668)
);

CKINVDCx11_ASAP7_75t_R g10669 ( 
.A(n_8702),
.Y(n_10669)
);

HB1xp67_ASAP7_75t_L g10670 ( 
.A(n_9474),
.Y(n_10670)
);

BUFx10_ASAP7_75t_L g10671 ( 
.A(n_8504),
.Y(n_10671)
);

INVx2_ASAP7_75t_SL g10672 ( 
.A(n_9040),
.Y(n_10672)
);

INVx1_ASAP7_75t_L g10673 ( 
.A(n_8600),
.Y(n_10673)
);

AND2x2_ASAP7_75t_L g10674 ( 
.A(n_9567),
.B(n_8037),
.Y(n_10674)
);

CKINVDCx5p33_ASAP7_75t_R g10675 ( 
.A(n_9370),
.Y(n_10675)
);

INVx1_ASAP7_75t_L g10676 ( 
.A(n_8600),
.Y(n_10676)
);

INVx6_ASAP7_75t_L g10677 ( 
.A(n_8257),
.Y(n_10677)
);

OAI21x1_ASAP7_75t_L g10678 ( 
.A1(n_8839),
.A2(n_7068),
.B(n_7062),
.Y(n_10678)
);

AOI22xp5_ASAP7_75t_L g10679 ( 
.A1(n_8511),
.A2(n_7681),
.B1(n_7376),
.B2(n_7010),
.Y(n_10679)
);

BUFx12f_ASAP7_75t_L g10680 ( 
.A(n_8504),
.Y(n_10680)
);

AO21x1_ASAP7_75t_L g10681 ( 
.A1(n_8400),
.A2(n_7337),
.B(n_7330),
.Y(n_10681)
);

BUFx6f_ASAP7_75t_L g10682 ( 
.A(n_8211),
.Y(n_10682)
);

OAI21x1_ASAP7_75t_L g10683 ( 
.A1(n_8839),
.A2(n_7068),
.B(n_7062),
.Y(n_10683)
);

INVx1_ASAP7_75t_L g10684 ( 
.A(n_8600),
.Y(n_10684)
);

OAI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_8980),
.A2(n_7993),
.B(n_7892),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_8601),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_8601),
.Y(n_10687)
);

INVx1_ASAP7_75t_L g10688 ( 
.A(n_8601),
.Y(n_10688)
);

INVx2_ASAP7_75t_SL g10689 ( 
.A(n_9040),
.Y(n_10689)
);

CKINVDCx5p33_ASAP7_75t_R g10690 ( 
.A(n_9370),
.Y(n_10690)
);

AND2x2_ASAP7_75t_L g10691 ( 
.A(n_9567),
.B(n_8037),
.Y(n_10691)
);

INVx1_ASAP7_75t_L g10692 ( 
.A(n_8608),
.Y(n_10692)
);

INVx3_ASAP7_75t_L g10693 ( 
.A(n_8561),
.Y(n_10693)
);

AOI21x1_ASAP7_75t_L g10694 ( 
.A1(n_8145),
.A2(n_7477),
.B(n_7432),
.Y(n_10694)
);

OAI22xp33_ASAP7_75t_SL g10695 ( 
.A1(n_8866),
.A2(n_7483),
.B1(n_7681),
.B2(n_7848),
.Y(n_10695)
);

AO21x1_ASAP7_75t_SL g10696 ( 
.A1(n_8620),
.A2(n_7337),
.B(n_7330),
.Y(n_10696)
);

INVx3_ASAP7_75t_L g10697 ( 
.A(n_8561),
.Y(n_10697)
);

BUFx2_ASAP7_75t_L g10698 ( 
.A(n_8577),
.Y(n_10698)
);

AOI22xp5_ASAP7_75t_L g10699 ( 
.A1(n_8998),
.A2(n_7376),
.B1(n_7010),
.B2(n_7892),
.Y(n_10699)
);

INVx2_ASAP7_75t_L g10700 ( 
.A(n_9259),
.Y(n_10700)
);

INVx1_ASAP7_75t_L g10701 ( 
.A(n_8608),
.Y(n_10701)
);

BUFx10_ASAP7_75t_L g10702 ( 
.A(n_8834),
.Y(n_10702)
);

HB1xp67_ASAP7_75t_L g10703 ( 
.A(n_9474),
.Y(n_10703)
);

CKINVDCx16_ASAP7_75t_R g10704 ( 
.A(n_8257),
.Y(n_10704)
);

OAI21x1_ASAP7_75t_L g10705 ( 
.A1(n_8849),
.A2(n_7068),
.B(n_7062),
.Y(n_10705)
);

BUFx2_ASAP7_75t_L g10706 ( 
.A(n_8577),
.Y(n_10706)
);

INVx4_ASAP7_75t_L g10707 ( 
.A(n_9427),
.Y(n_10707)
);

OAI22xp5_ASAP7_75t_L g10708 ( 
.A1(n_8889),
.A2(n_8647),
.B1(n_8400),
.B2(n_8643),
.Y(n_10708)
);

INVx2_ASAP7_75t_L g10709 ( 
.A(n_9259),
.Y(n_10709)
);

INVx4_ASAP7_75t_L g10710 ( 
.A(n_9427),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_L g10711 ( 
.A(n_8931),
.B(n_7330),
.Y(n_10711)
);

INVx1_ASAP7_75t_L g10712 ( 
.A(n_8608),
.Y(n_10712)
);

HB1xp67_ASAP7_75t_L g10713 ( 
.A(n_9530),
.Y(n_10713)
);

INVx4_ASAP7_75t_L g10714 ( 
.A(n_9427),
.Y(n_10714)
);

AOI22xp33_ASAP7_75t_L g10715 ( 
.A1(n_8370),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10715)
);

INVx2_ASAP7_75t_L g10716 ( 
.A(n_9261),
.Y(n_10716)
);

OAI21x1_ASAP7_75t_L g10717 ( 
.A1(n_9544),
.A2(n_7091),
.B(n_7068),
.Y(n_10717)
);

CKINVDCx14_ASAP7_75t_R g10718 ( 
.A(n_9043),
.Y(n_10718)
);

INVx1_ASAP7_75t_L g10719 ( 
.A(n_8629),
.Y(n_10719)
);

INVx2_ASAP7_75t_L g10720 ( 
.A(n_9261),
.Y(n_10720)
);

OAI21x1_ASAP7_75t_L g10721 ( 
.A1(n_8911),
.A2(n_7092),
.B(n_7091),
.Y(n_10721)
);

CKINVDCx6p67_ASAP7_75t_R g10722 ( 
.A(n_8602),
.Y(n_10722)
);

HB1xp67_ASAP7_75t_L g10723 ( 
.A(n_9530),
.Y(n_10723)
);

BUFx2_ASAP7_75t_SL g10724 ( 
.A(n_8272),
.Y(n_10724)
);

AND2x2_ASAP7_75t_L g10725 ( 
.A(n_8309),
.B(n_8037),
.Y(n_10725)
);

INVx2_ASAP7_75t_L g10726 ( 
.A(n_9261),
.Y(n_10726)
);

AO21x1_ASAP7_75t_SL g10727 ( 
.A1(n_8575),
.A2(n_7337),
.B(n_7226),
.Y(n_10727)
);

INVx1_ASAP7_75t_SL g10728 ( 
.A(n_9010),
.Y(n_10728)
);

INVx2_ASAP7_75t_L g10729 ( 
.A(n_8561),
.Y(n_10729)
);

INVx2_ASAP7_75t_SL g10730 ( 
.A(n_9427),
.Y(n_10730)
);

OR2x6_ASAP7_75t_L g10731 ( 
.A(n_8202),
.B(n_6965),
.Y(n_10731)
);

OA21x2_ASAP7_75t_L g10732 ( 
.A1(n_8706),
.A2(n_7015),
.B(n_7003),
.Y(n_10732)
);

INVx2_ASAP7_75t_SL g10733 ( 
.A(n_9427),
.Y(n_10733)
);

INVx1_ASAP7_75t_L g10734 ( 
.A(n_8629),
.Y(n_10734)
);

BUFx8_ASAP7_75t_L g10735 ( 
.A(n_8674),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_8629),
.Y(n_10736)
);

INVx2_ASAP7_75t_L g10737 ( 
.A(n_8561),
.Y(n_10737)
);

CKINVDCx11_ASAP7_75t_R g10738 ( 
.A(n_8702),
.Y(n_10738)
);

AOI22xp33_ASAP7_75t_SL g10739 ( 
.A1(n_8866),
.A2(n_7483),
.B1(n_7795),
.B2(n_7739),
.Y(n_10739)
);

INVx2_ASAP7_75t_L g10740 ( 
.A(n_9249),
.Y(n_10740)
);

INVx1_ASAP7_75t_L g10741 ( 
.A(n_8660),
.Y(n_10741)
);

INVx6_ASAP7_75t_L g10742 ( 
.A(n_8704),
.Y(n_10742)
);

HB1xp67_ASAP7_75t_L g10743 ( 
.A(n_9530),
.Y(n_10743)
);

INVx1_ASAP7_75t_SL g10744 ( 
.A(n_9034),
.Y(n_10744)
);

INVx2_ASAP7_75t_L g10745 ( 
.A(n_9249),
.Y(n_10745)
);

AOI22xp33_ASAP7_75t_SL g10746 ( 
.A1(n_8866),
.A2(n_7483),
.B1(n_7795),
.B2(n_7739),
.Y(n_10746)
);

OAI21xp33_ASAP7_75t_L g10747 ( 
.A1(n_8575),
.A2(n_7047),
.B(n_7578),
.Y(n_10747)
);

INVx2_ASAP7_75t_L g10748 ( 
.A(n_9249),
.Y(n_10748)
);

INVx2_ASAP7_75t_L g10749 ( 
.A(n_9257),
.Y(n_10749)
);

CKINVDCx20_ASAP7_75t_R g10750 ( 
.A(n_9520),
.Y(n_10750)
);

AOI22xp33_ASAP7_75t_L g10751 ( 
.A1(n_8486),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10751)
);

INVx2_ASAP7_75t_L g10752 ( 
.A(n_9257),
.Y(n_10752)
);

BUFx4_ASAP7_75t_SL g10753 ( 
.A(n_9049),
.Y(n_10753)
);

CKINVDCx6p67_ASAP7_75t_R g10754 ( 
.A(n_8602),
.Y(n_10754)
);

INVx3_ASAP7_75t_L g10755 ( 
.A(n_9077),
.Y(n_10755)
);

CKINVDCx5p33_ASAP7_75t_R g10756 ( 
.A(n_9520),
.Y(n_10756)
);

AOI22xp33_ASAP7_75t_L g10757 ( 
.A1(n_8486),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10757)
);

AOI22xp33_ASAP7_75t_SL g10758 ( 
.A1(n_8143),
.A2(n_7483),
.B1(n_7866),
.B2(n_7739),
.Y(n_10758)
);

BUFx6f_ASAP7_75t_SL g10759 ( 
.A(n_8630),
.Y(n_10759)
);

HB1xp67_ASAP7_75t_L g10760 ( 
.A(n_8221),
.Y(n_10760)
);

AOI21x1_ASAP7_75t_L g10761 ( 
.A1(n_8145),
.A2(n_7502),
.B(n_7477),
.Y(n_10761)
);

INVx1_ASAP7_75t_L g10762 ( 
.A(n_8660),
.Y(n_10762)
);

NOR2xp33_ASAP7_75t_L g10763 ( 
.A(n_8834),
.B(n_7312),
.Y(n_10763)
);

AO21x1_ASAP7_75t_SL g10764 ( 
.A1(n_8667),
.A2(n_7226),
.B(n_7221),
.Y(n_10764)
);

AND2x2_ASAP7_75t_L g10765 ( 
.A(n_8309),
.B(n_8037),
.Y(n_10765)
);

INVx1_ASAP7_75t_L g10766 ( 
.A(n_8660),
.Y(n_10766)
);

INVx1_ASAP7_75t_L g10767 ( 
.A(n_8670),
.Y(n_10767)
);

OAI21x1_ASAP7_75t_L g10768 ( 
.A1(n_9544),
.A2(n_7092),
.B(n_7091),
.Y(n_10768)
);

BUFx3_ASAP7_75t_L g10769 ( 
.A(n_9427),
.Y(n_10769)
);

AND2x2_ASAP7_75t_L g10770 ( 
.A(n_8309),
.B(n_8042),
.Y(n_10770)
);

INVx2_ASAP7_75t_L g10771 ( 
.A(n_9257),
.Y(n_10771)
);

BUFx6f_ASAP7_75t_L g10772 ( 
.A(n_8211),
.Y(n_10772)
);

CKINVDCx5p33_ASAP7_75t_R g10773 ( 
.A(n_9049),
.Y(n_10773)
);

AOI22xp33_ASAP7_75t_L g10774 ( 
.A1(n_8617),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10774)
);

AOI22xp33_ASAP7_75t_L g10775 ( 
.A1(n_8617),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10775)
);

AND2x2_ASAP7_75t_L g10776 ( 
.A(n_8312),
.B(n_8042),
.Y(n_10776)
);

CKINVDCx11_ASAP7_75t_R g10777 ( 
.A(n_8272),
.Y(n_10777)
);

HB1xp67_ASAP7_75t_L g10778 ( 
.A(n_8221),
.Y(n_10778)
);

INVx1_ASAP7_75t_L g10779 ( 
.A(n_8670),
.Y(n_10779)
);

OAI22xp33_ASAP7_75t_L g10780 ( 
.A1(n_8551),
.A2(n_8049),
.B1(n_8023),
.B2(n_7848),
.Y(n_10780)
);

INVx2_ASAP7_75t_L g10781 ( 
.A(n_8512),
.Y(n_10781)
);

OAI22xp5_ASAP7_75t_L g10782 ( 
.A1(n_8889),
.A2(n_7304),
.B1(n_7513),
.B2(n_6998),
.Y(n_10782)
);

NAND2xp5_ASAP7_75t_L g10783 ( 
.A(n_8931),
.B(n_7047),
.Y(n_10783)
);

AOI21x1_ASAP7_75t_L g10784 ( 
.A1(n_8145),
.A2(n_7519),
.B(n_7502),
.Y(n_10784)
);

INVx1_ASAP7_75t_L g10785 ( 
.A(n_8670),
.Y(n_10785)
);

OAI22xp33_ASAP7_75t_L g10786 ( 
.A1(n_8551),
.A2(n_8023),
.B1(n_8049),
.B2(n_7483),
.Y(n_10786)
);

AOI21x1_ASAP7_75t_L g10787 ( 
.A1(n_8156),
.A2(n_7519),
.B(n_7502),
.Y(n_10787)
);

INVx3_ASAP7_75t_L g10788 ( 
.A(n_9077),
.Y(n_10788)
);

AND2x4_ASAP7_75t_L g10789 ( 
.A(n_8720),
.B(n_9144),
.Y(n_10789)
);

INVx1_ASAP7_75t_L g10790 ( 
.A(n_8676),
.Y(n_10790)
);

AOI22xp33_ASAP7_75t_SL g10791 ( 
.A1(n_8143),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_10791)
);

OR2x2_ASAP7_75t_L g10792 ( 
.A(n_8301),
.B(n_7209),
.Y(n_10792)
);

INVx2_ASAP7_75t_SL g10793 ( 
.A(n_9427),
.Y(n_10793)
);

INVx1_ASAP7_75t_L g10794 ( 
.A(n_8676),
.Y(n_10794)
);

INVx2_ASAP7_75t_L g10795 ( 
.A(n_8512),
.Y(n_10795)
);

AND2x2_ASAP7_75t_L g10796 ( 
.A(n_8312),
.B(n_8042),
.Y(n_10796)
);

OR2x2_ASAP7_75t_L g10797 ( 
.A(n_8301),
.B(n_7209),
.Y(n_10797)
);

INVx1_ASAP7_75t_L g10798 ( 
.A(n_8676),
.Y(n_10798)
);

BUFx6f_ASAP7_75t_L g10799 ( 
.A(n_8360),
.Y(n_10799)
);

AOI22xp33_ASAP7_75t_L g10800 ( 
.A1(n_9514),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10800)
);

OAI22xp33_ASAP7_75t_L g10801 ( 
.A1(n_8604),
.A2(n_9000),
.B1(n_8745),
.B2(n_8529),
.Y(n_10801)
);

INVx1_ASAP7_75t_L g10802 ( 
.A(n_8683),
.Y(n_10802)
);

OAI21x1_ASAP7_75t_L g10803 ( 
.A1(n_8911),
.A2(n_7092),
.B(n_7091),
.Y(n_10803)
);

INVx1_ASAP7_75t_L g10804 ( 
.A(n_8683),
.Y(n_10804)
);

HB1xp67_ASAP7_75t_L g10805 ( 
.A(n_8236),
.Y(n_10805)
);

INVx1_ASAP7_75t_L g10806 ( 
.A(n_8683),
.Y(n_10806)
);

OR2x2_ASAP7_75t_L g10807 ( 
.A(n_8311),
.B(n_7209),
.Y(n_10807)
);

OAI21x1_ASAP7_75t_SL g10808 ( 
.A1(n_8143),
.A2(n_7080),
.B(n_7065),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_8685),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_8685),
.Y(n_10810)
);

AOI22xp5_ASAP7_75t_L g10811 ( 
.A1(n_8998),
.A2(n_7892),
.B1(n_6998),
.B2(n_6962),
.Y(n_10811)
);

INVx1_ASAP7_75t_L g10812 ( 
.A(n_8685),
.Y(n_10812)
);

INVx1_ASAP7_75t_L g10813 ( 
.A(n_8689),
.Y(n_10813)
);

AND2x4_ASAP7_75t_L g10814 ( 
.A(n_8720),
.B(n_8042),
.Y(n_10814)
);

INVx1_ASAP7_75t_L g10815 ( 
.A(n_8689),
.Y(n_10815)
);

AOI22xp33_ASAP7_75t_L g10816 ( 
.A1(n_9514),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10816)
);

BUFx4f_ASAP7_75t_SL g10817 ( 
.A(n_9034),
.Y(n_10817)
);

AOI22xp33_ASAP7_75t_L g10818 ( 
.A1(n_9514),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_8689),
.Y(n_10819)
);

CKINVDCx5p33_ASAP7_75t_R g10820 ( 
.A(n_9356),
.Y(n_10820)
);

AND2x2_ASAP7_75t_L g10821 ( 
.A(n_8312),
.B(n_8068),
.Y(n_10821)
);

BUFx10_ASAP7_75t_L g10822 ( 
.A(n_8704),
.Y(n_10822)
);

INVx1_ASAP7_75t_L g10823 ( 
.A(n_8696),
.Y(n_10823)
);

INVx2_ASAP7_75t_L g10824 ( 
.A(n_8512),
.Y(n_10824)
);

AOI22xp33_ASAP7_75t_L g10825 ( 
.A1(n_9514),
.A2(n_7230),
.B1(n_7286),
.B2(n_7245),
.Y(n_10825)
);

INVx2_ASAP7_75t_L g10826 ( 
.A(n_8512),
.Y(n_10826)
);

INVx2_ASAP7_75t_L g10827 ( 
.A(n_8512),
.Y(n_10827)
);

INVx1_ASAP7_75t_L g10828 ( 
.A(n_8696),
.Y(n_10828)
);

HB1xp67_ASAP7_75t_L g10829 ( 
.A(n_8236),
.Y(n_10829)
);

INVx1_ASAP7_75t_L g10830 ( 
.A(n_8696),
.Y(n_10830)
);

NAND2x1p5_ASAP7_75t_L g10831 ( 
.A(n_9508),
.B(n_7834),
.Y(n_10831)
);

INVx2_ASAP7_75t_L g10832 ( 
.A(n_8138),
.Y(n_10832)
);

INVx1_ASAP7_75t_L g10833 ( 
.A(n_8701),
.Y(n_10833)
);

NAND2x1p5_ASAP7_75t_L g10834 ( 
.A(n_9508),
.B(n_7834),
.Y(n_10834)
);

AND2x2_ASAP7_75t_L g10835 ( 
.A(n_8482),
.B(n_8068),
.Y(n_10835)
);

INVx2_ASAP7_75t_L g10836 ( 
.A(n_8138),
.Y(n_10836)
);

OAI22x1_ASAP7_75t_L g10837 ( 
.A1(n_8485),
.A2(n_7859),
.B1(n_7258),
.B2(n_7259),
.Y(n_10837)
);

BUFx2_ASAP7_75t_L g10838 ( 
.A(n_8577),
.Y(n_10838)
);

AO21x1_ASAP7_75t_SL g10839 ( 
.A1(n_8667),
.A2(n_7226),
.B(n_7221),
.Y(n_10839)
);

NAND2xp5_ASAP7_75t_L g10840 ( 
.A(n_9023),
.B(n_7047),
.Y(n_10840)
);

INVx1_ASAP7_75t_L g10841 ( 
.A(n_8701),
.Y(n_10841)
);

OAI22xp33_ASAP7_75t_L g10842 ( 
.A1(n_8604),
.A2(n_7304),
.B1(n_7356),
.B2(n_7351),
.Y(n_10842)
);

AOI22xp33_ASAP7_75t_L g10843 ( 
.A1(n_9514),
.A2(n_7286),
.B1(n_7332),
.B2(n_7296),
.Y(n_10843)
);

OAI21x1_ASAP7_75t_L g10844 ( 
.A1(n_8405),
.A2(n_7092),
.B(n_7091),
.Y(n_10844)
);

INVxp67_ASAP7_75t_L g10845 ( 
.A(n_8606),
.Y(n_10845)
);

AOI22xp33_ASAP7_75t_L g10846 ( 
.A1(n_9543),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10846)
);

BUFx8_ASAP7_75t_L g10847 ( 
.A(n_8715),
.Y(n_10847)
);

INVx2_ASAP7_75t_L g10848 ( 
.A(n_8138),
.Y(n_10848)
);

AO21x1_ASAP7_75t_L g10849 ( 
.A1(n_9345),
.A2(n_7228),
.B(n_7221),
.Y(n_10849)
);

BUFx3_ASAP7_75t_L g10850 ( 
.A(n_8968),
.Y(n_10850)
);

INVx1_ASAP7_75t_L g10851 ( 
.A(n_8701),
.Y(n_10851)
);

BUFx2_ASAP7_75t_L g10852 ( 
.A(n_8577),
.Y(n_10852)
);

INVx1_ASAP7_75t_L g10853 ( 
.A(n_8710),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_8710),
.Y(n_10854)
);

OAI21x1_ASAP7_75t_L g10855 ( 
.A1(n_8911),
.A2(n_7092),
.B(n_7091),
.Y(n_10855)
);

AND2x2_ASAP7_75t_L g10856 ( 
.A(n_8482),
.B(n_8068),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_8710),
.Y(n_10857)
);

INVx4_ASAP7_75t_L g10858 ( 
.A(n_9111),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_8719),
.Y(n_10859)
);

OAI22xp5_ASAP7_75t_L g10860 ( 
.A1(n_8606),
.A2(n_7304),
.B1(n_7513),
.B2(n_6962),
.Y(n_10860)
);

BUFx4f_ASAP7_75t_SL g10861 ( 
.A(n_9204),
.Y(n_10861)
);

AOI22xp33_ASAP7_75t_SL g10862 ( 
.A1(n_8138),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_10862)
);

NAND2x1p5_ASAP7_75t_L g10863 ( 
.A(n_9512),
.B(n_7834),
.Y(n_10863)
);

BUFx6f_ASAP7_75t_L g10864 ( 
.A(n_8360),
.Y(n_10864)
);

AOI21x1_ASAP7_75t_L g10865 ( 
.A1(n_8156),
.A2(n_8157),
.B(n_9093),
.Y(n_10865)
);

BUFx2_ASAP7_75t_L g10866 ( 
.A(n_8577),
.Y(n_10866)
);

AO21x2_ASAP7_75t_L g10867 ( 
.A1(n_8189),
.A2(n_6934),
.B(n_6932),
.Y(n_10867)
);

INVx1_ASAP7_75t_L g10868 ( 
.A(n_8719),
.Y(n_10868)
);

INVx2_ASAP7_75t_L g10869 ( 
.A(n_8138),
.Y(n_10869)
);

BUFx3_ASAP7_75t_L g10870 ( 
.A(n_9111),
.Y(n_10870)
);

HB1xp67_ASAP7_75t_L g10871 ( 
.A(n_8292),
.Y(n_10871)
);

NAND2xp5_ASAP7_75t_L g10872 ( 
.A(n_9023),
.B(n_9030),
.Y(n_10872)
);

AND2x2_ASAP7_75t_L g10873 ( 
.A(n_8482),
.B(n_8068),
.Y(n_10873)
);

INVx1_ASAP7_75t_L g10874 ( 
.A(n_8719),
.Y(n_10874)
);

INVx1_ASAP7_75t_L g10875 ( 
.A(n_8721),
.Y(n_10875)
);

INVx1_ASAP7_75t_SL g10876 ( 
.A(n_9204),
.Y(n_10876)
);

INVx2_ASAP7_75t_SL g10877 ( 
.A(n_8246),
.Y(n_10877)
);

INVx1_ASAP7_75t_L g10878 ( 
.A(n_8721),
.Y(n_10878)
);

BUFx6f_ASAP7_75t_L g10879 ( 
.A(n_8360),
.Y(n_10879)
);

INVx2_ASAP7_75t_L g10880 ( 
.A(n_8138),
.Y(n_10880)
);

HB1xp67_ASAP7_75t_L g10881 ( 
.A(n_8292),
.Y(n_10881)
);

AOI22xp33_ASAP7_75t_L g10882 ( 
.A1(n_9543),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10882)
);

INVx6_ASAP7_75t_L g10883 ( 
.A(n_8704),
.Y(n_10883)
);

INVx2_ASAP7_75t_L g10884 ( 
.A(n_8144),
.Y(n_10884)
);

INVx11_ASAP7_75t_L g10885 ( 
.A(n_9111),
.Y(n_10885)
);

NOR2xp33_ASAP7_75t_L g10886 ( 
.A(n_8492),
.B(n_7312),
.Y(n_10886)
);

INVx2_ASAP7_75t_L g10887 ( 
.A(n_8144),
.Y(n_10887)
);

INVx2_ASAP7_75t_L g10888 ( 
.A(n_8144),
.Y(n_10888)
);

INVx4_ASAP7_75t_L g10889 ( 
.A(n_9414),
.Y(n_10889)
);

AND2x2_ASAP7_75t_L g10890 ( 
.A(n_8213),
.B(n_8090),
.Y(n_10890)
);

INVx1_ASAP7_75t_L g10891 ( 
.A(n_8721),
.Y(n_10891)
);

AOI22xp33_ASAP7_75t_L g10892 ( 
.A1(n_9543),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10892)
);

NAND2x1p5_ASAP7_75t_L g10893 ( 
.A(n_9512),
.B(n_7834),
.Y(n_10893)
);

INVx1_ASAP7_75t_L g10894 ( 
.A(n_8723),
.Y(n_10894)
);

OAI22xp33_ASAP7_75t_L g10895 ( 
.A1(n_9000),
.A2(n_7356),
.B1(n_7366),
.B2(n_7351),
.Y(n_10895)
);

INVx1_ASAP7_75t_L g10896 ( 
.A(n_8723),
.Y(n_10896)
);

AO21x1_ASAP7_75t_L g10897 ( 
.A1(n_9345),
.A2(n_7255),
.B(n_7228),
.Y(n_10897)
);

INVx1_ASAP7_75t_L g10898 ( 
.A(n_8723),
.Y(n_10898)
);

CKINVDCx20_ASAP7_75t_R g10899 ( 
.A(n_9276),
.Y(n_10899)
);

OAI21x1_ASAP7_75t_L g10900 ( 
.A1(n_8405),
.A2(n_7141),
.B(n_7092),
.Y(n_10900)
);

INVxp67_ASAP7_75t_L g10901 ( 
.A(n_8669),
.Y(n_10901)
);

INVx1_ASAP7_75t_L g10902 ( 
.A(n_8730),
.Y(n_10902)
);

OAI22xp5_ASAP7_75t_L g10903 ( 
.A1(n_8669),
.A2(n_7513),
.B1(n_7767),
.B2(n_8030),
.Y(n_10903)
);

OAI22xp5_ASAP7_75t_L g10904 ( 
.A1(n_8755),
.A2(n_7767),
.B1(n_8035),
.B2(n_8030),
.Y(n_10904)
);

INVx1_ASAP7_75t_L g10905 ( 
.A(n_8730),
.Y(n_10905)
);

NAND2x1p5_ASAP7_75t_L g10906 ( 
.A(n_9512),
.B(n_7834),
.Y(n_10906)
);

INVx1_ASAP7_75t_L g10907 ( 
.A(n_8730),
.Y(n_10907)
);

INVx1_ASAP7_75t_L g10908 ( 
.A(n_8743),
.Y(n_10908)
);

NAND2x1p5_ASAP7_75t_L g10909 ( 
.A(n_8151),
.B(n_7834),
.Y(n_10909)
);

AOI22xp33_ASAP7_75t_L g10910 ( 
.A1(n_9543),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10910)
);

AOI22xp33_ASAP7_75t_SL g10911 ( 
.A1(n_8144),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_10911)
);

CKINVDCx5p33_ASAP7_75t_R g10912 ( 
.A(n_9356),
.Y(n_10912)
);

AOI22xp33_ASAP7_75t_L g10913 ( 
.A1(n_9543),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10913)
);

OAI21x1_ASAP7_75t_SL g10914 ( 
.A1(n_8151),
.A2(n_7402),
.B(n_8090),
.Y(n_10914)
);

INVx1_ASAP7_75t_L g10915 ( 
.A(n_8743),
.Y(n_10915)
);

OR2x6_ASAP7_75t_L g10916 ( 
.A(n_8202),
.B(n_6965),
.Y(n_10916)
);

INVx1_ASAP7_75t_L g10917 ( 
.A(n_8743),
.Y(n_10917)
);

INVx2_ASAP7_75t_SL g10918 ( 
.A(n_8246),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_8758),
.Y(n_10919)
);

INVx2_ASAP7_75t_L g10920 ( 
.A(n_8144),
.Y(n_10920)
);

AO21x2_ASAP7_75t_L g10921 ( 
.A1(n_8189),
.A2(n_6934),
.B(n_6932),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_8758),
.Y(n_10922)
);

BUFx2_ASAP7_75t_R g10923 ( 
.A(n_8956),
.Y(n_10923)
);

AND2x2_ASAP7_75t_L g10924 ( 
.A(n_8213),
.B(n_8090),
.Y(n_10924)
);

AOI22xp33_ASAP7_75t_L g10925 ( 
.A1(n_9002),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10925)
);

BUFx6f_ASAP7_75t_L g10926 ( 
.A(n_8360),
.Y(n_10926)
);

AOI22xp33_ASAP7_75t_L g10927 ( 
.A1(n_9002),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10927)
);

INVx1_ASAP7_75t_L g10928 ( 
.A(n_8758),
.Y(n_10928)
);

OA21x2_ASAP7_75t_L g10929 ( 
.A1(n_9062),
.A2(n_7015),
.B(n_7003),
.Y(n_10929)
);

NAND2x1p5_ASAP7_75t_L g10930 ( 
.A(n_8151),
.B(n_7834),
.Y(n_10930)
);

INVx1_ASAP7_75t_L g10931 ( 
.A(n_8763),
.Y(n_10931)
);

BUFx6f_ASAP7_75t_L g10932 ( 
.A(n_8360),
.Y(n_10932)
);

OAI22xp5_ASAP7_75t_SL g10933 ( 
.A1(n_8492),
.A2(n_7312),
.B1(n_7382),
.B2(n_7326),
.Y(n_10933)
);

AOI22xp33_ASAP7_75t_SL g10934 ( 
.A1(n_8144),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_10934)
);

INVx2_ASAP7_75t_L g10935 ( 
.A(n_8940),
.Y(n_10935)
);

BUFx6f_ASAP7_75t_L g10936 ( 
.A(n_8360),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_8763),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_8763),
.Y(n_10938)
);

INVx2_ASAP7_75t_L g10939 ( 
.A(n_8940),
.Y(n_10939)
);

AO21x1_ASAP7_75t_L g10940 ( 
.A1(n_8909),
.A2(n_7255),
.B(n_7228),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_8786),
.Y(n_10941)
);

INVx2_ASAP7_75t_L g10942 ( 
.A(n_8940),
.Y(n_10942)
);

AND2x2_ASAP7_75t_L g10943 ( 
.A(n_8213),
.B(n_8090),
.Y(n_10943)
);

INVx1_ASAP7_75t_L g10944 ( 
.A(n_8786),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_8786),
.Y(n_10945)
);

INVx2_ASAP7_75t_L g10946 ( 
.A(n_8948),
.Y(n_10946)
);

INVx2_ASAP7_75t_L g10947 ( 
.A(n_8948),
.Y(n_10947)
);

BUFx3_ASAP7_75t_L g10948 ( 
.A(n_9414),
.Y(n_10948)
);

OA21x2_ASAP7_75t_L g10949 ( 
.A1(n_9062),
.A2(n_7015),
.B(n_7003),
.Y(n_10949)
);

INVx1_ASAP7_75t_L g10950 ( 
.A(n_8790),
.Y(n_10950)
);

INVx1_ASAP7_75t_L g10951 ( 
.A(n_8790),
.Y(n_10951)
);

INVx5_ASAP7_75t_L g10952 ( 
.A(n_9358),
.Y(n_10952)
);

INVx1_ASAP7_75t_L g10953 ( 
.A(n_8790),
.Y(n_10953)
);

CKINVDCx20_ASAP7_75t_R g10954 ( 
.A(n_9276),
.Y(n_10954)
);

INVx1_ASAP7_75t_L g10955 ( 
.A(n_8791),
.Y(n_10955)
);

OR2x2_ASAP7_75t_L g10956 ( 
.A(n_8311),
.B(n_7921),
.Y(n_10956)
);

INVx4_ASAP7_75t_L g10957 ( 
.A(n_9414),
.Y(n_10957)
);

AOI22xp33_ASAP7_75t_L g10958 ( 
.A1(n_8653),
.A2(n_8872),
.B1(n_8880),
.B2(n_9550),
.Y(n_10958)
);

AND2x4_ASAP7_75t_L g10959 ( 
.A(n_9144),
.B(n_8093),
.Y(n_10959)
);

BUFx2_ASAP7_75t_SL g10960 ( 
.A(n_8630),
.Y(n_10960)
);

BUFx3_ASAP7_75t_L g10961 ( 
.A(n_8630),
.Y(n_10961)
);

INVx3_ASAP7_75t_L g10962 ( 
.A(n_9077),
.Y(n_10962)
);

INVx2_ASAP7_75t_L g10963 ( 
.A(n_8948),
.Y(n_10963)
);

HB1xp67_ASAP7_75t_L g10964 ( 
.A(n_8359),
.Y(n_10964)
);

AND2x2_ASAP7_75t_L g10965 ( 
.A(n_8890),
.B(n_8093),
.Y(n_10965)
);

AOI22xp33_ASAP7_75t_SL g10966 ( 
.A1(n_8297),
.A2(n_8640),
.B1(n_8621),
.B2(n_9125),
.Y(n_10966)
);

INVx2_ASAP7_75t_L g10967 ( 
.A(n_9232),
.Y(n_10967)
);

INVx1_ASAP7_75t_L g10968 ( 
.A(n_8791),
.Y(n_10968)
);

INVx6_ASAP7_75t_L g10969 ( 
.A(n_8704),
.Y(n_10969)
);

INVx1_ASAP7_75t_SL g10970 ( 
.A(n_9291),
.Y(n_10970)
);

INVx1_ASAP7_75t_SL g10971 ( 
.A(n_9291),
.Y(n_10971)
);

OAI21xp5_ASAP7_75t_L g10972 ( 
.A1(n_8901),
.A2(n_7143),
.B(n_7751),
.Y(n_10972)
);

AOI22xp33_ASAP7_75t_L g10973 ( 
.A1(n_8653),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10973)
);

BUFx2_ASAP7_75t_L g10974 ( 
.A(n_8572),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_8791),
.Y(n_10975)
);

INVx3_ASAP7_75t_L g10976 ( 
.A(n_8164),
.Y(n_10976)
);

INVx1_ASAP7_75t_L g10977 ( 
.A(n_8804),
.Y(n_10977)
);

OAI22xp5_ASAP7_75t_L g10978 ( 
.A1(n_8755),
.A2(n_8030),
.B1(n_8052),
.B2(n_8035),
.Y(n_10978)
);

INVx1_ASAP7_75t_L g10979 ( 
.A(n_8804),
.Y(n_10979)
);

OR2x2_ASAP7_75t_L g10980 ( 
.A(n_8131),
.B(n_7921),
.Y(n_10980)
);

OAI21x1_ASAP7_75t_L g10981 ( 
.A1(n_8405),
.A2(n_7150),
.B(n_7141),
.Y(n_10981)
);

INVx1_ASAP7_75t_L g10982 ( 
.A(n_8804),
.Y(n_10982)
);

INVx1_ASAP7_75t_L g10983 ( 
.A(n_8970),
.Y(n_10983)
);

INVx1_ASAP7_75t_L g10984 ( 
.A(n_8970),
.Y(n_10984)
);

BUFx6f_ASAP7_75t_L g10985 ( 
.A(n_8360),
.Y(n_10985)
);

INVx2_ASAP7_75t_L g10986 ( 
.A(n_9232),
.Y(n_10986)
);

INVx1_ASAP7_75t_L g10987 ( 
.A(n_8970),
.Y(n_10987)
);

INVx2_ASAP7_75t_L g10988 ( 
.A(n_9232),
.Y(n_10988)
);

INVx2_ASAP7_75t_SL g10989 ( 
.A(n_8246),
.Y(n_10989)
);

OAI21x1_ASAP7_75t_L g10990 ( 
.A1(n_8371),
.A2(n_7150),
.B(n_7141),
.Y(n_10990)
);

AOI22xp33_ASAP7_75t_L g10991 ( 
.A1(n_8872),
.A2(n_7296),
.B1(n_7372),
.B2(n_7332),
.Y(n_10991)
);

AOI21x1_ASAP7_75t_L g10992 ( 
.A1(n_8156),
.A2(n_7534),
.B(n_7519),
.Y(n_10992)
);

INVx1_ASAP7_75t_L g10993 ( 
.A(n_8989),
.Y(n_10993)
);

BUFx2_ASAP7_75t_L g10994 ( 
.A(n_8572),
.Y(n_10994)
);

AOI21x1_ASAP7_75t_L g10995 ( 
.A1(n_8156),
.A2(n_7535),
.B(n_7534),
.Y(n_10995)
);

INVx1_ASAP7_75t_L g10996 ( 
.A(n_8989),
.Y(n_10996)
);

BUFx6f_ASAP7_75t_L g10997 ( 
.A(n_8360),
.Y(n_10997)
);

OAI21x1_ASAP7_75t_L g10998 ( 
.A1(n_8371),
.A2(n_7150),
.B(n_7141),
.Y(n_10998)
);

BUFx3_ASAP7_75t_L g10999 ( 
.A(n_8780),
.Y(n_10999)
);

AO21x1_ASAP7_75t_SL g11000 ( 
.A1(n_9368),
.A2(n_7287),
.B(n_7271),
.Y(n_11000)
);

OAI21x1_ASAP7_75t_L g11001 ( 
.A1(n_8371),
.A2(n_7150),
.B(n_7141),
.Y(n_11001)
);

INVx2_ASAP7_75t_L g11002 ( 
.A(n_9233),
.Y(n_11002)
);

AOI22xp5_ASAP7_75t_L g11003 ( 
.A1(n_9171),
.A2(n_7533),
.B1(n_7751),
.B2(n_7720),
.Y(n_11003)
);

AOI21xp5_ASAP7_75t_L g11004 ( 
.A1(n_8437),
.A2(n_7751),
.B(n_7806),
.Y(n_11004)
);

INVx6_ASAP7_75t_L g11005 ( 
.A(n_8704),
.Y(n_11005)
);

INVx1_ASAP7_75t_L g11006 ( 
.A(n_8989),
.Y(n_11006)
);

INVx1_ASAP7_75t_L g11007 ( 
.A(n_9007),
.Y(n_11007)
);

INVx1_ASAP7_75t_L g11008 ( 
.A(n_9007),
.Y(n_11008)
);

INVx2_ASAP7_75t_L g11009 ( 
.A(n_9233),
.Y(n_11009)
);

INVx1_ASAP7_75t_L g11010 ( 
.A(n_9007),
.Y(n_11010)
);

INVx1_ASAP7_75t_L g11011 ( 
.A(n_9016),
.Y(n_11011)
);

INVx1_ASAP7_75t_L g11012 ( 
.A(n_9016),
.Y(n_11012)
);

AND2x2_ASAP7_75t_L g11013 ( 
.A(n_8890),
.B(n_8093),
.Y(n_11013)
);

NAND2x1_ASAP7_75t_L g11014 ( 
.A(n_8260),
.B(n_8093),
.Y(n_11014)
);

INVx2_ASAP7_75t_L g11015 ( 
.A(n_9233),
.Y(n_11015)
);

INVx1_ASAP7_75t_L g11016 ( 
.A(n_9016),
.Y(n_11016)
);

AND2x2_ASAP7_75t_L g11017 ( 
.A(n_8890),
.B(n_8098),
.Y(n_11017)
);

BUFx2_ASAP7_75t_L g11018 ( 
.A(n_8572),
.Y(n_11018)
);

BUFx3_ASAP7_75t_L g11019 ( 
.A(n_8780),
.Y(n_11019)
);

INVx6_ASAP7_75t_L g11020 ( 
.A(n_8704),
.Y(n_11020)
);

INVx6_ASAP7_75t_L g11021 ( 
.A(n_8711),
.Y(n_11021)
);

INVx1_ASAP7_75t_L g11022 ( 
.A(n_9018),
.Y(n_11022)
);

INVx1_ASAP7_75t_SL g11023 ( 
.A(n_9303),
.Y(n_11023)
);

INVx2_ASAP7_75t_L g11024 ( 
.A(n_10458),
.Y(n_11024)
);

HB1xp67_ASAP7_75t_L g11025 ( 
.A(n_9677),
.Y(n_11025)
);

NAND2xp5_ASAP7_75t_L g11026 ( 
.A(n_9820),
.B(n_10050),
.Y(n_11026)
);

INVx1_ASAP7_75t_L g11027 ( 
.A(n_9581),
.Y(n_11027)
);

INVx2_ASAP7_75t_L g11028 ( 
.A(n_10458),
.Y(n_11028)
);

INVx2_ASAP7_75t_L g11029 ( 
.A(n_10458),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_9581),
.Y(n_11030)
);

OA21x2_ASAP7_75t_L g11031 ( 
.A1(n_10187),
.A2(n_8568),
.B(n_8208),
.Y(n_11031)
);

AND2x4_ASAP7_75t_L g11032 ( 
.A(n_9687),
.B(n_8246),
.Y(n_11032)
);

NOR2xp33_ASAP7_75t_L g11033 ( 
.A(n_9677),
.B(n_9303),
.Y(n_11033)
);

AOI222xp33_ASAP7_75t_L g11034 ( 
.A1(n_10557),
.A2(n_9017),
.B1(n_9008),
.B2(n_8901),
.C1(n_8860),
.C2(n_9563),
.Y(n_11034)
);

INVx2_ASAP7_75t_L g11035 ( 
.A(n_10458),
.Y(n_11035)
);

INVx2_ASAP7_75t_L g11036 ( 
.A(n_10458),
.Y(n_11036)
);

INVx1_ASAP7_75t_L g11037 ( 
.A(n_9582),
.Y(n_11037)
);

CKINVDCx5p33_ASAP7_75t_R g11038 ( 
.A(n_9821),
.Y(n_11038)
);

BUFx6f_ASAP7_75t_L g11039 ( 
.A(n_9657),
.Y(n_11039)
);

HB1xp67_ASAP7_75t_L g11040 ( 
.A(n_10147),
.Y(n_11040)
);

BUFx6f_ASAP7_75t_L g11041 ( 
.A(n_9657),
.Y(n_11041)
);

AOI21x1_ASAP7_75t_L g11042 ( 
.A1(n_9758),
.A2(n_8992),
.B(n_8978),
.Y(n_11042)
);

INVx2_ASAP7_75t_L g11043 ( 
.A(n_10458),
.Y(n_11043)
);

OAI21xp5_ASAP7_75t_L g11044 ( 
.A1(n_9882),
.A2(n_8593),
.B(n_8569),
.Y(n_11044)
);

NAND2xp5_ASAP7_75t_L g11045 ( 
.A(n_10187),
.B(n_9075),
.Y(n_11045)
);

AO21x2_ASAP7_75t_L g11046 ( 
.A1(n_9654),
.A2(n_8908),
.B(n_9407),
.Y(n_11046)
);

BUFx3_ASAP7_75t_L g11047 ( 
.A(n_9947),
.Y(n_11047)
);

AOI22xp33_ASAP7_75t_L g11048 ( 
.A1(n_9903),
.A2(n_8880),
.B1(n_9135),
.B2(n_9131),
.Y(n_11048)
);

INVx1_ASAP7_75t_L g11049 ( 
.A(n_9582),
.Y(n_11049)
);

INVx3_ASAP7_75t_L g11050 ( 
.A(n_9687),
.Y(n_11050)
);

INVx2_ASAP7_75t_L g11051 ( 
.A(n_10517),
.Y(n_11051)
);

BUFx2_ASAP7_75t_L g11052 ( 
.A(n_9799),
.Y(n_11052)
);

INVx1_ASAP7_75t_L g11053 ( 
.A(n_9583),
.Y(n_11053)
);

INVx4_ASAP7_75t_SL g11054 ( 
.A(n_9657),
.Y(n_11054)
);

INVx2_ASAP7_75t_L g11055 ( 
.A(n_10517),
.Y(n_11055)
);

OAI21x1_ASAP7_75t_L g11056 ( 
.A1(n_10143),
.A2(n_8264),
.B(n_8258),
.Y(n_11056)
);

HB1xp67_ASAP7_75t_L g11057 ( 
.A(n_10147),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_9583),
.Y(n_11058)
);

INVx2_ASAP7_75t_L g11059 ( 
.A(n_10517),
.Y(n_11059)
);

INVx1_ASAP7_75t_L g11060 ( 
.A(n_9586),
.Y(n_11060)
);

INVx2_ASAP7_75t_L g11061 ( 
.A(n_10517),
.Y(n_11061)
);

AND2x2_ASAP7_75t_L g11062 ( 
.A(n_10108),
.B(n_8952),
.Y(n_11062)
);

HB1xp67_ASAP7_75t_L g11063 ( 
.A(n_10157),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_9586),
.Y(n_11064)
);

INVx1_ASAP7_75t_L g11065 ( 
.A(n_9593),
.Y(n_11065)
);

HB1xp67_ASAP7_75t_L g11066 ( 
.A(n_10157),
.Y(n_11066)
);

INVx1_ASAP7_75t_L g11067 ( 
.A(n_9593),
.Y(n_11067)
);

INVx2_ASAP7_75t_L g11068 ( 
.A(n_10517),
.Y(n_11068)
);

OA21x2_ASAP7_75t_L g11069 ( 
.A1(n_10407),
.A2(n_8568),
.B(n_8208),
.Y(n_11069)
);

OA21x2_ASAP7_75t_L g11070 ( 
.A1(n_10407),
.A2(n_8568),
.B(n_8208),
.Y(n_11070)
);

INVx3_ASAP7_75t_L g11071 ( 
.A(n_9687),
.Y(n_11071)
);

INVx1_ASAP7_75t_SL g11072 ( 
.A(n_10274),
.Y(n_11072)
);

HB1xp67_ASAP7_75t_L g11073 ( 
.A(n_10171),
.Y(n_11073)
);

INVx2_ASAP7_75t_L g11074 ( 
.A(n_10517),
.Y(n_11074)
);

HB1xp67_ASAP7_75t_L g11075 ( 
.A(n_10171),
.Y(n_11075)
);

HB1xp67_ASAP7_75t_L g11076 ( 
.A(n_10215),
.Y(n_11076)
);

OR2x2_ASAP7_75t_L g11077 ( 
.A(n_10872),
.B(n_8314),
.Y(n_11077)
);

BUFx6f_ASAP7_75t_L g11078 ( 
.A(n_9665),
.Y(n_11078)
);

HB1xp67_ASAP7_75t_L g11079 ( 
.A(n_10215),
.Y(n_11079)
);

INVx1_ASAP7_75t_L g11080 ( 
.A(n_9596),
.Y(n_11080)
);

OA21x2_ASAP7_75t_L g11081 ( 
.A1(n_9855),
.A2(n_8189),
.B(n_8282),
.Y(n_11081)
);

AOI22xp5_ASAP7_75t_SL g11082 ( 
.A1(n_10347),
.A2(n_7350),
.B1(n_7381),
.B2(n_8806),
.Y(n_11082)
);

OR2x2_ASAP7_75t_L g11083 ( 
.A(n_10872),
.B(n_8314),
.Y(n_11083)
);

INVx2_ASAP7_75t_L g11084 ( 
.A(n_9670),
.Y(n_11084)
);

INVx3_ASAP7_75t_L g11085 ( 
.A(n_9687),
.Y(n_11085)
);

NAND2xp5_ASAP7_75t_L g11086 ( 
.A(n_9688),
.B(n_9075),
.Y(n_11086)
);

INVxp67_ASAP7_75t_L g11087 ( 
.A(n_10487),
.Y(n_11087)
);

INVx2_ASAP7_75t_L g11088 ( 
.A(n_9670),
.Y(n_11088)
);

INVx2_ASAP7_75t_L g11089 ( 
.A(n_9670),
.Y(n_11089)
);

AND2x2_ASAP7_75t_L g11090 ( 
.A(n_10108),
.B(n_8952),
.Y(n_11090)
);

INVx1_ASAP7_75t_L g11091 ( 
.A(n_9596),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_9600),
.Y(n_11092)
);

AND2x2_ASAP7_75t_L g11093 ( 
.A(n_9758),
.B(n_8952),
.Y(n_11093)
);

AND2x2_ASAP7_75t_L g11094 ( 
.A(n_9879),
.B(n_8972),
.Y(n_11094)
);

NAND2x1p5_ASAP7_75t_L g11095 ( 
.A(n_9759),
.B(n_8780),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_9600),
.Y(n_11096)
);

OAI21x1_ASAP7_75t_L g11097 ( 
.A1(n_10143),
.A2(n_8264),
.B(n_8258),
.Y(n_11097)
);

INVx2_ASAP7_75t_L g11098 ( 
.A(n_9670),
.Y(n_11098)
);

AND2x2_ASAP7_75t_L g11099 ( 
.A(n_9879),
.B(n_8972),
.Y(n_11099)
);

INVx2_ASAP7_75t_L g11100 ( 
.A(n_9722),
.Y(n_11100)
);

AND2x2_ASAP7_75t_L g11101 ( 
.A(n_10704),
.B(n_8972),
.Y(n_11101)
);

INVx1_ASAP7_75t_L g11102 ( 
.A(n_9603),
.Y(n_11102)
);

INVx2_ASAP7_75t_SL g11103 ( 
.A(n_10080),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_9603),
.Y(n_11104)
);

INVx1_ASAP7_75t_L g11105 ( 
.A(n_9609),
.Y(n_11105)
);

INVx1_ASAP7_75t_L g11106 ( 
.A(n_9609),
.Y(n_11106)
);

INVx1_ASAP7_75t_L g11107 ( 
.A(n_9610),
.Y(n_11107)
);

INVx1_ASAP7_75t_L g11108 ( 
.A(n_9610),
.Y(n_11108)
);

INVx2_ASAP7_75t_L g11109 ( 
.A(n_9722),
.Y(n_11109)
);

INVx1_ASAP7_75t_L g11110 ( 
.A(n_9611),
.Y(n_11110)
);

INVx1_ASAP7_75t_L g11111 ( 
.A(n_9611),
.Y(n_11111)
);

INVx2_ASAP7_75t_L g11112 ( 
.A(n_9722),
.Y(n_11112)
);

INVx1_ASAP7_75t_SL g11113 ( 
.A(n_10274),
.Y(n_11113)
);

INVx2_ASAP7_75t_L g11114 ( 
.A(n_9722),
.Y(n_11114)
);

INVxp67_ASAP7_75t_SL g11115 ( 
.A(n_9625),
.Y(n_11115)
);

INVx2_ASAP7_75t_L g11116 ( 
.A(n_9766),
.Y(n_11116)
);

INVx1_ASAP7_75t_L g11117 ( 
.A(n_9612),
.Y(n_11117)
);

INVx2_ASAP7_75t_L g11118 ( 
.A(n_9766),
.Y(n_11118)
);

INVx1_ASAP7_75t_L g11119 ( 
.A(n_9612),
.Y(n_11119)
);

OAI21xp5_ASAP7_75t_L g11120 ( 
.A1(n_9882),
.A2(n_8593),
.B(n_8569),
.Y(n_11120)
);

NAND2xp5_ASAP7_75t_L g11121 ( 
.A(n_9688),
.B(n_9082),
.Y(n_11121)
);

INVx1_ASAP7_75t_L g11122 ( 
.A(n_9614),
.Y(n_11122)
);

OAI21xp5_ASAP7_75t_L g11123 ( 
.A1(n_10246),
.A2(n_9171),
.B(n_8591),
.Y(n_11123)
);

AO21x2_ASAP7_75t_L g11124 ( 
.A1(n_9654),
.A2(n_8908),
.B(n_9407),
.Y(n_11124)
);

INVx2_ASAP7_75t_L g11125 ( 
.A(n_9766),
.Y(n_11125)
);

INVx1_ASAP7_75t_L g11126 ( 
.A(n_9614),
.Y(n_11126)
);

BUFx2_ASAP7_75t_L g11127 ( 
.A(n_9799),
.Y(n_11127)
);

INVx1_ASAP7_75t_L g11128 ( 
.A(n_9619),
.Y(n_11128)
);

OR2x2_ASAP7_75t_L g11129 ( 
.A(n_9778),
.B(n_8417),
.Y(n_11129)
);

BUFx3_ASAP7_75t_L g11130 ( 
.A(n_9947),
.Y(n_11130)
);

INVx2_ASAP7_75t_L g11131 ( 
.A(n_9766),
.Y(n_11131)
);

BUFx2_ASAP7_75t_SL g11132 ( 
.A(n_10242),
.Y(n_11132)
);

INVx2_ASAP7_75t_L g11133 ( 
.A(n_9806),
.Y(n_11133)
);

INVx1_ASAP7_75t_L g11134 ( 
.A(n_9619),
.Y(n_11134)
);

AND2x2_ASAP7_75t_L g11135 ( 
.A(n_10704),
.B(n_8979),
.Y(n_11135)
);

INVx1_ASAP7_75t_L g11136 ( 
.A(n_9622),
.Y(n_11136)
);

AND2x2_ASAP7_75t_L g11137 ( 
.A(n_9702),
.B(n_8979),
.Y(n_11137)
);

NAND2xp5_ASAP7_75t_L g11138 ( 
.A(n_9807),
.B(n_9082),
.Y(n_11138)
);

OAI21x1_ASAP7_75t_L g11139 ( 
.A1(n_10053),
.A2(n_8264),
.B(n_8258),
.Y(n_11139)
);

INVxp33_ASAP7_75t_L g11140 ( 
.A(n_9708),
.Y(n_11140)
);

INVx1_ASAP7_75t_L g11141 ( 
.A(n_9622),
.Y(n_11141)
);

INVx1_ASAP7_75t_L g11142 ( 
.A(n_9623),
.Y(n_11142)
);

BUFx3_ASAP7_75t_L g11143 ( 
.A(n_9947),
.Y(n_11143)
);

INVx2_ASAP7_75t_L g11144 ( 
.A(n_9806),
.Y(n_11144)
);

INVx1_ASAP7_75t_L g11145 ( 
.A(n_9623),
.Y(n_11145)
);

AO21x2_ASAP7_75t_L g11146 ( 
.A1(n_9855),
.A2(n_9195),
.B(n_9017),
.Y(n_11146)
);

AOI21xp33_ASAP7_75t_L g11147 ( 
.A1(n_10164),
.A2(n_9235),
.B(n_8226),
.Y(n_11147)
);

OR2x2_ASAP7_75t_L g11148 ( 
.A(n_9778),
.B(n_8417),
.Y(n_11148)
);

INVx1_ASAP7_75t_L g11149 ( 
.A(n_9624),
.Y(n_11149)
);

INVx2_ASAP7_75t_SL g11150 ( 
.A(n_10080),
.Y(n_11150)
);

OAI21x1_ASAP7_75t_L g11151 ( 
.A1(n_10053),
.A2(n_9093),
.B(n_8387),
.Y(n_11151)
);

BUFx6f_ASAP7_75t_L g11152 ( 
.A(n_9665),
.Y(n_11152)
);

INVx1_ASAP7_75t_L g11153 ( 
.A(n_9624),
.Y(n_11153)
);

BUFx3_ASAP7_75t_L g11154 ( 
.A(n_10051),
.Y(n_11154)
);

HB1xp67_ASAP7_75t_L g11155 ( 
.A(n_9806),
.Y(n_11155)
);

BUFx3_ASAP7_75t_L g11156 ( 
.A(n_10051),
.Y(n_11156)
);

INVx1_ASAP7_75t_L g11157 ( 
.A(n_9628),
.Y(n_11157)
);

INVx2_ASAP7_75t_L g11158 ( 
.A(n_9806),
.Y(n_11158)
);

AND2x2_ASAP7_75t_L g11159 ( 
.A(n_9702),
.B(n_9998),
.Y(n_11159)
);

NAND2xp5_ASAP7_75t_L g11160 ( 
.A(n_9807),
.B(n_9118),
.Y(n_11160)
);

INVxp33_ASAP7_75t_L g11161 ( 
.A(n_9708),
.Y(n_11161)
);

INVx2_ASAP7_75t_L g11162 ( 
.A(n_9835),
.Y(n_11162)
);

INVx2_ASAP7_75t_L g11163 ( 
.A(n_9835),
.Y(n_11163)
);

BUFx3_ASAP7_75t_L g11164 ( 
.A(n_10051),
.Y(n_11164)
);

INVx2_ASAP7_75t_L g11165 ( 
.A(n_9835),
.Y(n_11165)
);

BUFx6f_ASAP7_75t_L g11166 ( 
.A(n_9665),
.Y(n_11166)
);

INVx2_ASAP7_75t_L g11167 ( 
.A(n_9835),
.Y(n_11167)
);

CKINVDCx5p33_ASAP7_75t_R g11168 ( 
.A(n_10522),
.Y(n_11168)
);

INVx1_ASAP7_75t_L g11169 ( 
.A(n_9628),
.Y(n_11169)
);

INVx1_ASAP7_75t_L g11170 ( 
.A(n_9633),
.Y(n_11170)
);

INVx1_ASAP7_75t_L g11171 ( 
.A(n_9633),
.Y(n_11171)
);

INVx2_ASAP7_75t_L g11172 ( 
.A(n_9839),
.Y(n_11172)
);

OR2x2_ASAP7_75t_L g11173 ( 
.A(n_9815),
.B(n_8430),
.Y(n_11173)
);

INVx1_ASAP7_75t_L g11174 ( 
.A(n_9636),
.Y(n_11174)
);

BUFx3_ASAP7_75t_L g11175 ( 
.A(n_10082),
.Y(n_11175)
);

AND2x2_ASAP7_75t_L g11176 ( 
.A(n_9702),
.B(n_8979),
.Y(n_11176)
);

INVx1_ASAP7_75t_L g11177 ( 
.A(n_9636),
.Y(n_11177)
);

INVx2_ASAP7_75t_L g11178 ( 
.A(n_9839),
.Y(n_11178)
);

NAND2xp5_ASAP7_75t_L g11179 ( 
.A(n_9718),
.B(n_9118),
.Y(n_11179)
);

BUFx3_ASAP7_75t_L g11180 ( 
.A(n_10082),
.Y(n_11180)
);

AOI21x1_ASAP7_75t_L g11181 ( 
.A1(n_9650),
.A2(n_8992),
.B(n_8978),
.Y(n_11181)
);

NOR2x1_ASAP7_75t_R g11182 ( 
.A(n_9823),
.B(n_7312),
.Y(n_11182)
);

NAND2xp5_ASAP7_75t_L g11183 ( 
.A(n_9718),
.B(n_9008),
.Y(n_11183)
);

INVx1_ASAP7_75t_L g11184 ( 
.A(n_9640),
.Y(n_11184)
);

INVx1_ASAP7_75t_L g11185 ( 
.A(n_9640),
.Y(n_11185)
);

OAI21xp5_ASAP7_75t_L g11186 ( 
.A1(n_10246),
.A2(n_8591),
.B(n_8437),
.Y(n_11186)
);

HB1xp67_ASAP7_75t_L g11187 ( 
.A(n_9839),
.Y(n_11187)
);

INVx1_ASAP7_75t_L g11188 ( 
.A(n_9647),
.Y(n_11188)
);

HB1xp67_ASAP7_75t_L g11189 ( 
.A(n_9839),
.Y(n_11189)
);

INVx2_ASAP7_75t_SL g11190 ( 
.A(n_10671),
.Y(n_11190)
);

INVx1_ASAP7_75t_L g11191 ( 
.A(n_9647),
.Y(n_11191)
);

INVx2_ASAP7_75t_L g11192 ( 
.A(n_9843),
.Y(n_11192)
);

INVx1_ASAP7_75t_L g11193 ( 
.A(n_9661),
.Y(n_11193)
);

BUFx6f_ASAP7_75t_L g11194 ( 
.A(n_9823),
.Y(n_11194)
);

BUFx3_ASAP7_75t_L g11195 ( 
.A(n_10082),
.Y(n_11195)
);

INVx3_ASAP7_75t_L g11196 ( 
.A(n_9769),
.Y(n_11196)
);

INVx2_ASAP7_75t_L g11197 ( 
.A(n_9843),
.Y(n_11197)
);

BUFx6f_ASAP7_75t_L g11198 ( 
.A(n_9823),
.Y(n_11198)
);

NAND2xp5_ASAP7_75t_L g11199 ( 
.A(n_10270),
.B(n_9030),
.Y(n_11199)
);

INVx1_ASAP7_75t_SL g11200 ( 
.A(n_10342),
.Y(n_11200)
);

AND2x4_ASAP7_75t_L g11201 ( 
.A(n_9769),
.B(n_8259),
.Y(n_11201)
);

OAI21xp5_ASAP7_75t_L g11202 ( 
.A1(n_10292),
.A2(n_9287),
.B(n_8909),
.Y(n_11202)
);

AOI22xp33_ASAP7_75t_L g11203 ( 
.A1(n_10557),
.A2(n_9135),
.B1(n_9131),
.B2(n_8986),
.Y(n_11203)
);

AO21x1_ASAP7_75t_SL g11204 ( 
.A1(n_11003),
.A2(n_9368),
.B(n_9363),
.Y(n_11204)
);

INVx2_ASAP7_75t_L g11205 ( 
.A(n_9843),
.Y(n_11205)
);

INVx2_ASAP7_75t_L g11206 ( 
.A(n_9843),
.Y(n_11206)
);

INVx1_ASAP7_75t_L g11207 ( 
.A(n_9661),
.Y(n_11207)
);

INVx2_ASAP7_75t_L g11208 ( 
.A(n_9857),
.Y(n_11208)
);

INVx1_ASAP7_75t_L g11209 ( 
.A(n_9662),
.Y(n_11209)
);

INVx1_ASAP7_75t_L g11210 ( 
.A(n_9662),
.Y(n_11210)
);

INVx2_ASAP7_75t_L g11211 ( 
.A(n_9857),
.Y(n_11211)
);

INVx2_ASAP7_75t_L g11212 ( 
.A(n_9857),
.Y(n_11212)
);

INVx1_ASAP7_75t_L g11213 ( 
.A(n_9666),
.Y(n_11213)
);

OAI21x1_ASAP7_75t_L g11214 ( 
.A1(n_9826),
.A2(n_9093),
.B(n_8387),
.Y(n_11214)
);

INVx2_ASAP7_75t_L g11215 ( 
.A(n_9857),
.Y(n_11215)
);

BUFx3_ASAP7_75t_L g11216 ( 
.A(n_9799),
.Y(n_11216)
);

NAND3xp33_ASAP7_75t_L g11217 ( 
.A(n_10252),
.B(n_8745),
.C(n_8278),
.Y(n_11217)
);

INVx2_ASAP7_75t_L g11218 ( 
.A(n_9805),
.Y(n_11218)
);

AND2x2_ASAP7_75t_L g11219 ( 
.A(n_9998),
.B(n_9088),
.Y(n_11219)
);

INVx1_ASAP7_75t_L g11220 ( 
.A(n_9666),
.Y(n_11220)
);

INVx2_ASAP7_75t_L g11221 ( 
.A(n_9805),
.Y(n_11221)
);

BUFx6f_ASAP7_75t_L g11222 ( 
.A(n_9708),
.Y(n_11222)
);

INVx1_ASAP7_75t_L g11223 ( 
.A(n_9667),
.Y(n_11223)
);

INVx1_ASAP7_75t_L g11224 ( 
.A(n_9667),
.Y(n_11224)
);

INVx2_ASAP7_75t_L g11225 ( 
.A(n_9805),
.Y(n_11225)
);

NAND2xp5_ASAP7_75t_L g11226 ( 
.A(n_10270),
.B(n_10277),
.Y(n_11226)
);

OAI21xp5_ASAP7_75t_L g11227 ( 
.A1(n_10292),
.A2(n_9287),
.B(n_8278),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_9673),
.Y(n_11228)
);

INVx1_ASAP7_75t_L g11229 ( 
.A(n_9673),
.Y(n_11229)
);

INVx1_ASAP7_75t_L g11230 ( 
.A(n_9682),
.Y(n_11230)
);

HB1xp67_ASAP7_75t_L g11231 ( 
.A(n_10974),
.Y(n_11231)
);

INVx1_ASAP7_75t_L g11232 ( 
.A(n_9682),
.Y(n_11232)
);

AND2x2_ASAP7_75t_L g11233 ( 
.A(n_10527),
.B(n_9088),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_9684),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_9684),
.Y(n_11235)
);

INVx1_ASAP7_75t_SL g11236 ( 
.A(n_10342),
.Y(n_11236)
);

INVx3_ASAP7_75t_L g11237 ( 
.A(n_9769),
.Y(n_11237)
);

OAI221xp5_ASAP7_75t_L g11238 ( 
.A1(n_10089),
.A2(n_9039),
.B1(n_9139),
.B2(n_9100),
.C(n_9069),
.Y(n_11238)
);

INVx1_ASAP7_75t_L g11239 ( 
.A(n_9686),
.Y(n_11239)
);

INVx1_ASAP7_75t_L g11240 ( 
.A(n_9686),
.Y(n_11240)
);

OAI21x1_ASAP7_75t_L g11241 ( 
.A1(n_9826),
.A2(n_8387),
.B(n_8828),
.Y(n_11241)
);

INVx1_ASAP7_75t_L g11242 ( 
.A(n_9698),
.Y(n_11242)
);

INVxp33_ASAP7_75t_L g11243 ( 
.A(n_9708),
.Y(n_11243)
);

HB1xp67_ASAP7_75t_L g11244 ( 
.A(n_10974),
.Y(n_11244)
);

AO21x1_ASAP7_75t_L g11245 ( 
.A1(n_9632),
.A2(n_8406),
.B(n_8594),
.Y(n_11245)
);

INVx1_ASAP7_75t_L g11246 ( 
.A(n_9698),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_9707),
.Y(n_11247)
);

INVx2_ASAP7_75t_L g11248 ( 
.A(n_9805),
.Y(n_11248)
);

OR2x6_ASAP7_75t_L g11249 ( 
.A(n_9626),
.B(n_8780),
.Y(n_11249)
);

INVx1_ASAP7_75t_L g11250 ( 
.A(n_9707),
.Y(n_11250)
);

CKINVDCx20_ASAP7_75t_R g11251 ( 
.A(n_9621),
.Y(n_11251)
);

INVx2_ASAP7_75t_L g11252 ( 
.A(n_10123),
.Y(n_11252)
);

AND2x4_ASAP7_75t_L g11253 ( 
.A(n_9769),
.B(n_8259),
.Y(n_11253)
);

AOI22xp33_ASAP7_75t_L g11254 ( 
.A1(n_10642),
.A2(n_9135),
.B1(n_9131),
.B2(n_8986),
.Y(n_11254)
);

INVx1_ASAP7_75t_SL g11255 ( 
.A(n_10376),
.Y(n_11255)
);

OAI22xp33_ASAP7_75t_L g11256 ( 
.A1(n_10485),
.A2(n_9432),
.B1(n_8745),
.B2(n_8476),
.Y(n_11256)
);

INVx1_ASAP7_75t_L g11257 ( 
.A(n_9711),
.Y(n_11257)
);

OAI21x1_ASAP7_75t_L g11258 ( 
.A1(n_10495),
.A2(n_8892),
.B(n_8828),
.Y(n_11258)
);

INVx1_ASAP7_75t_L g11259 ( 
.A(n_9711),
.Y(n_11259)
);

INVx1_ASAP7_75t_L g11260 ( 
.A(n_9714),
.Y(n_11260)
);

INVx1_ASAP7_75t_L g11261 ( 
.A(n_9714),
.Y(n_11261)
);

OAI21x1_ASAP7_75t_L g11262 ( 
.A1(n_10495),
.A2(n_8892),
.B(n_8828),
.Y(n_11262)
);

INVx2_ASAP7_75t_L g11263 ( 
.A(n_10123),
.Y(n_11263)
);

INVx1_ASAP7_75t_L g11264 ( 
.A(n_9723),
.Y(n_11264)
);

INVx2_ASAP7_75t_L g11265 ( 
.A(n_10123),
.Y(n_11265)
);

OAI21x1_ASAP7_75t_L g11266 ( 
.A1(n_10495),
.A2(n_8892),
.B(n_9062),
.Y(n_11266)
);

INVx1_ASAP7_75t_L g11267 ( 
.A(n_9723),
.Y(n_11267)
);

INVx2_ASAP7_75t_L g11268 ( 
.A(n_10123),
.Y(n_11268)
);

OAI21xp5_ASAP7_75t_L g11269 ( 
.A1(n_10477),
.A2(n_9117),
.B(n_8760),
.Y(n_11269)
);

INVx1_ASAP7_75t_L g11270 ( 
.A(n_9728),
.Y(n_11270)
);

INVx2_ASAP7_75t_L g11271 ( 
.A(n_10169),
.Y(n_11271)
);

INVx1_ASAP7_75t_L g11272 ( 
.A(n_9728),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_9738),
.Y(n_11273)
);

BUFx2_ASAP7_75t_SL g11274 ( 
.A(n_10328),
.Y(n_11274)
);

INVx1_ASAP7_75t_L g11275 ( 
.A(n_9738),
.Y(n_11275)
);

OAI21x1_ASAP7_75t_L g11276 ( 
.A1(n_9650),
.A2(n_8281),
.B(n_8460),
.Y(n_11276)
);

INVx2_ASAP7_75t_L g11277 ( 
.A(n_10169),
.Y(n_11277)
);

INVx1_ASAP7_75t_L g11278 ( 
.A(n_9739),
.Y(n_11278)
);

AND2x2_ASAP7_75t_L g11279 ( 
.A(n_10527),
.B(n_9088),
.Y(n_11279)
);

INVx1_ASAP7_75t_L g11280 ( 
.A(n_9739),
.Y(n_11280)
);

AOI21x1_ASAP7_75t_L g11281 ( 
.A1(n_9589),
.A2(n_8992),
.B(n_8978),
.Y(n_11281)
);

INVx1_ASAP7_75t_L g11282 ( 
.A(n_9740),
.Y(n_11282)
);

AND2x4_ASAP7_75t_SL g11283 ( 
.A(n_10822),
.B(n_8780),
.Y(n_11283)
);

HB1xp67_ASAP7_75t_L g11284 ( 
.A(n_10994),
.Y(n_11284)
);

INVx1_ASAP7_75t_L g11285 ( 
.A(n_9740),
.Y(n_11285)
);

INVx2_ASAP7_75t_L g11286 ( 
.A(n_10169),
.Y(n_11286)
);

AOI21x1_ASAP7_75t_L g11287 ( 
.A1(n_9589),
.A2(n_9606),
.B(n_10410),
.Y(n_11287)
);

INVx1_ASAP7_75t_SL g11288 ( 
.A(n_10376),
.Y(n_11288)
);

AO21x2_ASAP7_75t_L g11289 ( 
.A1(n_10329),
.A2(n_10040),
.B(n_9899),
.Y(n_11289)
);

INVx2_ASAP7_75t_L g11290 ( 
.A(n_10169),
.Y(n_11290)
);

INVx1_ASAP7_75t_L g11291 ( 
.A(n_9741),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_9741),
.Y(n_11292)
);

INVx1_ASAP7_75t_L g11293 ( 
.A(n_9745),
.Y(n_11293)
);

INVx2_ASAP7_75t_L g11294 ( 
.A(n_10186),
.Y(n_11294)
);

INVx2_ASAP7_75t_SL g11295 ( 
.A(n_10671),
.Y(n_11295)
);

OA21x2_ASAP7_75t_L g11296 ( 
.A1(n_9784),
.A2(n_8282),
.B(n_8281),
.Y(n_11296)
);

NAND2xp5_ASAP7_75t_L g11297 ( 
.A(n_10277),
.B(n_9039),
.Y(n_11297)
);

INVx3_ASAP7_75t_L g11298 ( 
.A(n_10125),
.Y(n_11298)
);

INVx2_ASAP7_75t_L g11299 ( 
.A(n_10186),
.Y(n_11299)
);

INVx2_ASAP7_75t_L g11300 ( 
.A(n_10186),
.Y(n_11300)
);

INVx2_ASAP7_75t_L g11301 ( 
.A(n_10186),
.Y(n_11301)
);

INVx2_ASAP7_75t_L g11302 ( 
.A(n_10189),
.Y(n_11302)
);

INVx1_ASAP7_75t_L g11303 ( 
.A(n_9745),
.Y(n_11303)
);

INVx1_ASAP7_75t_L g11304 ( 
.A(n_9749),
.Y(n_11304)
);

AO21x1_ASAP7_75t_L g11305 ( 
.A1(n_9658),
.A2(n_8406),
.B(n_8594),
.Y(n_11305)
);

BUFx3_ASAP7_75t_L g11306 ( 
.A(n_9799),
.Y(n_11306)
);

INVx2_ASAP7_75t_L g11307 ( 
.A(n_10189),
.Y(n_11307)
);

INVx2_ASAP7_75t_L g11308 ( 
.A(n_10189),
.Y(n_11308)
);

INVx1_ASAP7_75t_L g11309 ( 
.A(n_9749),
.Y(n_11309)
);

INVx2_ASAP7_75t_L g11310 ( 
.A(n_10189),
.Y(n_11310)
);

INVx2_ASAP7_75t_L g11311 ( 
.A(n_10198),
.Y(n_11311)
);

INVx1_ASAP7_75t_L g11312 ( 
.A(n_9750),
.Y(n_11312)
);

INVx1_ASAP7_75t_L g11313 ( 
.A(n_9750),
.Y(n_11313)
);

INVx1_ASAP7_75t_SL g11314 ( 
.A(n_10388),
.Y(n_11314)
);

INVx2_ASAP7_75t_L g11315 ( 
.A(n_10198),
.Y(n_11315)
);

INVx2_ASAP7_75t_L g11316 ( 
.A(n_10198),
.Y(n_11316)
);

INVx3_ASAP7_75t_L g11317 ( 
.A(n_10125),
.Y(n_11317)
);

INVx2_ASAP7_75t_L g11318 ( 
.A(n_10198),
.Y(n_11318)
);

INVx1_ASAP7_75t_L g11319 ( 
.A(n_9752),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_9752),
.Y(n_11320)
);

INVx2_ASAP7_75t_L g11321 ( 
.A(n_10205),
.Y(n_11321)
);

INVx2_ASAP7_75t_L g11322 ( 
.A(n_10205),
.Y(n_11322)
);

AOI22xp33_ASAP7_75t_L g11323 ( 
.A1(n_10642),
.A2(n_10698),
.B1(n_10706),
.B2(n_10663),
.Y(n_11323)
);

AND2x4_ASAP7_75t_L g11324 ( 
.A(n_10399),
.B(n_8259),
.Y(n_11324)
);

CKINVDCx6p67_ASAP7_75t_R g11325 ( 
.A(n_10059),
.Y(n_11325)
);

NAND2xp5_ASAP7_75t_L g11326 ( 
.A(n_10353),
.B(n_9069),
.Y(n_11326)
);

INVx1_ASAP7_75t_L g11327 ( 
.A(n_9753),
.Y(n_11327)
);

INVx2_ASAP7_75t_L g11328 ( 
.A(n_10205),
.Y(n_11328)
);

AOI22xp5_ASAP7_75t_L g11329 ( 
.A1(n_10663),
.A2(n_8548),
.B1(n_8616),
.B2(n_9550),
.Y(n_11329)
);

INVx1_ASAP7_75t_L g11330 ( 
.A(n_9753),
.Y(n_11330)
);

HB1xp67_ASAP7_75t_SL g11331 ( 
.A(n_9735),
.Y(n_11331)
);

OAI22xp5_ASAP7_75t_L g11332 ( 
.A1(n_10485),
.A2(n_8548),
.B1(n_8616),
.B2(n_9166),
.Y(n_11332)
);

CKINVDCx5p33_ASAP7_75t_R g11333 ( 
.A(n_10523),
.Y(n_11333)
);

OAI21x1_ASAP7_75t_L g11334 ( 
.A1(n_9606),
.A2(n_8281),
.B(n_8460),
.Y(n_11334)
);

AND2x2_ASAP7_75t_L g11335 ( 
.A(n_10590),
.B(n_9097),
.Y(n_11335)
);

INVx1_ASAP7_75t_L g11336 ( 
.A(n_9754),
.Y(n_11336)
);

INVx2_ASAP7_75t_L g11337 ( 
.A(n_10205),
.Y(n_11337)
);

INVx2_ASAP7_75t_L g11338 ( 
.A(n_10251),
.Y(n_11338)
);

HB1xp67_ASAP7_75t_L g11339 ( 
.A(n_10994),
.Y(n_11339)
);

INVx1_ASAP7_75t_L g11340 ( 
.A(n_9754),
.Y(n_11340)
);

INVx2_ASAP7_75t_L g11341 ( 
.A(n_10251),
.Y(n_11341)
);

AND2x2_ASAP7_75t_L g11342 ( 
.A(n_10590),
.B(n_9097),
.Y(n_11342)
);

AO21x2_ASAP7_75t_L g11343 ( 
.A1(n_10329),
.A2(n_9195),
.B(n_8760),
.Y(n_11343)
);

INVx2_ASAP7_75t_L g11344 ( 
.A(n_10251),
.Y(n_11344)
);

INVx2_ASAP7_75t_L g11345 ( 
.A(n_10251),
.Y(n_11345)
);

NOR2xp33_ASAP7_75t_L g11346 ( 
.A(n_10347),
.B(n_9556),
.Y(n_11346)
);

INVx2_ASAP7_75t_L g11347 ( 
.A(n_10259),
.Y(n_11347)
);

INVx1_ASAP7_75t_L g11348 ( 
.A(n_9756),
.Y(n_11348)
);

INVx1_ASAP7_75t_L g11349 ( 
.A(n_9756),
.Y(n_11349)
);

OA21x2_ASAP7_75t_L g11350 ( 
.A1(n_9784),
.A2(n_9789),
.B(n_9788),
.Y(n_11350)
);

INVx1_ASAP7_75t_L g11351 ( 
.A(n_9762),
.Y(n_11351)
);

INVx1_ASAP7_75t_L g11352 ( 
.A(n_9762),
.Y(n_11352)
);

INVx2_ASAP7_75t_L g11353 ( 
.A(n_10259),
.Y(n_11353)
);

NAND2xp5_ASAP7_75t_L g11354 ( 
.A(n_10353),
.B(n_9100),
.Y(n_11354)
);

INVx8_ASAP7_75t_L g11355 ( 
.A(n_10093),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_9763),
.Y(n_11356)
);

AND2x2_ASAP7_75t_L g11357 ( 
.A(n_9834),
.B(n_9097),
.Y(n_11357)
);

INVx1_ASAP7_75t_L g11358 ( 
.A(n_9763),
.Y(n_11358)
);

INVx1_ASAP7_75t_L g11359 ( 
.A(n_9772),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_9772),
.Y(n_11360)
);

BUFx2_ASAP7_75t_L g11361 ( 
.A(n_10301),
.Y(n_11361)
);

OAI21x1_ASAP7_75t_L g11362 ( 
.A1(n_10173),
.A2(n_8495),
.B(n_8460),
.Y(n_11362)
);

INVx2_ASAP7_75t_SL g11363 ( 
.A(n_10671),
.Y(n_11363)
);

OAI21x1_ASAP7_75t_L g11364 ( 
.A1(n_10173),
.A2(n_8495),
.B(n_8397),
.Y(n_11364)
);

INVx1_ASAP7_75t_L g11365 ( 
.A(n_9773),
.Y(n_11365)
);

HB1xp67_ASAP7_75t_L g11366 ( 
.A(n_11018),
.Y(n_11366)
);

INVx1_ASAP7_75t_L g11367 ( 
.A(n_9773),
.Y(n_11367)
);

AND2x2_ASAP7_75t_L g11368 ( 
.A(n_9834),
.B(n_9198),
.Y(n_11368)
);

INVx2_ASAP7_75t_L g11369 ( 
.A(n_10259),
.Y(n_11369)
);

INVx2_ASAP7_75t_L g11370 ( 
.A(n_10259),
.Y(n_11370)
);

AOI222xp33_ASAP7_75t_L g11371 ( 
.A1(n_10698),
.A2(n_8860),
.B1(n_9563),
.B2(n_9139),
.C1(n_9505),
.C2(n_9491),
.Y(n_11371)
);

INVx1_ASAP7_75t_L g11372 ( 
.A(n_9780),
.Y(n_11372)
);

INVx1_ASAP7_75t_L g11373 ( 
.A(n_9780),
.Y(n_11373)
);

BUFx3_ASAP7_75t_L g11374 ( 
.A(n_10680),
.Y(n_11374)
);

INVx3_ASAP7_75t_L g11375 ( 
.A(n_10125),
.Y(n_11375)
);

NAND2xp5_ASAP7_75t_L g11376 ( 
.A(n_10366),
.B(n_9117),
.Y(n_11376)
);

HB1xp67_ASAP7_75t_L g11377 ( 
.A(n_11018),
.Y(n_11377)
);

INVx1_ASAP7_75t_L g11378 ( 
.A(n_9787),
.Y(n_11378)
);

AOI22xp33_ASAP7_75t_L g11379 ( 
.A1(n_10706),
.A2(n_9135),
.B1(n_9131),
.B2(n_8986),
.Y(n_11379)
);

NOR2x1_ASAP7_75t_R g11380 ( 
.A(n_9696),
.B(n_7326),
.Y(n_11380)
);

AOI21xp5_ASAP7_75t_L g11381 ( 
.A1(n_10164),
.A2(n_8173),
.B(n_8556),
.Y(n_11381)
);

INVx1_ASAP7_75t_L g11382 ( 
.A(n_9787),
.Y(n_11382)
);

INVx1_ASAP7_75t_L g11383 ( 
.A(n_9790),
.Y(n_11383)
);

BUFx2_ASAP7_75t_SL g11384 ( 
.A(n_10372),
.Y(n_11384)
);

INVx2_ASAP7_75t_L g11385 ( 
.A(n_10267),
.Y(n_11385)
);

INVx3_ASAP7_75t_L g11386 ( 
.A(n_10125),
.Y(n_11386)
);

INVx1_ASAP7_75t_L g11387 ( 
.A(n_9790),
.Y(n_11387)
);

INVx2_ASAP7_75t_L g11388 ( 
.A(n_10267),
.Y(n_11388)
);

NAND2xp5_ASAP7_75t_SL g11389 ( 
.A(n_10665),
.B(n_9566),
.Y(n_11389)
);

INVx1_ASAP7_75t_L g11390 ( 
.A(n_9791),
.Y(n_11390)
);

OAI21x1_ASAP7_75t_L g11391 ( 
.A1(n_10217),
.A2(n_8495),
.B(n_8397),
.Y(n_11391)
);

INVx1_ASAP7_75t_L g11392 ( 
.A(n_9791),
.Y(n_11392)
);

INVx2_ASAP7_75t_L g11393 ( 
.A(n_10267),
.Y(n_11393)
);

AOI22xp33_ASAP7_75t_SL g11394 ( 
.A1(n_10838),
.A2(n_8297),
.B1(n_8640),
.B2(n_8621),
.Y(n_11394)
);

HB1xp67_ASAP7_75t_SL g11395 ( 
.A(n_9735),
.Y(n_11395)
);

OAI21x1_ASAP7_75t_L g11396 ( 
.A1(n_10217),
.A2(n_8397),
.B(n_9246),
.Y(n_11396)
);

INVx1_ASAP7_75t_L g11397 ( 
.A(n_9793),
.Y(n_11397)
);

INVx2_ASAP7_75t_L g11398 ( 
.A(n_10267),
.Y(n_11398)
);

INVx2_ASAP7_75t_SL g11399 ( 
.A(n_10671),
.Y(n_11399)
);

INVx2_ASAP7_75t_L g11400 ( 
.A(n_10271),
.Y(n_11400)
);

BUFx3_ASAP7_75t_L g11401 ( 
.A(n_10680),
.Y(n_11401)
);

AO21x1_ASAP7_75t_L g11402 ( 
.A1(n_10801),
.A2(n_8826),
.B(n_8740),
.Y(n_11402)
);

INVx1_ASAP7_75t_L g11403 ( 
.A(n_9793),
.Y(n_11403)
);

INVx2_ASAP7_75t_L g11404 ( 
.A(n_10271),
.Y(n_11404)
);

OA21x2_ASAP7_75t_L g11405 ( 
.A1(n_9784),
.A2(n_9789),
.B(n_9788),
.Y(n_11405)
);

HB1xp67_ASAP7_75t_L g11406 ( 
.A(n_9607),
.Y(n_11406)
);

HB1xp67_ASAP7_75t_L g11407 ( 
.A(n_9915),
.Y(n_11407)
);

AND2x2_ASAP7_75t_L g11408 ( 
.A(n_10650),
.B(n_9198),
.Y(n_11408)
);

AND2x4_ASAP7_75t_L g11409 ( 
.A(n_10399),
.B(n_8259),
.Y(n_11409)
);

BUFx3_ASAP7_75t_L g11410 ( 
.A(n_10680),
.Y(n_11410)
);

INVx1_ASAP7_75t_L g11411 ( 
.A(n_9796),
.Y(n_11411)
);

HB1xp67_ASAP7_75t_L g11412 ( 
.A(n_9950),
.Y(n_11412)
);

INVx2_ASAP7_75t_L g11413 ( 
.A(n_10271),
.Y(n_11413)
);

INVx1_ASAP7_75t_L g11414 ( 
.A(n_9796),
.Y(n_11414)
);

INVx2_ASAP7_75t_L g11415 ( 
.A(n_10271),
.Y(n_11415)
);

OR2x2_ASAP7_75t_L g11416 ( 
.A(n_9815),
.B(n_8430),
.Y(n_11416)
);

OA21x2_ASAP7_75t_L g11417 ( 
.A1(n_9788),
.A2(n_8282),
.B(n_8155),
.Y(n_11417)
);

INVx1_ASAP7_75t_L g11418 ( 
.A(n_9801),
.Y(n_11418)
);

OA21x2_ASAP7_75t_L g11419 ( 
.A1(n_9789),
.A2(n_8155),
.B(n_8266),
.Y(n_11419)
);

INVx2_ASAP7_75t_L g11420 ( 
.A(n_10306),
.Y(n_11420)
);

INVx1_ASAP7_75t_L g11421 ( 
.A(n_9801),
.Y(n_11421)
);

INVx1_ASAP7_75t_L g11422 ( 
.A(n_9812),
.Y(n_11422)
);

INVx2_ASAP7_75t_L g11423 ( 
.A(n_10306),
.Y(n_11423)
);

INVx2_ASAP7_75t_L g11424 ( 
.A(n_10306),
.Y(n_11424)
);

BUFx6f_ASAP7_75t_L g11425 ( 
.A(n_9708),
.Y(n_11425)
);

INVx3_ASAP7_75t_L g11426 ( 
.A(n_9708),
.Y(n_11426)
);

AND2x4_ASAP7_75t_L g11427 ( 
.A(n_10399),
.B(n_8346),
.Y(n_11427)
);

HB1xp67_ASAP7_75t_L g11428 ( 
.A(n_9734),
.Y(n_11428)
);

INVx1_ASAP7_75t_L g11429 ( 
.A(n_9812),
.Y(n_11429)
);

INVx2_ASAP7_75t_L g11430 ( 
.A(n_10306),
.Y(n_11430)
);

INVx2_ASAP7_75t_L g11431 ( 
.A(n_10314),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_10314),
.Y(n_11432)
);

INVx1_ASAP7_75t_L g11433 ( 
.A(n_9816),
.Y(n_11433)
);

INVx2_ASAP7_75t_L g11434 ( 
.A(n_10314),
.Y(n_11434)
);

INVx1_ASAP7_75t_L g11435 ( 
.A(n_9816),
.Y(n_11435)
);

INVx1_ASAP7_75t_L g11436 ( 
.A(n_9819),
.Y(n_11436)
);

HB1xp67_ASAP7_75t_L g11437 ( 
.A(n_9802),
.Y(n_11437)
);

AND2x4_ASAP7_75t_SL g11438 ( 
.A(n_10822),
.B(n_8793),
.Y(n_11438)
);

INVx1_ASAP7_75t_SL g11439 ( 
.A(n_10388),
.Y(n_11439)
);

INVx1_ASAP7_75t_L g11440 ( 
.A(n_9819),
.Y(n_11440)
);

INVx1_ASAP7_75t_L g11441 ( 
.A(n_9825),
.Y(n_11441)
);

AND2x2_ASAP7_75t_L g11442 ( 
.A(n_10650),
.B(n_9198),
.Y(n_11442)
);

HB1xp67_ASAP7_75t_L g11443 ( 
.A(n_9824),
.Y(n_11443)
);

INVx2_ASAP7_75t_L g11444 ( 
.A(n_10314),
.Y(n_11444)
);

INVx1_ASAP7_75t_L g11445 ( 
.A(n_9825),
.Y(n_11445)
);

OAI21xp5_ASAP7_75t_L g11446 ( 
.A1(n_10477),
.A2(n_9006),
.B(n_8173),
.Y(n_11446)
);

OAI21x1_ASAP7_75t_L g11447 ( 
.A1(n_10516),
.A2(n_9246),
.B(n_8332),
.Y(n_11447)
);

INVx2_ASAP7_75t_L g11448 ( 
.A(n_10516),
.Y(n_11448)
);

INVx3_ASAP7_75t_L g11449 ( 
.A(n_9764),
.Y(n_11449)
);

OAI21x1_ASAP7_75t_L g11450 ( 
.A1(n_10516),
.A2(n_9246),
.B(n_8332),
.Y(n_11450)
);

INVx2_ASAP7_75t_L g11451 ( 
.A(n_10516),
.Y(n_11451)
);

BUFx3_ASAP7_75t_L g11452 ( 
.A(n_10093),
.Y(n_11452)
);

HB1xp67_ASAP7_75t_L g11453 ( 
.A(n_9831),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_9838),
.Y(n_11454)
);

INVx2_ASAP7_75t_L g11455 ( 
.A(n_10520),
.Y(n_11455)
);

AND2x4_ASAP7_75t_L g11456 ( 
.A(n_10399),
.B(n_8346),
.Y(n_11456)
);

AND2x2_ASAP7_75t_L g11457 ( 
.A(n_11020),
.B(n_9263),
.Y(n_11457)
);

AND2x2_ASAP7_75t_L g11458 ( 
.A(n_11020),
.B(n_9263),
.Y(n_11458)
);

OR2x6_ASAP7_75t_L g11459 ( 
.A(n_9626),
.B(n_8793),
.Y(n_11459)
);

BUFx3_ASAP7_75t_L g11460 ( 
.A(n_10093),
.Y(n_11460)
);

HB1xp67_ASAP7_75t_L g11461 ( 
.A(n_9893),
.Y(n_11461)
);

OAI21x1_ASAP7_75t_L g11462 ( 
.A1(n_10520),
.A2(n_8332),
.B(n_8323),
.Y(n_11462)
);

INVx1_ASAP7_75t_L g11463 ( 
.A(n_9838),
.Y(n_11463)
);

INVx2_ASAP7_75t_SL g11464 ( 
.A(n_9914),
.Y(n_11464)
);

INVx1_ASAP7_75t_L g11465 ( 
.A(n_9850),
.Y(n_11465)
);

INVx2_ASAP7_75t_L g11466 ( 
.A(n_10520),
.Y(n_11466)
);

OAI21x1_ASAP7_75t_L g11467 ( 
.A1(n_10520),
.A2(n_10609),
.B(n_10605),
.Y(n_11467)
);

HB1xp67_ASAP7_75t_L g11468 ( 
.A(n_9719),
.Y(n_11468)
);

INVx1_ASAP7_75t_L g11469 ( 
.A(n_9850),
.Y(n_11469)
);

INVx1_ASAP7_75t_L g11470 ( 
.A(n_9858),
.Y(n_11470)
);

AND2x2_ASAP7_75t_L g11471 ( 
.A(n_11020),
.B(n_9263),
.Y(n_11471)
);

AND2x2_ASAP7_75t_L g11472 ( 
.A(n_11020),
.B(n_9304),
.Y(n_11472)
);

INVx3_ASAP7_75t_L g11473 ( 
.A(n_9764),
.Y(n_11473)
);

INVx1_ASAP7_75t_L g11474 ( 
.A(n_9858),
.Y(n_11474)
);

INVx1_ASAP7_75t_L g11475 ( 
.A(n_9865),
.Y(n_11475)
);

AO21x1_ASAP7_75t_SL g11476 ( 
.A1(n_11003),
.A2(n_9363),
.B(n_9353),
.Y(n_11476)
);

AND2x2_ASAP7_75t_L g11477 ( 
.A(n_11020),
.B(n_9304),
.Y(n_11477)
);

INVx2_ASAP7_75t_L g11478 ( 
.A(n_10605),
.Y(n_11478)
);

INVx2_ASAP7_75t_L g11479 ( 
.A(n_10605),
.Y(n_11479)
);

OAI21xp5_ASAP7_75t_L g11480 ( 
.A1(n_10164),
.A2(n_9006),
.B(n_8280),
.Y(n_11480)
);

HB1xp67_ASAP7_75t_L g11481 ( 
.A(n_9719),
.Y(n_11481)
);

OAI21x1_ASAP7_75t_L g11482 ( 
.A1(n_10605),
.A2(n_8323),
.B(n_8850),
.Y(n_11482)
);

OR2x2_ASAP7_75t_L g11483 ( 
.A(n_9599),
.B(n_8434),
.Y(n_11483)
);

OR2x6_ASAP7_75t_L g11484 ( 
.A(n_9626),
.B(n_8793),
.Y(n_11484)
);

INVx1_ASAP7_75t_L g11485 ( 
.A(n_9865),
.Y(n_11485)
);

CKINVDCx14_ASAP7_75t_R g11486 ( 
.A(n_10718),
.Y(n_11486)
);

INVx1_ASAP7_75t_L g11487 ( 
.A(n_9868),
.Y(n_11487)
);

INVx1_ASAP7_75t_L g11488 ( 
.A(n_9868),
.Y(n_11488)
);

INVx2_ASAP7_75t_L g11489 ( 
.A(n_10609),
.Y(n_11489)
);

INVx2_ASAP7_75t_SL g11490 ( 
.A(n_9914),
.Y(n_11490)
);

AND2x4_ASAP7_75t_L g11491 ( 
.A(n_10399),
.B(n_10442),
.Y(n_11491)
);

INVx1_ASAP7_75t_L g11492 ( 
.A(n_9877),
.Y(n_11492)
);

INVxp67_ASAP7_75t_L g11493 ( 
.A(n_10487),
.Y(n_11493)
);

INVx2_ASAP7_75t_L g11494 ( 
.A(n_10609),
.Y(n_11494)
);

INVx2_ASAP7_75t_L g11495 ( 
.A(n_10609),
.Y(n_11495)
);

OA21x2_ASAP7_75t_L g11496 ( 
.A1(n_9808),
.A2(n_8155),
.B(n_8266),
.Y(n_11496)
);

INVx2_ASAP7_75t_L g11497 ( 
.A(n_10616),
.Y(n_11497)
);

INVx2_ASAP7_75t_L g11498 ( 
.A(n_10616),
.Y(n_11498)
);

INVx2_ASAP7_75t_L g11499 ( 
.A(n_10616),
.Y(n_11499)
);

INVx2_ASAP7_75t_L g11500 ( 
.A(n_10616),
.Y(n_11500)
);

AO21x2_ASAP7_75t_L g11501 ( 
.A1(n_10040),
.A2(n_8850),
.B(n_8157),
.Y(n_11501)
);

OAI21x1_ASAP7_75t_L g11502 ( 
.A1(n_10625),
.A2(n_10636),
.B(n_10627),
.Y(n_11502)
);

INVx2_ASAP7_75t_L g11503 ( 
.A(n_10625),
.Y(n_11503)
);

OAI21x1_ASAP7_75t_L g11504 ( 
.A1(n_10625),
.A2(n_8323),
.B(n_8305),
.Y(n_11504)
);

INVx1_ASAP7_75t_L g11505 ( 
.A(n_9877),
.Y(n_11505)
);

INVx1_ASAP7_75t_L g11506 ( 
.A(n_9878),
.Y(n_11506)
);

AND2x2_ASAP7_75t_L g11507 ( 
.A(n_11021),
.B(n_9304),
.Y(n_11507)
);

HB1xp67_ASAP7_75t_L g11508 ( 
.A(n_9591),
.Y(n_11508)
);

INVx1_ASAP7_75t_L g11509 ( 
.A(n_9878),
.Y(n_11509)
);

INVx2_ASAP7_75t_L g11510 ( 
.A(n_10625),
.Y(n_11510)
);

INVx5_ASAP7_75t_L g11511 ( 
.A(n_9764),
.Y(n_11511)
);

AND2x2_ASAP7_75t_L g11512 ( 
.A(n_11021),
.B(n_9430),
.Y(n_11512)
);

BUFx6f_ASAP7_75t_L g11513 ( 
.A(n_9764),
.Y(n_11513)
);

OAI21x1_ASAP7_75t_L g11514 ( 
.A1(n_10627),
.A2(n_8305),
.B(n_8453),
.Y(n_11514)
);

AND2x4_ASAP7_75t_L g11515 ( 
.A(n_10399),
.B(n_10442),
.Y(n_11515)
);

INVx1_ASAP7_75t_L g11516 ( 
.A(n_9885),
.Y(n_11516)
);

OAI21x1_ASAP7_75t_L g11517 ( 
.A1(n_10627),
.A2(n_8305),
.B(n_8453),
.Y(n_11517)
);

INVx1_ASAP7_75t_L g11518 ( 
.A(n_9885),
.Y(n_11518)
);

BUFx4f_ASAP7_75t_SL g11519 ( 
.A(n_10102),
.Y(n_11519)
);

INVx3_ASAP7_75t_L g11520 ( 
.A(n_9764),
.Y(n_11520)
);

OAI21x1_ASAP7_75t_L g11521 ( 
.A1(n_10627),
.A2(n_8453),
.B(n_9175),
.Y(n_11521)
);

INVx2_ASAP7_75t_L g11522 ( 
.A(n_10636),
.Y(n_11522)
);

INVx2_ASAP7_75t_L g11523 ( 
.A(n_10636),
.Y(n_11523)
);

CKINVDCx5p33_ASAP7_75t_R g11524 ( 
.A(n_10546),
.Y(n_11524)
);

HB1xp67_ASAP7_75t_L g11525 ( 
.A(n_9591),
.Y(n_11525)
);

INVx1_ASAP7_75t_L g11526 ( 
.A(n_9892),
.Y(n_11526)
);

INVx2_ASAP7_75t_L g11527 ( 
.A(n_10636),
.Y(n_11527)
);

OR2x2_ASAP7_75t_L g11528 ( 
.A(n_9599),
.B(n_8434),
.Y(n_11528)
);

INVx1_ASAP7_75t_L g11529 ( 
.A(n_9892),
.Y(n_11529)
);

INVx1_ASAP7_75t_L g11530 ( 
.A(n_9902),
.Y(n_11530)
);

OA21x2_ASAP7_75t_L g11531 ( 
.A1(n_9808),
.A2(n_8266),
.B(n_8157),
.Y(n_11531)
);

AND2x4_ASAP7_75t_L g11532 ( 
.A(n_10399),
.B(n_8346),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_9902),
.Y(n_11533)
);

INVx2_ASAP7_75t_L g11534 ( 
.A(n_10693),
.Y(n_11534)
);

OAI21x1_ASAP7_75t_L g11535 ( 
.A1(n_10693),
.A2(n_9176),
.B(n_9175),
.Y(n_11535)
);

INVx1_ASAP7_75t_L g11536 ( 
.A(n_9905),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_9905),
.Y(n_11537)
);

INVx1_ASAP7_75t_L g11538 ( 
.A(n_9907),
.Y(n_11538)
);

OAI21xp5_ASAP7_75t_L g11539 ( 
.A1(n_10164),
.A2(n_8280),
.B(n_8223),
.Y(n_11539)
);

INVx1_ASAP7_75t_L g11540 ( 
.A(n_9907),
.Y(n_11540)
);

AO21x2_ASAP7_75t_L g11541 ( 
.A1(n_9818),
.A2(n_9899),
.B(n_10509),
.Y(n_11541)
);

AO21x2_ASAP7_75t_L g11542 ( 
.A1(n_9818),
.A2(n_8157),
.B(n_9398),
.Y(n_11542)
);

INVx2_ASAP7_75t_L g11543 ( 
.A(n_10693),
.Y(n_11543)
);

INVx2_ASAP7_75t_L g11544 ( 
.A(n_10693),
.Y(n_11544)
);

INVx2_ASAP7_75t_L g11545 ( 
.A(n_10697),
.Y(n_11545)
);

AO21x1_ASAP7_75t_SL g11546 ( 
.A1(n_10972),
.A2(n_9353),
.B(n_8134),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_9912),
.Y(n_11547)
);

AOI21x1_ASAP7_75t_L g11548 ( 
.A1(n_10410),
.A2(n_9115),
.B(n_9012),
.Y(n_11548)
);

BUFx2_ASAP7_75t_L g11549 ( 
.A(n_10301),
.Y(n_11549)
);

AND2x2_ASAP7_75t_L g11550 ( 
.A(n_11021),
.B(n_9430),
.Y(n_11550)
);

INVx2_ASAP7_75t_L g11551 ( 
.A(n_10697),
.Y(n_11551)
);

INVx1_ASAP7_75t_L g11552 ( 
.A(n_9912),
.Y(n_11552)
);

INVx1_ASAP7_75t_L g11553 ( 
.A(n_9917),
.Y(n_11553)
);

INVx2_ASAP7_75t_L g11554 ( 
.A(n_10697),
.Y(n_11554)
);

INVx2_ASAP7_75t_L g11555 ( 
.A(n_10697),
.Y(n_11555)
);

AOI22xp33_ASAP7_75t_L g11556 ( 
.A1(n_10838),
.A2(n_9135),
.B1(n_9131),
.B2(n_8986),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_9917),
.Y(n_11557)
);

INVx2_ASAP7_75t_L g11558 ( 
.A(n_10333),
.Y(n_11558)
);

INVx2_ASAP7_75t_L g11559 ( 
.A(n_10333),
.Y(n_11559)
);

INVx1_ASAP7_75t_L g11560 ( 
.A(n_9921),
.Y(n_11560)
);

HB1xp67_ASAP7_75t_L g11561 ( 
.A(n_9590),
.Y(n_11561)
);

HB1xp67_ASAP7_75t_L g11562 ( 
.A(n_9590),
.Y(n_11562)
);

INVx2_ASAP7_75t_L g11563 ( 
.A(n_10333),
.Y(n_11563)
);

INVx1_ASAP7_75t_L g11564 ( 
.A(n_9921),
.Y(n_11564)
);

INVx2_ASAP7_75t_L g11565 ( 
.A(n_10333),
.Y(n_11565)
);

INVx2_ASAP7_75t_L g11566 ( 
.A(n_10422),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_9929),
.Y(n_11567)
);

INVx1_ASAP7_75t_L g11568 ( 
.A(n_9929),
.Y(n_11568)
);

OAI21x1_ASAP7_75t_L g11569 ( 
.A1(n_10405),
.A2(n_9176),
.B(n_9175),
.Y(n_11569)
);

AND2x2_ASAP7_75t_L g11570 ( 
.A(n_10742),
.B(n_9430),
.Y(n_11570)
);

INVx2_ASAP7_75t_L g11571 ( 
.A(n_10422),
.Y(n_11571)
);

INVx1_ASAP7_75t_L g11572 ( 
.A(n_9938),
.Y(n_11572)
);

BUFx2_ASAP7_75t_L g11573 ( 
.A(n_10301),
.Y(n_11573)
);

INVx2_ASAP7_75t_L g11574 ( 
.A(n_10422),
.Y(n_11574)
);

INVx2_ASAP7_75t_L g11575 ( 
.A(n_10422),
.Y(n_11575)
);

INVx1_ASAP7_75t_L g11576 ( 
.A(n_9938),
.Y(n_11576)
);

HB1xp67_ASAP7_75t_L g11577 ( 
.A(n_9590),
.Y(n_11577)
);

HB1xp67_ASAP7_75t_L g11578 ( 
.A(n_9590),
.Y(n_11578)
);

AOI21xp5_ASAP7_75t_L g11579 ( 
.A1(n_10164),
.A2(n_8556),
.B(n_8549),
.Y(n_11579)
);

INVx5_ASAP7_75t_SL g11580 ( 
.A(n_9695),
.Y(n_11580)
);

INVx1_ASAP7_75t_L g11581 ( 
.A(n_9942),
.Y(n_11581)
);

CKINVDCx11_ASAP7_75t_R g11582 ( 
.A(n_9608),
.Y(n_11582)
);

INVx2_ASAP7_75t_L g11583 ( 
.A(n_10425),
.Y(n_11583)
);

INVx1_ASAP7_75t_L g11584 ( 
.A(n_9942),
.Y(n_11584)
);

INVx1_ASAP7_75t_L g11585 ( 
.A(n_9943),
.Y(n_11585)
);

AND2x4_ASAP7_75t_L g11586 ( 
.A(n_10442),
.B(n_10952),
.Y(n_11586)
);

AO31x2_ASAP7_75t_L g11587 ( 
.A1(n_10509),
.A2(n_9432),
.A3(n_8851),
.B(n_8904),
.Y(n_11587)
);

INVx1_ASAP7_75t_L g11588 ( 
.A(n_9943),
.Y(n_11588)
);

HB1xp67_ASAP7_75t_L g11589 ( 
.A(n_9618),
.Y(n_11589)
);

OAI22xp5_ASAP7_75t_L g11590 ( 
.A1(n_10665),
.A2(n_9166),
.B1(n_8549),
.B2(n_8566),
.Y(n_11590)
);

OR2x2_ASAP7_75t_L g11591 ( 
.A(n_10980),
.B(n_8466),
.Y(n_11591)
);

INVx3_ASAP7_75t_L g11592 ( 
.A(n_9764),
.Y(n_11592)
);

AND2x4_ASAP7_75t_L g11593 ( 
.A(n_10442),
.B(n_8346),
.Y(n_11593)
);

INVx2_ASAP7_75t_L g11594 ( 
.A(n_10425),
.Y(n_11594)
);

INVx1_ASAP7_75t_L g11595 ( 
.A(n_9944),
.Y(n_11595)
);

INVx1_ASAP7_75t_L g11596 ( 
.A(n_9944),
.Y(n_11596)
);

BUFx2_ASAP7_75t_L g11597 ( 
.A(n_10301),
.Y(n_11597)
);

INVx4_ASAP7_75t_SL g11598 ( 
.A(n_9743),
.Y(n_11598)
);

AND2x2_ASAP7_75t_L g11599 ( 
.A(n_11021),
.B(n_8490),
.Y(n_11599)
);

INVx1_ASAP7_75t_L g11600 ( 
.A(n_9952),
.Y(n_11600)
);

INVx1_ASAP7_75t_L g11601 ( 
.A(n_9952),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_9955),
.Y(n_11602)
);

INVx1_ASAP7_75t_L g11603 ( 
.A(n_9955),
.Y(n_11603)
);

INVx3_ASAP7_75t_L g11604 ( 
.A(n_10229),
.Y(n_11604)
);

OAI21x1_ASAP7_75t_L g11605 ( 
.A1(n_10405),
.A2(n_9206),
.B(n_9176),
.Y(n_11605)
);

OAI22xp5_ASAP7_75t_L g11606 ( 
.A1(n_10366),
.A2(n_8566),
.B1(n_8806),
.B2(n_8609),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_9962),
.Y(n_11607)
);

INVx2_ASAP7_75t_SL g11608 ( 
.A(n_10677),
.Y(n_11608)
);

AND2x4_ASAP7_75t_L g11609 ( 
.A(n_10442),
.B(n_8366),
.Y(n_11609)
);

INVx2_ASAP7_75t_L g11610 ( 
.A(n_10425),
.Y(n_11610)
);

INVx1_ASAP7_75t_L g11611 ( 
.A(n_9962),
.Y(n_11611)
);

INVx3_ASAP7_75t_L g11612 ( 
.A(n_10229),
.Y(n_11612)
);

AOI22xp33_ASAP7_75t_L g11613 ( 
.A1(n_10852),
.A2(n_8986),
.B1(n_8985),
.B2(n_8182),
.Y(n_11613)
);

HB1xp67_ASAP7_75t_L g11614 ( 
.A(n_9634),
.Y(n_11614)
);

HB1xp67_ASAP7_75t_L g11615 ( 
.A(n_9689),
.Y(n_11615)
);

INVx2_ASAP7_75t_L g11616 ( 
.A(n_10425),
.Y(n_11616)
);

AND2x2_ASAP7_75t_L g11617 ( 
.A(n_11021),
.B(n_8490),
.Y(n_11617)
);

INVx1_ASAP7_75t_L g11618 ( 
.A(n_9964),
.Y(n_11618)
);

OR2x6_ASAP7_75t_L g11619 ( 
.A(n_9626),
.B(n_8793),
.Y(n_11619)
);

INVx1_ASAP7_75t_L g11620 ( 
.A(n_9964),
.Y(n_11620)
);

INVx1_ASAP7_75t_L g11621 ( 
.A(n_9975),
.Y(n_11621)
);

INVx1_ASAP7_75t_L g11622 ( 
.A(n_9975),
.Y(n_11622)
);

AND2x2_ASAP7_75t_L g11623 ( 
.A(n_10742),
.B(n_8490),
.Y(n_11623)
);

HB1xp67_ASAP7_75t_L g11624 ( 
.A(n_9690),
.Y(n_11624)
);

BUFx3_ASAP7_75t_L g11625 ( 
.A(n_10102),
.Y(n_11625)
);

INVx1_ASAP7_75t_L g11626 ( 
.A(n_9978),
.Y(n_11626)
);

AND2x2_ASAP7_75t_L g11627 ( 
.A(n_10742),
.B(n_8510),
.Y(n_11627)
);

INVx1_ASAP7_75t_L g11628 ( 
.A(n_9978),
.Y(n_11628)
);

AND2x4_ASAP7_75t_L g11629 ( 
.A(n_10442),
.B(n_8366),
.Y(n_11629)
);

INVx3_ASAP7_75t_L g11630 ( 
.A(n_10229),
.Y(n_11630)
);

INVx1_ASAP7_75t_L g11631 ( 
.A(n_9981),
.Y(n_11631)
);

NAND2xp5_ASAP7_75t_L g11632 ( 
.A(n_10439),
.B(n_9529),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_9981),
.Y(n_11633)
);

INVx2_ASAP7_75t_L g11634 ( 
.A(n_10432),
.Y(n_11634)
);

OAI22xp5_ASAP7_75t_L g11635 ( 
.A1(n_10439),
.A2(n_8609),
.B1(n_8614),
.B2(n_9442),
.Y(n_11635)
);

NAND2xp5_ASAP7_75t_L g11636 ( 
.A(n_10455),
.B(n_9529),
.Y(n_11636)
);

INVxp33_ASAP7_75t_SL g11637 ( 
.A(n_10561),
.Y(n_11637)
);

AND2x2_ASAP7_75t_L g11638 ( 
.A(n_10742),
.B(n_8510),
.Y(n_11638)
);

AO31x2_ASAP7_75t_L g11639 ( 
.A1(n_10455),
.A2(n_9432),
.A3(n_8851),
.B(n_8904),
.Y(n_11639)
);

NOR2xp33_ASAP7_75t_L g11640 ( 
.A(n_10263),
.B(n_9556),
.Y(n_11640)
);

OR2x2_ASAP7_75t_L g11641 ( 
.A(n_10980),
.B(n_8466),
.Y(n_11641)
);

A2O1A1Ixp33_ASAP7_75t_L g11642 ( 
.A1(n_10852),
.A2(n_8727),
.B(n_9566),
.C(n_8476),
.Y(n_11642)
);

OAI21x1_ASAP7_75t_L g11643 ( 
.A1(n_10580),
.A2(n_9209),
.B(n_9206),
.Y(n_11643)
);

INVxp67_ASAP7_75t_L g11644 ( 
.A(n_10501),
.Y(n_11644)
);

INVx2_ASAP7_75t_L g11645 ( 
.A(n_10432),
.Y(n_11645)
);

INVx1_ASAP7_75t_L g11646 ( 
.A(n_9989),
.Y(n_11646)
);

INVx1_ASAP7_75t_L g11647 ( 
.A(n_9989),
.Y(n_11647)
);

INVx2_ASAP7_75t_L g11648 ( 
.A(n_10432),
.Y(n_11648)
);

INVx2_ASAP7_75t_L g11649 ( 
.A(n_10432),
.Y(n_11649)
);

INVx2_ASAP7_75t_L g11650 ( 
.A(n_10441),
.Y(n_11650)
);

HB1xp67_ASAP7_75t_L g11651 ( 
.A(n_9715),
.Y(n_11651)
);

INVx2_ASAP7_75t_SL g11652 ( 
.A(n_10677),
.Y(n_11652)
);

INVx3_ASAP7_75t_L g11653 ( 
.A(n_10255),
.Y(n_11653)
);

NOR2xp33_ASAP7_75t_L g11654 ( 
.A(n_10263),
.B(n_7381),
.Y(n_11654)
);

CKINVDCx5p33_ASAP7_75t_R g11655 ( 
.A(n_10566),
.Y(n_11655)
);

CKINVDCx5p33_ASAP7_75t_R g11656 ( 
.A(n_10570),
.Y(n_11656)
);

INVx1_ASAP7_75t_L g11657 ( 
.A(n_10000),
.Y(n_11657)
);

INVx1_ASAP7_75t_L g11658 ( 
.A(n_10000),
.Y(n_11658)
);

BUFx3_ASAP7_75t_L g11659 ( 
.A(n_10102),
.Y(n_11659)
);

INVx2_ASAP7_75t_L g11660 ( 
.A(n_10441),
.Y(n_11660)
);

INVx2_ASAP7_75t_L g11661 ( 
.A(n_10441),
.Y(n_11661)
);

INVx1_ASAP7_75t_L g11662 ( 
.A(n_10007),
.Y(n_11662)
);

CKINVDCx5p33_ASAP7_75t_R g11663 ( 
.A(n_10669),
.Y(n_11663)
);

OAI21x1_ASAP7_75t_L g11664 ( 
.A1(n_10580),
.A2(n_9854),
.B(n_10026),
.Y(n_11664)
);

OR2x2_ASAP7_75t_L g11665 ( 
.A(n_10473),
.B(n_8131),
.Y(n_11665)
);

AOI22xp5_ASAP7_75t_L g11666 ( 
.A1(n_10866),
.A2(n_8656),
.B1(n_8657),
.B2(n_9310),
.Y(n_11666)
);

HB1xp67_ASAP7_75t_L g11667 ( 
.A(n_9732),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_10007),
.Y(n_11668)
);

INVx2_ASAP7_75t_L g11669 ( 
.A(n_10441),
.Y(n_11669)
);

HB1xp67_ASAP7_75t_L g11670 ( 
.A(n_10760),
.Y(n_11670)
);

INVx2_ASAP7_75t_SL g11671 ( 
.A(n_10677),
.Y(n_11671)
);

OR2x2_ASAP7_75t_L g11672 ( 
.A(n_10473),
.B(n_8146),
.Y(n_11672)
);

INVx1_ASAP7_75t_L g11673 ( 
.A(n_10010),
.Y(n_11673)
);

INVx1_ASAP7_75t_L g11674 ( 
.A(n_10010),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_10471),
.Y(n_11675)
);

INVx1_ASAP7_75t_L g11676 ( 
.A(n_10013),
.Y(n_11676)
);

INVx2_ASAP7_75t_L g11677 ( 
.A(n_10471),
.Y(n_11677)
);

AND2x4_ASAP7_75t_SL g11678 ( 
.A(n_10822),
.B(n_8793),
.Y(n_11678)
);

INVx2_ASAP7_75t_SL g11679 ( 
.A(n_10677),
.Y(n_11679)
);

INVx1_ASAP7_75t_L g11680 ( 
.A(n_10013),
.Y(n_11680)
);

AND2x4_ASAP7_75t_L g11681 ( 
.A(n_10442),
.B(n_8366),
.Y(n_11681)
);

HB1xp67_ASAP7_75t_L g11682 ( 
.A(n_10778),
.Y(n_11682)
);

BUFx6f_ASAP7_75t_L g11683 ( 
.A(n_9703),
.Y(n_11683)
);

AND2x4_ASAP7_75t_L g11684 ( 
.A(n_10952),
.B(n_8366),
.Y(n_11684)
);

INVx1_ASAP7_75t_L g11685 ( 
.A(n_10014),
.Y(n_11685)
);

INVxp67_ASAP7_75t_L g11686 ( 
.A(n_10501),
.Y(n_11686)
);

INVx1_ASAP7_75t_L g11687 ( 
.A(n_10014),
.Y(n_11687)
);

AND2x2_ASAP7_75t_L g11688 ( 
.A(n_10742),
.B(n_8510),
.Y(n_11688)
);

AO21x2_ASAP7_75t_L g11689 ( 
.A1(n_10940),
.A2(n_10629),
.B(n_10620),
.Y(n_11689)
);

OA21x2_ASAP7_75t_L g11690 ( 
.A1(n_9808),
.A2(n_8149),
.B(n_8625),
.Y(n_11690)
);

INVx1_ASAP7_75t_L g11691 ( 
.A(n_10022),
.Y(n_11691)
);

INVx2_ASAP7_75t_L g11692 ( 
.A(n_10471),
.Y(n_11692)
);

INVx2_ASAP7_75t_L g11693 ( 
.A(n_10471),
.Y(n_11693)
);

AND2x2_ASAP7_75t_L g11694 ( 
.A(n_10883),
.B(n_9352),
.Y(n_11694)
);

INVx1_ASAP7_75t_L g11695 ( 
.A(n_10022),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_10030),
.Y(n_11696)
);

INVx1_ASAP7_75t_L g11697 ( 
.A(n_10030),
.Y(n_11697)
);

INVx1_ASAP7_75t_L g11698 ( 
.A(n_10031),
.Y(n_11698)
);

OAI21x1_ASAP7_75t_L g11699 ( 
.A1(n_9854),
.A2(n_9209),
.B(n_9206),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_10031),
.Y(n_11700)
);

INVx1_ASAP7_75t_L g11701 ( 
.A(n_10032),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_10032),
.Y(n_11702)
);

NAND2xp5_ASAP7_75t_L g11703 ( 
.A(n_10529),
.B(n_8959),
.Y(n_11703)
);

AOI22xp5_ASAP7_75t_L g11704 ( 
.A1(n_10866),
.A2(n_8656),
.B1(n_8657),
.B2(n_9310),
.Y(n_11704)
);

AOI22xp33_ASAP7_75t_L g11705 ( 
.A1(n_10529),
.A2(n_8985),
.B1(n_8182),
.B2(n_8245),
.Y(n_11705)
);

INVx1_ASAP7_75t_SL g11706 ( 
.A(n_10514),
.Y(n_11706)
);

HB1xp67_ASAP7_75t_L g11707 ( 
.A(n_10805),
.Y(n_11707)
);

INVx2_ASAP7_75t_L g11708 ( 
.A(n_10489),
.Y(n_11708)
);

INVx1_ASAP7_75t_L g11709 ( 
.A(n_10041),
.Y(n_11709)
);

BUFx3_ASAP7_75t_L g11710 ( 
.A(n_9608),
.Y(n_11710)
);

AOI22xp33_ASAP7_75t_L g11711 ( 
.A1(n_9974),
.A2(n_8985),
.B1(n_8182),
.B2(n_8245),
.Y(n_11711)
);

INVx2_ASAP7_75t_L g11712 ( 
.A(n_10489),
.Y(n_11712)
);

AOI22xp33_ASAP7_75t_L g11713 ( 
.A1(n_9803),
.A2(n_8985),
.B1(n_8182),
.B2(n_8245),
.Y(n_11713)
);

OAI22xp33_ASAP7_75t_L g11714 ( 
.A1(n_9652),
.A2(n_8614),
.B1(n_9482),
.B2(n_8935),
.Y(n_11714)
);

OR2x2_ASAP7_75t_L g11715 ( 
.A(n_10956),
.B(n_10978),
.Y(n_11715)
);

INVx1_ASAP7_75t_L g11716 ( 
.A(n_10041),
.Y(n_11716)
);

NAND2x1p5_ASAP7_75t_L g11717 ( 
.A(n_9759),
.B(n_9783),
.Y(n_11717)
);

AND2x2_ASAP7_75t_L g11718 ( 
.A(n_10883),
.B(n_9352),
.Y(n_11718)
);

CKINVDCx5p33_ASAP7_75t_R g11719 ( 
.A(n_10738),
.Y(n_11719)
);

OAI21xp5_ASAP7_75t_L g11720 ( 
.A1(n_10685),
.A2(n_8299),
.B(n_8223),
.Y(n_11720)
);

INVx1_ASAP7_75t_L g11721 ( 
.A(n_10094),
.Y(n_11721)
);

AOI22xp33_ASAP7_75t_L g11722 ( 
.A1(n_10685),
.A2(n_8985),
.B1(n_8182),
.B2(n_8245),
.Y(n_11722)
);

INVx2_ASAP7_75t_SL g11723 ( 
.A(n_10677),
.Y(n_11723)
);

INVx1_ASAP7_75t_L g11724 ( 
.A(n_10094),
.Y(n_11724)
);

INVx2_ASAP7_75t_L g11725 ( 
.A(n_10489),
.Y(n_11725)
);

INVx2_ASAP7_75t_L g11726 ( 
.A(n_10489),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_10098),
.Y(n_11727)
);

INVx2_ASAP7_75t_SL g11728 ( 
.A(n_10885),
.Y(n_11728)
);

INVx1_ASAP7_75t_L g11729 ( 
.A(n_10098),
.Y(n_11729)
);

HB1xp67_ASAP7_75t_L g11730 ( 
.A(n_10829),
.Y(n_11730)
);

INVx1_ASAP7_75t_L g11731 ( 
.A(n_10101),
.Y(n_11731)
);

INVx1_ASAP7_75t_L g11732 ( 
.A(n_10101),
.Y(n_11732)
);

OAI21x1_ASAP7_75t_L g11733 ( 
.A1(n_10026),
.A2(n_9221),
.B(n_9209),
.Y(n_11733)
);

INVx2_ASAP7_75t_L g11734 ( 
.A(n_10867),
.Y(n_11734)
);

INVx2_ASAP7_75t_SL g11735 ( 
.A(n_10885),
.Y(n_11735)
);

INVx2_ASAP7_75t_L g11736 ( 
.A(n_10867),
.Y(n_11736)
);

INVx1_ASAP7_75t_L g11737 ( 
.A(n_10104),
.Y(n_11737)
);

INVx2_ASAP7_75t_L g11738 ( 
.A(n_10867),
.Y(n_11738)
);

INVx1_ASAP7_75t_L g11739 ( 
.A(n_10104),
.Y(n_11739)
);

OAI21x1_ASAP7_75t_L g11740 ( 
.A1(n_9876),
.A2(n_9221),
.B(n_8411),
.Y(n_11740)
);

OAI21x1_ASAP7_75t_L g11741 ( 
.A1(n_9876),
.A2(n_9221),
.B(n_8411),
.Y(n_11741)
);

INVx2_ASAP7_75t_L g11742 ( 
.A(n_10867),
.Y(n_11742)
);

NOR2x1_ASAP7_75t_SL g11743 ( 
.A(n_11000),
.B(n_9035),
.Y(n_11743)
);

INVx2_ASAP7_75t_SL g11744 ( 
.A(n_10702),
.Y(n_11744)
);

NAND2xp5_ASAP7_75t_L g11745 ( 
.A(n_9792),
.B(n_8959),
.Y(n_11745)
);

AO21x1_ASAP7_75t_L g11746 ( 
.A1(n_10429),
.A2(n_8826),
.B(n_8740),
.Y(n_11746)
);

INVx3_ASAP7_75t_L g11747 ( 
.A(n_10255),
.Y(n_11747)
);

INVx1_ASAP7_75t_L g11748 ( 
.A(n_10109),
.Y(n_11748)
);

HB1xp67_ASAP7_75t_L g11749 ( 
.A(n_10871),
.Y(n_11749)
);

A2O1A1Ixp33_ASAP7_75t_L g11750 ( 
.A1(n_9862),
.A2(n_8727),
.B(n_9306),
.C(n_8734),
.Y(n_11750)
);

BUFx3_ASAP7_75t_L g11751 ( 
.A(n_9932),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_10109),
.Y(n_11752)
);

OAI21x1_ASAP7_75t_L g11753 ( 
.A1(n_9880),
.A2(n_9923),
.B(n_9701),
.Y(n_11753)
);

OR2x2_ASAP7_75t_L g11754 ( 
.A(n_10956),
.B(n_8146),
.Y(n_11754)
);

BUFx2_ASAP7_75t_L g11755 ( 
.A(n_9935),
.Y(n_11755)
);

INVxp67_ASAP7_75t_R g11756 ( 
.A(n_10933),
.Y(n_11756)
);

INVxp67_ASAP7_75t_SL g11757 ( 
.A(n_9625),
.Y(n_11757)
);

INVx3_ASAP7_75t_L g11758 ( 
.A(n_10255),
.Y(n_11758)
);

INVx1_ASAP7_75t_L g11759 ( 
.A(n_10112),
.Y(n_11759)
);

OAI22xp5_ASAP7_75t_L g11760 ( 
.A1(n_10923),
.A2(n_9442),
.B1(n_9035),
.B2(n_9076),
.Y(n_11760)
);

AND2x4_ASAP7_75t_SL g11761 ( 
.A(n_10822),
.B(n_8851),
.Y(n_11761)
);

INVx2_ASAP7_75t_L g11762 ( 
.A(n_10921),
.Y(n_11762)
);

INVx2_ASAP7_75t_L g11763 ( 
.A(n_10921),
.Y(n_11763)
);

HB1xp67_ASAP7_75t_L g11764 ( 
.A(n_10881),
.Y(n_11764)
);

INVx2_ASAP7_75t_L g11765 ( 
.A(n_10921),
.Y(n_11765)
);

INVx1_ASAP7_75t_L g11766 ( 
.A(n_10112),
.Y(n_11766)
);

INVx2_ASAP7_75t_L g11767 ( 
.A(n_10921),
.Y(n_11767)
);

INVx2_ASAP7_75t_L g11768 ( 
.A(n_10729),
.Y(n_11768)
);

INVx1_ASAP7_75t_L g11769 ( 
.A(n_10119),
.Y(n_11769)
);

NAND2x1p5_ASAP7_75t_L g11770 ( 
.A(n_9759),
.B(n_8851),
.Y(n_11770)
);

AND2x2_ASAP7_75t_L g11771 ( 
.A(n_10883),
.B(n_9396),
.Y(n_11771)
);

INVx1_ASAP7_75t_L g11772 ( 
.A(n_10119),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_10120),
.Y(n_11773)
);

INVx1_ASAP7_75t_L g11774 ( 
.A(n_10120),
.Y(n_11774)
);

OAI21xp5_ASAP7_75t_L g11775 ( 
.A1(n_9617),
.A2(n_9809),
.B(n_9797),
.Y(n_11775)
);

INVx1_ASAP7_75t_L g11776 ( 
.A(n_10127),
.Y(n_11776)
);

NOR2xp33_ASAP7_75t_L g11777 ( 
.A(n_10278),
.B(n_7776),
.Y(n_11777)
);

AND2x2_ASAP7_75t_L g11778 ( 
.A(n_10883),
.B(n_9396),
.Y(n_11778)
);

AO21x2_ASAP7_75t_L g11779 ( 
.A1(n_10940),
.A2(n_10629),
.B(n_10620),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_10127),
.Y(n_11780)
);

OR2x2_ASAP7_75t_L g11781 ( 
.A(n_10978),
.B(n_8163),
.Y(n_11781)
);

INVx2_ASAP7_75t_L g11782 ( 
.A(n_10729),
.Y(n_11782)
);

OAI22xp33_ASAP7_75t_L g11783 ( 
.A1(n_9652),
.A2(n_9482),
.B1(n_8829),
.B2(n_8935),
.Y(n_11783)
);

INVx6_ASAP7_75t_L g11784 ( 
.A(n_9932),
.Y(n_11784)
);

INVx1_ASAP7_75t_L g11785 ( 
.A(n_10130),
.Y(n_11785)
);

INVx2_ASAP7_75t_L g11786 ( 
.A(n_10729),
.Y(n_11786)
);

INVx1_ASAP7_75t_L g11787 ( 
.A(n_10130),
.Y(n_11787)
);

HB1xp67_ASAP7_75t_L g11788 ( 
.A(n_10964),
.Y(n_11788)
);

BUFx2_ASAP7_75t_L g11789 ( 
.A(n_9935),
.Y(n_11789)
);

OAI21xp5_ASAP7_75t_L g11790 ( 
.A1(n_9617),
.A2(n_8299),
.B(n_8779),
.Y(n_11790)
);

INVxp67_ASAP7_75t_L g11791 ( 
.A(n_10724),
.Y(n_11791)
);

INVx1_ASAP7_75t_L g11792 ( 
.A(n_10136),
.Y(n_11792)
);

INVx1_ASAP7_75t_L g11793 ( 
.A(n_10136),
.Y(n_11793)
);

INVx3_ASAP7_75t_L g11794 ( 
.A(n_9592),
.Y(n_11794)
);

INVx1_ASAP7_75t_L g11795 ( 
.A(n_10146),
.Y(n_11795)
);

AO31x2_ASAP7_75t_L g11796 ( 
.A1(n_10519),
.A2(n_8904),
.A3(n_9060),
.B(n_8851),
.Y(n_11796)
);

AND2x4_ASAP7_75t_L g11797 ( 
.A(n_10952),
.B(n_8378),
.Y(n_11797)
);

INVx2_ASAP7_75t_SL g11798 ( 
.A(n_10702),
.Y(n_11798)
);

INVx1_ASAP7_75t_L g11799 ( 
.A(n_10146),
.Y(n_11799)
);

HB1xp67_ASAP7_75t_L g11800 ( 
.A(n_10713),
.Y(n_11800)
);

NAND2xp5_ASAP7_75t_L g11801 ( 
.A(n_9792),
.B(n_8572),
.Y(n_11801)
);

HB1xp67_ASAP7_75t_L g11802 ( 
.A(n_10723),
.Y(n_11802)
);

NAND2xp5_ASAP7_75t_L g11803 ( 
.A(n_10628),
.B(n_8572),
.Y(n_11803)
);

INVx2_ASAP7_75t_L g11804 ( 
.A(n_10737),
.Y(n_11804)
);

OAI21xp5_ASAP7_75t_L g11805 ( 
.A1(n_9797),
.A2(n_8800),
.B(n_8779),
.Y(n_11805)
);

HB1xp67_ASAP7_75t_L g11806 ( 
.A(n_10743),
.Y(n_11806)
);

OR2x6_ASAP7_75t_L g11807 ( 
.A(n_9856),
.B(n_8904),
.Y(n_11807)
);

INVx2_ASAP7_75t_L g11808 ( 
.A(n_10737),
.Y(n_11808)
);

INVx2_ASAP7_75t_L g11809 ( 
.A(n_10737),
.Y(n_11809)
);

AOI21x1_ASAP7_75t_L g11810 ( 
.A1(n_9727),
.A2(n_9115),
.B(n_9012),
.Y(n_11810)
);

INVx2_ASAP7_75t_L g11811 ( 
.A(n_9888),
.Y(n_11811)
);

INVx1_ASAP7_75t_L g11812 ( 
.A(n_10153),
.Y(n_11812)
);

NAND2xp5_ASAP7_75t_L g11813 ( 
.A(n_10116),
.B(n_8572),
.Y(n_11813)
);

BUFx3_ASAP7_75t_L g11814 ( 
.A(n_9932),
.Y(n_11814)
);

AND2x2_ASAP7_75t_L g11815 ( 
.A(n_10883),
.B(n_8164),
.Y(n_11815)
);

BUFx2_ASAP7_75t_L g11816 ( 
.A(n_9935),
.Y(n_11816)
);

BUFx4f_ASAP7_75t_SL g11817 ( 
.A(n_9695),
.Y(n_11817)
);

NAND2x1p5_ASAP7_75t_L g11818 ( 
.A(n_9759),
.B(n_8904),
.Y(n_11818)
);

AOI21x1_ASAP7_75t_L g11819 ( 
.A1(n_9727),
.A2(n_9115),
.B(n_9012),
.Y(n_11819)
);

INVx1_ASAP7_75t_L g11820 ( 
.A(n_10153),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_10156),
.Y(n_11821)
);

HB1xp67_ASAP7_75t_L g11822 ( 
.A(n_10156),
.Y(n_11822)
);

AND2x4_ASAP7_75t_L g11823 ( 
.A(n_10952),
.B(n_8378),
.Y(n_11823)
);

INVx2_ASAP7_75t_L g11824 ( 
.A(n_9888),
.Y(n_11824)
);

INVx2_ASAP7_75t_L g11825 ( 
.A(n_9888),
.Y(n_11825)
);

NAND2xp5_ASAP7_75t_L g11826 ( 
.A(n_10116),
.B(n_8572),
.Y(n_11826)
);

INVx1_ASAP7_75t_L g11827 ( 
.A(n_10166),
.Y(n_11827)
);

INVx1_ASAP7_75t_L g11828 ( 
.A(n_10166),
.Y(n_11828)
);

OAI21xp5_ASAP7_75t_L g11829 ( 
.A1(n_9809),
.A2(n_8800),
.B(n_8769),
.Y(n_11829)
);

NOR2xp33_ASAP7_75t_L g11830 ( 
.A(n_10278),
.B(n_7899),
.Y(n_11830)
);

AOI21x1_ASAP7_75t_L g11831 ( 
.A1(n_9890),
.A2(n_9923),
.B(n_9598),
.Y(n_11831)
);

AND2x4_ASAP7_75t_L g11832 ( 
.A(n_10952),
.B(n_9631),
.Y(n_11832)
);

INVx2_ASAP7_75t_L g11833 ( 
.A(n_9888),
.Y(n_11833)
);

INVx1_ASAP7_75t_L g11834 ( 
.A(n_10172),
.Y(n_11834)
);

INVx1_ASAP7_75t_L g11835 ( 
.A(n_10172),
.Y(n_11835)
);

AND2x4_ASAP7_75t_L g11836 ( 
.A(n_10952),
.B(n_8378),
.Y(n_11836)
);

OR2x2_ASAP7_75t_L g11837 ( 
.A(n_10272),
.B(n_8163),
.Y(n_11837)
);

INVx1_ASAP7_75t_SL g11838 ( 
.A(n_10514),
.Y(n_11838)
);

AOI22xp33_ASAP7_75t_L g11839 ( 
.A1(n_10348),
.A2(n_8182),
.B1(n_8245),
.B2(n_8226),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_10176),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_9949),
.Y(n_11841)
);

AO21x2_ASAP7_75t_L g11842 ( 
.A1(n_10849),
.A2(n_9413),
.B(n_9398),
.Y(n_11842)
);

OAI21x1_ASAP7_75t_L g11843 ( 
.A1(n_9880),
.A2(n_8411),
.B(n_8734),
.Y(n_11843)
);

BUFx2_ASAP7_75t_L g11844 ( 
.A(n_9935),
.Y(n_11844)
);

AND2x2_ASAP7_75t_L g11845 ( 
.A(n_10969),
.B(n_8164),
.Y(n_11845)
);

INVx2_ASAP7_75t_L g11846 ( 
.A(n_9949),
.Y(n_11846)
);

BUFx2_ASAP7_75t_L g11847 ( 
.A(n_10018),
.Y(n_11847)
);

AOI22xp33_ASAP7_75t_L g11848 ( 
.A1(n_10651),
.A2(n_8245),
.B1(n_8226),
.B2(n_9199),
.Y(n_11848)
);

INVx2_ASAP7_75t_L g11849 ( 
.A(n_9949),
.Y(n_11849)
);

INVx1_ASAP7_75t_L g11850 ( 
.A(n_10176),
.Y(n_11850)
);

INVx2_ASAP7_75t_L g11851 ( 
.A(n_9949),
.Y(n_11851)
);

INVx2_ASAP7_75t_L g11852 ( 
.A(n_9960),
.Y(n_11852)
);

AO21x1_ASAP7_75t_SL g11853 ( 
.A1(n_10972),
.A2(n_8134),
.B(n_8624),
.Y(n_11853)
);

INVx2_ASAP7_75t_L g11854 ( 
.A(n_9960),
.Y(n_11854)
);

INVx1_ASAP7_75t_L g11855 ( 
.A(n_10177),
.Y(n_11855)
);

NAND2xp5_ASAP7_75t_L g11856 ( 
.A(n_10202),
.B(n_8572),
.Y(n_11856)
);

INVx3_ASAP7_75t_L g11857 ( 
.A(n_9592),
.Y(n_11857)
);

OAI22xp5_ASAP7_75t_L g11858 ( 
.A1(n_10923),
.A2(n_10958),
.B1(n_10429),
.B2(n_10337),
.Y(n_11858)
);

INVx1_ASAP7_75t_L g11859 ( 
.A(n_10177),
.Y(n_11859)
);

INVx2_ASAP7_75t_SL g11860 ( 
.A(n_10702),
.Y(n_11860)
);

OAI22xp5_ASAP7_75t_L g11861 ( 
.A1(n_10337),
.A2(n_9862),
.B1(n_9760),
.B2(n_9781),
.Y(n_11861)
);

OAI222xp33_ASAP7_75t_L g11862 ( 
.A1(n_10699),
.A2(n_9109),
.B1(n_8944),
.B2(n_8666),
.C1(n_8673),
.C2(n_8716),
.Y(n_11862)
);

AOI21x1_ASAP7_75t_L g11863 ( 
.A1(n_9890),
.A2(n_9266),
.B(n_9190),
.Y(n_11863)
);

INVx1_ASAP7_75t_L g11864 ( 
.A(n_10188),
.Y(n_11864)
);

AND2x2_ASAP7_75t_L g11865 ( 
.A(n_10969),
.B(n_8164),
.Y(n_11865)
);

OAI21xp5_ASAP7_75t_L g11866 ( 
.A1(n_10708),
.A2(n_8769),
.B(n_9167),
.Y(n_11866)
);

INVx2_ASAP7_75t_L g11867 ( 
.A(n_9960),
.Y(n_11867)
);

AO21x2_ASAP7_75t_L g11868 ( 
.A1(n_10849),
.A2(n_9413),
.B(n_9398),
.Y(n_11868)
);

NAND2xp5_ASAP7_75t_L g11869 ( 
.A(n_10202),
.B(n_8576),
.Y(n_11869)
);

OA21x2_ASAP7_75t_L g11870 ( 
.A1(n_9829),
.A2(n_8149),
.B(n_8625),
.Y(n_11870)
);

INVx2_ASAP7_75t_L g11871 ( 
.A(n_9960),
.Y(n_11871)
);

INVx1_ASAP7_75t_L g11872 ( 
.A(n_10188),
.Y(n_11872)
);

BUFx2_ASAP7_75t_L g11873 ( 
.A(n_10018),
.Y(n_11873)
);

INVx2_ASAP7_75t_L g11874 ( 
.A(n_9994),
.Y(n_11874)
);

INVx1_ASAP7_75t_L g11875 ( 
.A(n_10192),
.Y(n_11875)
);

INVx1_ASAP7_75t_L g11876 ( 
.A(n_10192),
.Y(n_11876)
);

INVx4_ASAP7_75t_L g11877 ( 
.A(n_9759),
.Y(n_11877)
);

INVx1_ASAP7_75t_L g11878 ( 
.A(n_10199),
.Y(n_11878)
);

NOR2xp33_ASAP7_75t_L g11879 ( 
.A(n_10018),
.B(n_7899),
.Y(n_11879)
);

INVx3_ASAP7_75t_L g11880 ( 
.A(n_9592),
.Y(n_11880)
);

INVx1_ASAP7_75t_L g11881 ( 
.A(n_10199),
.Y(n_11881)
);

OAI221xp5_ASAP7_75t_L g11882 ( 
.A1(n_10368),
.A2(n_9505),
.B1(n_9491),
.B2(n_8624),
.C(n_9167),
.Y(n_11882)
);

AND2x2_ASAP7_75t_L g11883 ( 
.A(n_10969),
.B(n_8164),
.Y(n_11883)
);

INVx2_ASAP7_75t_L g11884 ( 
.A(n_9994),
.Y(n_11884)
);

AND2x2_ASAP7_75t_L g11885 ( 
.A(n_10969),
.B(n_8164),
.Y(n_11885)
);

INVx2_ASAP7_75t_L g11886 ( 
.A(n_9994),
.Y(n_11886)
);

AND2x2_ASAP7_75t_L g11887 ( 
.A(n_10969),
.B(n_8203),
.Y(n_11887)
);

INVx1_ASAP7_75t_L g11888 ( 
.A(n_10200),
.Y(n_11888)
);

OAI21x1_ASAP7_75t_L g11889 ( 
.A1(n_9701),
.A2(n_9418),
.B(n_8603),
.Y(n_11889)
);

A2O1A1Ixp33_ASAP7_75t_L g11890 ( 
.A1(n_10699),
.A2(n_9306),
.B(n_9109),
.C(n_8944),
.Y(n_11890)
);

AND2x2_ASAP7_75t_L g11891 ( 
.A(n_11005),
.B(n_8203),
.Y(n_11891)
);

BUFx3_ASAP7_75t_L g11892 ( 
.A(n_9932),
.Y(n_11892)
);

OR2x2_ASAP7_75t_L g11893 ( 
.A(n_10272),
.B(n_9042),
.Y(n_11893)
);

OAI21x1_ASAP7_75t_L g11894 ( 
.A1(n_9958),
.A2(n_9418),
.B(n_8603),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_10200),
.Y(n_11895)
);

HB1xp67_ASAP7_75t_L g11896 ( 
.A(n_10218),
.Y(n_11896)
);

CKINVDCx8_ASAP7_75t_R g11897 ( 
.A(n_10724),
.Y(n_11897)
);

AND2x4_ASAP7_75t_L g11898 ( 
.A(n_10952),
.B(n_8378),
.Y(n_11898)
);

OR2x6_ASAP7_75t_L g11899 ( 
.A(n_9856),
.B(n_9060),
.Y(n_11899)
);

NAND2xp5_ASAP7_75t_L g11900 ( 
.A(n_10254),
.B(n_8576),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_10218),
.Y(n_11901)
);

INVx3_ASAP7_75t_L g11902 ( 
.A(n_9620),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_10220),
.Y(n_11903)
);

HB1xp67_ASAP7_75t_L g11904 ( 
.A(n_10220),
.Y(n_11904)
);

AND2x2_ASAP7_75t_L g11905 ( 
.A(n_11005),
.B(n_8203),
.Y(n_11905)
);

AND2x2_ASAP7_75t_L g11906 ( 
.A(n_11005),
.B(n_8203),
.Y(n_11906)
);

BUFx2_ASAP7_75t_L g11907 ( 
.A(n_10018),
.Y(n_11907)
);

OAI21x1_ASAP7_75t_L g11908 ( 
.A1(n_9958),
.A2(n_9418),
.B(n_8603),
.Y(n_11908)
);

INVx2_ASAP7_75t_L g11909 ( 
.A(n_9994),
.Y(n_11909)
);

INVx1_ASAP7_75t_L g11910 ( 
.A(n_10226),
.Y(n_11910)
);

NAND2xp5_ASAP7_75t_L g11911 ( 
.A(n_10254),
.B(n_8576),
.Y(n_11911)
);

INVx1_ASAP7_75t_L g11912 ( 
.A(n_10226),
.Y(n_11912)
);

BUFx2_ASAP7_75t_L g11913 ( 
.A(n_9992),
.Y(n_11913)
);

HB1xp67_ASAP7_75t_L g11914 ( 
.A(n_10234),
.Y(n_11914)
);

INVx1_ASAP7_75t_L g11915 ( 
.A(n_10234),
.Y(n_11915)
);

OAI21x1_ASAP7_75t_L g11916 ( 
.A1(n_9958),
.A2(n_10705),
.B(n_10637),
.Y(n_11916)
);

AND2x2_ASAP7_75t_L g11917 ( 
.A(n_11005),
.B(n_8203),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_10236),
.Y(n_11918)
);

INVx1_ASAP7_75t_L g11919 ( 
.A(n_10236),
.Y(n_11919)
);

INVx2_ASAP7_75t_L g11920 ( 
.A(n_10049),
.Y(n_11920)
);

BUFx4f_ASAP7_75t_L g11921 ( 
.A(n_9703),
.Y(n_11921)
);

AO21x2_ASAP7_75t_L g11922 ( 
.A1(n_10897),
.A2(n_9413),
.B(n_9398),
.Y(n_11922)
);

INVx1_ASAP7_75t_L g11923 ( 
.A(n_10238),
.Y(n_11923)
);

OAI21x1_ASAP7_75t_L g11924 ( 
.A1(n_10637),
.A2(n_8320),
.B(n_8796),
.Y(n_11924)
);

INVx2_ASAP7_75t_L g11925 ( 
.A(n_10049),
.Y(n_11925)
);

INVx2_ASAP7_75t_L g11926 ( 
.A(n_10049),
.Y(n_11926)
);

BUFx2_ASAP7_75t_L g11927 ( 
.A(n_9992),
.Y(n_11927)
);

INVx1_ASAP7_75t_L g11928 ( 
.A(n_10238),
.Y(n_11928)
);

OAI21x1_ASAP7_75t_L g11929 ( 
.A1(n_10705),
.A2(n_8320),
.B(n_8796),
.Y(n_11929)
);

INVx1_ASAP7_75t_L g11930 ( 
.A(n_10239),
.Y(n_11930)
);

HB1xp67_ASAP7_75t_L g11931 ( 
.A(n_10239),
.Y(n_11931)
);

INVx1_ASAP7_75t_L g11932 ( 
.A(n_10241),
.Y(n_11932)
);

INVxp67_ASAP7_75t_SL g11933 ( 
.A(n_10897),
.Y(n_11933)
);

OR2x2_ASAP7_75t_L g11934 ( 
.A(n_10840),
.B(n_9042),
.Y(n_11934)
);

INVx1_ASAP7_75t_L g11935 ( 
.A(n_10241),
.Y(n_11935)
);

INVx2_ASAP7_75t_L g11936 ( 
.A(n_10049),
.Y(n_11936)
);

INVx2_ASAP7_75t_L g11937 ( 
.A(n_10052),
.Y(n_11937)
);

INVx1_ASAP7_75t_L g11938 ( 
.A(n_10243),
.Y(n_11938)
);

INVx2_ASAP7_75t_L g11939 ( 
.A(n_10052),
.Y(n_11939)
);

OAI21x1_ASAP7_75t_SL g11940 ( 
.A1(n_9896),
.A2(n_8260),
.B(n_8796),
.Y(n_11940)
);

INVx1_ASAP7_75t_L g11941 ( 
.A(n_10243),
.Y(n_11941)
);

INVx4_ASAP7_75t_L g11942 ( 
.A(n_9759),
.Y(n_11942)
);

HB1xp67_ASAP7_75t_L g11943 ( 
.A(n_10245),
.Y(n_11943)
);

INVx1_ASAP7_75t_L g11944 ( 
.A(n_10245),
.Y(n_11944)
);

INVx2_ASAP7_75t_SL g11945 ( 
.A(n_10702),
.Y(n_11945)
);

NAND2xp5_ASAP7_75t_L g11946 ( 
.A(n_10503),
.B(n_8576),
.Y(n_11946)
);

INVx1_ASAP7_75t_L g11947 ( 
.A(n_10249),
.Y(n_11947)
);

A2O1A1Ixp33_ASAP7_75t_L g11948 ( 
.A1(n_9699),
.A2(n_8873),
.B(n_8994),
.C(n_8859),
.Y(n_11948)
);

HB1xp67_ASAP7_75t_L g11949 ( 
.A(n_10249),
.Y(n_11949)
);

AND2x4_ASAP7_75t_L g11950 ( 
.A(n_9631),
.B(n_8455),
.Y(n_11950)
);

INVx1_ASAP7_75t_L g11951 ( 
.A(n_10253),
.Y(n_11951)
);

INVx2_ASAP7_75t_L g11952 ( 
.A(n_10052),
.Y(n_11952)
);

BUFx2_ASAP7_75t_L g11953 ( 
.A(n_9992),
.Y(n_11953)
);

INVx1_ASAP7_75t_L g11954 ( 
.A(n_10253),
.Y(n_11954)
);

AOI21x1_ASAP7_75t_L g11955 ( 
.A1(n_9584),
.A2(n_9266),
.B(n_9190),
.Y(n_11955)
);

INVx1_ASAP7_75t_L g11956 ( 
.A(n_10256),
.Y(n_11956)
);

INVx1_ASAP7_75t_L g11957 ( 
.A(n_10256),
.Y(n_11957)
);

INVx1_ASAP7_75t_L g11958 ( 
.A(n_10261),
.Y(n_11958)
);

INVx2_ASAP7_75t_L g11959 ( 
.A(n_10052),
.Y(n_11959)
);

AND2x4_ASAP7_75t_L g11960 ( 
.A(n_9584),
.B(n_8455),
.Y(n_11960)
);

AND2x2_ASAP7_75t_L g11961 ( 
.A(n_11005),
.B(n_8203),
.Y(n_11961)
);

NAND2xp5_ASAP7_75t_L g11962 ( 
.A(n_10503),
.B(n_8576),
.Y(n_11962)
);

INVx1_ASAP7_75t_L g11963 ( 
.A(n_10261),
.Y(n_11963)
);

BUFx2_ASAP7_75t_L g11964 ( 
.A(n_9992),
.Y(n_11964)
);

OA21x2_ASAP7_75t_L g11965 ( 
.A1(n_9829),
.A2(n_8149),
.B(n_8625),
.Y(n_11965)
);

BUFx2_ASAP7_75t_L g11966 ( 
.A(n_10028),
.Y(n_11966)
);

INVx2_ASAP7_75t_L g11967 ( 
.A(n_10336),
.Y(n_11967)
);

INVx1_ASAP7_75t_L g11968 ( 
.A(n_10262),
.Y(n_11968)
);

INVx6_ASAP7_75t_L g11969 ( 
.A(n_10028),
.Y(n_11969)
);

BUFx6f_ASAP7_75t_L g11970 ( 
.A(n_9703),
.Y(n_11970)
);

INVx1_ASAP7_75t_L g11971 ( 
.A(n_10262),
.Y(n_11971)
);

AND2x2_ASAP7_75t_L g11972 ( 
.A(n_10420),
.B(n_8216),
.Y(n_11972)
);

INVx1_ASAP7_75t_L g11973 ( 
.A(n_10264),
.Y(n_11973)
);

INVxp67_ASAP7_75t_L g11974 ( 
.A(n_9969),
.Y(n_11974)
);

INVx1_ASAP7_75t_L g11975 ( 
.A(n_10264),
.Y(n_11975)
);

INVx1_ASAP7_75t_L g11976 ( 
.A(n_10266),
.Y(n_11976)
);

BUFx6f_ASAP7_75t_L g11977 ( 
.A(n_9620),
.Y(n_11977)
);

INVx1_ASAP7_75t_L g11978 ( 
.A(n_10266),
.Y(n_11978)
);

BUFx10_ASAP7_75t_L g11979 ( 
.A(n_9856),
.Y(n_11979)
);

INVxp67_ASAP7_75t_SL g11980 ( 
.A(n_10681),
.Y(n_11980)
);

HB1xp67_ASAP7_75t_L g11981 ( 
.A(n_10276),
.Y(n_11981)
);

CKINVDCx20_ASAP7_75t_R g11982 ( 
.A(n_9676),
.Y(n_11982)
);

AO21x2_ASAP7_75t_L g11983 ( 
.A1(n_9996),
.A2(n_9413),
.B(n_9398),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_10276),
.Y(n_11984)
);

INVx2_ASAP7_75t_L g11985 ( 
.A(n_10336),
.Y(n_11985)
);

INVx2_ASAP7_75t_SL g11986 ( 
.A(n_10028),
.Y(n_11986)
);

BUFx6f_ASAP7_75t_L g11987 ( 
.A(n_9620),
.Y(n_11987)
);

INVx2_ASAP7_75t_L g11988 ( 
.A(n_10336),
.Y(n_11988)
);

INVx1_ASAP7_75t_L g11989 ( 
.A(n_10279),
.Y(n_11989)
);

INVxp67_ASAP7_75t_L g11990 ( 
.A(n_9969),
.Y(n_11990)
);

INVx2_ASAP7_75t_SL g11991 ( 
.A(n_10028),
.Y(n_11991)
);

INVx2_ASAP7_75t_SL g11992 ( 
.A(n_10043),
.Y(n_11992)
);

INVx2_ASAP7_75t_L g11993 ( 
.A(n_10339),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_10279),
.Y(n_11994)
);

INVx3_ASAP7_75t_L g11995 ( 
.A(n_9681),
.Y(n_11995)
);

INVx4_ASAP7_75t_SL g11996 ( 
.A(n_10321),
.Y(n_11996)
);

BUFx2_ASAP7_75t_L g11997 ( 
.A(n_10043),
.Y(n_11997)
);

INVx2_ASAP7_75t_L g11998 ( 
.A(n_10339),
.Y(n_11998)
);

OR2x2_ASAP7_75t_L g11999 ( 
.A(n_10840),
.B(n_8744),
.Y(n_11999)
);

INVx1_ASAP7_75t_L g12000 ( 
.A(n_10282),
.Y(n_12000)
);

AND2x2_ASAP7_75t_L g12001 ( 
.A(n_10420),
.B(n_8216),
.Y(n_12001)
);

INVx3_ASAP7_75t_L g12002 ( 
.A(n_9681),
.Y(n_12002)
);

INVx2_ASAP7_75t_L g12003 ( 
.A(n_10339),
.Y(n_12003)
);

NAND2xp5_ASAP7_75t_L g12004 ( 
.A(n_10497),
.B(n_8576),
.Y(n_12004)
);

OAI21xp5_ASAP7_75t_L g12005 ( 
.A1(n_10708),
.A2(n_8987),
.B(n_8971),
.Y(n_12005)
);

INVx1_ASAP7_75t_L g12006 ( 
.A(n_10282),
.Y(n_12006)
);

BUFx6f_ASAP7_75t_L g12007 ( 
.A(n_9681),
.Y(n_12007)
);

INVx1_ASAP7_75t_L g12008 ( 
.A(n_10286),
.Y(n_12008)
);

INVx1_ASAP7_75t_L g12009 ( 
.A(n_10286),
.Y(n_12009)
);

INVx1_ASAP7_75t_L g12010 ( 
.A(n_10289),
.Y(n_12010)
);

OA21x2_ASAP7_75t_L g12011 ( 
.A1(n_9829),
.A2(n_8463),
.B(n_8178),
.Y(n_12011)
);

AO21x2_ASAP7_75t_L g12012 ( 
.A1(n_9996),
.A2(n_9413),
.B(n_9027),
.Y(n_12012)
);

INVx1_ASAP7_75t_L g12013 ( 
.A(n_10289),
.Y(n_12013)
);

INVx1_ASAP7_75t_L g12014 ( 
.A(n_10291),
.Y(n_12014)
);

INVx1_ASAP7_75t_L g12015 ( 
.A(n_10291),
.Y(n_12015)
);

AND2x2_ASAP7_75t_L g12016 ( 
.A(n_10531),
.B(n_8216),
.Y(n_12016)
);

NOR2xp33_ASAP7_75t_L g12017 ( 
.A(n_10059),
.B(n_9339),
.Y(n_12017)
);

INVx1_ASAP7_75t_L g12018 ( 
.A(n_10307),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_10307),
.Y(n_12019)
);

INVx1_ASAP7_75t_L g12020 ( 
.A(n_10315),
.Y(n_12020)
);

NAND2xp5_ASAP7_75t_L g12021 ( 
.A(n_10497),
.B(n_8576),
.Y(n_12021)
);

BUFx2_ASAP7_75t_L g12022 ( 
.A(n_10043),
.Y(n_12022)
);

INVx2_ASAP7_75t_L g12023 ( 
.A(n_10343),
.Y(n_12023)
);

INVx1_ASAP7_75t_L g12024 ( 
.A(n_10315),
.Y(n_12024)
);

AND2x2_ASAP7_75t_L g12025 ( 
.A(n_10531),
.B(n_8216),
.Y(n_12025)
);

INVx1_ASAP7_75t_L g12026 ( 
.A(n_10319),
.Y(n_12026)
);

INVx2_ASAP7_75t_L g12027 ( 
.A(n_10343),
.Y(n_12027)
);

OR2x2_ASAP7_75t_L g12028 ( 
.A(n_10393),
.B(n_8744),
.Y(n_12028)
);

INVx1_ASAP7_75t_L g12029 ( 
.A(n_10319),
.Y(n_12029)
);

INVx3_ASAP7_75t_L g12030 ( 
.A(n_9717),
.Y(n_12030)
);

AOI22xp33_ASAP7_75t_SL g12031 ( 
.A1(n_10518),
.A2(n_8297),
.B1(n_8640),
.B2(n_8621),
.Y(n_12031)
);

INVx4_ASAP7_75t_L g12032 ( 
.A(n_9759),
.Y(n_12032)
);

BUFx3_ASAP7_75t_L g12033 ( 
.A(n_10043),
.Y(n_12033)
);

INVx1_ASAP7_75t_L g12034 ( 
.A(n_10326),
.Y(n_12034)
);

INVx1_ASAP7_75t_L g12035 ( 
.A(n_10326),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_10330),
.Y(n_12036)
);

AND2x2_ASAP7_75t_L g12037 ( 
.A(n_10564),
.B(n_8216),
.Y(n_12037)
);

INVx1_ASAP7_75t_L g12038 ( 
.A(n_10330),
.Y(n_12038)
);

OR2x2_ASAP7_75t_L g12039 ( 
.A(n_10393),
.B(n_8744),
.Y(n_12039)
);

INVx1_ASAP7_75t_L g12040 ( 
.A(n_10334),
.Y(n_12040)
);

AOI22xp33_ASAP7_75t_L g12041 ( 
.A1(n_10519),
.A2(n_8226),
.B1(n_9199),
.B2(n_8150),
.Y(n_12041)
);

INVx2_ASAP7_75t_L g12042 ( 
.A(n_10343),
.Y(n_12042)
);

BUFx12f_ASAP7_75t_L g12043 ( 
.A(n_10777),
.Y(n_12043)
);

AOI22xp33_ASAP7_75t_L g12044 ( 
.A1(n_10519),
.A2(n_8226),
.B1(n_9199),
.B2(n_8150),
.Y(n_12044)
);

INVx1_ASAP7_75t_L g12045 ( 
.A(n_10334),
.Y(n_12045)
);

NOR2x1_ASAP7_75t_SL g12046 ( 
.A(n_11000),
.B(n_8455),
.Y(n_12046)
);

BUFx2_ASAP7_75t_L g12047 ( 
.A(n_9717),
.Y(n_12047)
);

INVx1_ASAP7_75t_L g12048 ( 
.A(n_10349),
.Y(n_12048)
);

AND2x2_ASAP7_75t_L g12049 ( 
.A(n_10564),
.B(n_8216),
.Y(n_12049)
);

INVx2_ASAP7_75t_L g12050 ( 
.A(n_10344),
.Y(n_12050)
);

INVx2_ASAP7_75t_SL g12051 ( 
.A(n_9717),
.Y(n_12051)
);

INVx1_ASAP7_75t_L g12052 ( 
.A(n_10349),
.Y(n_12052)
);

AND2x2_ASAP7_75t_L g12053 ( 
.A(n_10619),
.B(n_8238),
.Y(n_12053)
);

BUFx4f_ASAP7_75t_SL g12054 ( 
.A(n_10400),
.Y(n_12054)
);

AO31x2_ASAP7_75t_L g12055 ( 
.A1(n_10535),
.A2(n_9277),
.A3(n_9500),
.B(n_9060),
.Y(n_12055)
);

AND2x2_ASAP7_75t_L g12056 ( 
.A(n_10619),
.B(n_8238),
.Y(n_12056)
);

INVx1_ASAP7_75t_L g12057 ( 
.A(n_10351),
.Y(n_12057)
);

INVx2_ASAP7_75t_SL g12058 ( 
.A(n_9736),
.Y(n_12058)
);

INVx2_ASAP7_75t_SL g12059 ( 
.A(n_9588),
.Y(n_12059)
);

AND2x2_ASAP7_75t_L g12060 ( 
.A(n_10624),
.B(n_8238),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_10351),
.Y(n_12061)
);

OAI21x1_ASAP7_75t_L g12062 ( 
.A1(n_10302),
.A2(n_8320),
.B(n_9486),
.Y(n_12062)
);

INVx1_ASAP7_75t_L g12063 ( 
.A(n_10352),
.Y(n_12063)
);

INVx4_ASAP7_75t_L g12064 ( 
.A(n_9783),
.Y(n_12064)
);

INVx3_ASAP7_75t_L g12065 ( 
.A(n_9736),
.Y(n_12065)
);

INVx1_ASAP7_75t_L g12066 ( 
.A(n_10352),
.Y(n_12066)
);

INVx1_ASAP7_75t_L g12067 ( 
.A(n_10356),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_10356),
.Y(n_12068)
);

INVx2_ASAP7_75t_L g12069 ( 
.A(n_10344),
.Y(n_12069)
);

INVx1_ASAP7_75t_L g12070 ( 
.A(n_10358),
.Y(n_12070)
);

INVx1_ASAP7_75t_L g12071 ( 
.A(n_10358),
.Y(n_12071)
);

INVxp67_ASAP7_75t_L g12072 ( 
.A(n_10641),
.Y(n_12072)
);

NAND2xp5_ASAP7_75t_L g12073 ( 
.A(n_10845),
.B(n_10901),
.Y(n_12073)
);

AND2x2_ASAP7_75t_L g12074 ( 
.A(n_10624),
.B(n_8238),
.Y(n_12074)
);

INVx2_ASAP7_75t_L g12075 ( 
.A(n_10344),
.Y(n_12075)
);

INVx2_ASAP7_75t_L g12076 ( 
.A(n_10355),
.Y(n_12076)
);

INVx2_ASAP7_75t_L g12077 ( 
.A(n_10355),
.Y(n_12077)
);

OAI21x1_ASAP7_75t_L g12078 ( 
.A1(n_10302),
.A2(n_9488),
.B(n_9486),
.Y(n_12078)
);

INVx1_ASAP7_75t_L g12079 ( 
.A(n_10360),
.Y(n_12079)
);

INVx1_ASAP7_75t_L g12080 ( 
.A(n_10360),
.Y(n_12080)
);

INVx2_ASAP7_75t_L g12081 ( 
.A(n_10355),
.Y(n_12081)
);

HB1xp67_ASAP7_75t_L g12082 ( 
.A(n_10362),
.Y(n_12082)
);

INVx1_ASAP7_75t_L g12083 ( 
.A(n_10362),
.Y(n_12083)
);

AND2x4_ASAP7_75t_L g12084 ( 
.A(n_9598),
.B(n_8455),
.Y(n_12084)
);

AOI22xp33_ASAP7_75t_L g12085 ( 
.A1(n_10521),
.A2(n_9199),
.B1(n_8150),
.B2(n_8571),
.Y(n_12085)
);

INVx1_ASAP7_75t_L g12086 ( 
.A(n_10364),
.Y(n_12086)
);

INVx1_ASAP7_75t_L g12087 ( 
.A(n_10364),
.Y(n_12087)
);

HB1xp67_ASAP7_75t_L g12088 ( 
.A(n_10367),
.Y(n_12088)
);

AOI22xp33_ASAP7_75t_L g12089 ( 
.A1(n_10521),
.A2(n_9199),
.B1(n_8150),
.B2(n_8571),
.Y(n_12089)
);

INVx2_ASAP7_75t_L g12090 ( 
.A(n_10359),
.Y(n_12090)
);

INVx1_ASAP7_75t_L g12091 ( 
.A(n_10367),
.Y(n_12091)
);

INVx1_ASAP7_75t_L g12092 ( 
.A(n_10373),
.Y(n_12092)
);

OA21x2_ASAP7_75t_L g12093 ( 
.A1(n_9840),
.A2(n_8463),
.B(n_8178),
.Y(n_12093)
);

INVx3_ASAP7_75t_L g12094 ( 
.A(n_9736),
.Y(n_12094)
);

AND2x2_ASAP7_75t_L g12095 ( 
.A(n_10672),
.B(n_10689),
.Y(n_12095)
);

HB1xp67_ASAP7_75t_L g12096 ( 
.A(n_10373),
.Y(n_12096)
);

INVx1_ASAP7_75t_L g12097 ( 
.A(n_10381),
.Y(n_12097)
);

INVx2_ASAP7_75t_L g12098 ( 
.A(n_10359),
.Y(n_12098)
);

INVx2_ASAP7_75t_L g12099 ( 
.A(n_10359),
.Y(n_12099)
);

INVx1_ASAP7_75t_L g12100 ( 
.A(n_10381),
.Y(n_12100)
);

OAI21x1_ASAP7_75t_L g12101 ( 
.A1(n_10345),
.A2(n_9488),
.B(n_9486),
.Y(n_12101)
);

INVx1_ASAP7_75t_L g12102 ( 
.A(n_10383),
.Y(n_12102)
);

BUFx2_ASAP7_75t_R g12103 ( 
.A(n_9637),
.Y(n_12103)
);

INVx2_ASAP7_75t_L g12104 ( 
.A(n_10382),
.Y(n_12104)
);

NAND2xp5_ASAP7_75t_L g12105 ( 
.A(n_10369),
.B(n_8576),
.Y(n_12105)
);

INVx2_ASAP7_75t_L g12106 ( 
.A(n_10382),
.Y(n_12106)
);

INVx2_ASAP7_75t_L g12107 ( 
.A(n_10382),
.Y(n_12107)
);

INVx1_ASAP7_75t_L g12108 ( 
.A(n_10383),
.Y(n_12108)
);

INVx1_ASAP7_75t_L g12109 ( 
.A(n_10397),
.Y(n_12109)
);

INVx2_ASAP7_75t_L g12110 ( 
.A(n_10392),
.Y(n_12110)
);

AND2x2_ASAP7_75t_L g12111 ( 
.A(n_10672),
.B(n_8238),
.Y(n_12111)
);

INVx1_ASAP7_75t_L g12112 ( 
.A(n_10397),
.Y(n_12112)
);

HB1xp67_ASAP7_75t_L g12113 ( 
.A(n_10401),
.Y(n_12113)
);

INVx1_ASAP7_75t_L g12114 ( 
.A(n_10401),
.Y(n_12114)
);

INVx2_ASAP7_75t_SL g12115 ( 
.A(n_9782),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_10408),
.Y(n_12116)
);

INVx1_ASAP7_75t_L g12117 ( 
.A(n_10408),
.Y(n_12117)
);

INVx1_ASAP7_75t_L g12118 ( 
.A(n_10411),
.Y(n_12118)
);

OAI21x1_ASAP7_75t_L g12119 ( 
.A1(n_10345),
.A2(n_9526),
.B(n_9488),
.Y(n_12119)
);

NAND2xp5_ASAP7_75t_L g12120 ( 
.A(n_10369),
.B(n_8912),
.Y(n_12120)
);

INVx2_ASAP7_75t_L g12121 ( 
.A(n_10392),
.Y(n_12121)
);

INVx1_ASAP7_75t_SL g12122 ( 
.A(n_10641),
.Y(n_12122)
);

INVx3_ASAP7_75t_L g12123 ( 
.A(n_9782),
.Y(n_12123)
);

OR2x2_ASAP7_75t_L g12124 ( 
.A(n_10402),
.B(n_8822),
.Y(n_12124)
);

AND2x2_ASAP7_75t_L g12125 ( 
.A(n_10689),
.B(n_8238),
.Y(n_12125)
);

INVx2_ASAP7_75t_L g12126 ( 
.A(n_10392),
.Y(n_12126)
);

INVx2_ASAP7_75t_L g12127 ( 
.A(n_10403),
.Y(n_12127)
);

BUFx3_ASAP7_75t_L g12128 ( 
.A(n_10645),
.Y(n_12128)
);

HB1xp67_ASAP7_75t_L g12129 ( 
.A(n_10411),
.Y(n_12129)
);

INVx1_ASAP7_75t_L g12130 ( 
.A(n_10412),
.Y(n_12130)
);

BUFx2_ASAP7_75t_L g12131 ( 
.A(n_9782),
.Y(n_12131)
);

NAND2xp5_ASAP7_75t_L g12132 ( 
.A(n_10404),
.B(n_8912),
.Y(n_12132)
);

AO21x1_ASAP7_75t_L g12133 ( 
.A1(n_10085),
.A2(n_9301),
.B(n_8930),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_10412),
.Y(n_12134)
);

INVx1_ASAP7_75t_L g12135 ( 
.A(n_10418),
.Y(n_12135)
);

INVx2_ASAP7_75t_L g12136 ( 
.A(n_10403),
.Y(n_12136)
);

OR2x2_ASAP7_75t_L g12137 ( 
.A(n_10402),
.B(n_8822),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_10418),
.Y(n_12138)
);

AND2x2_ASAP7_75t_L g12139 ( 
.A(n_10730),
.B(n_8256),
.Y(n_12139)
);

INVx2_ASAP7_75t_L g12140 ( 
.A(n_10403),
.Y(n_12140)
);

INVx2_ASAP7_75t_L g12141 ( 
.A(n_10413),
.Y(n_12141)
);

INVx1_ASAP7_75t_L g12142 ( 
.A(n_10431),
.Y(n_12142)
);

AND2x2_ASAP7_75t_L g12143 ( 
.A(n_10730),
.B(n_8256),
.Y(n_12143)
);

OR2x2_ASAP7_75t_L g12144 ( 
.A(n_10414),
.B(n_8822),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_10733),
.B(n_8256),
.Y(n_12145)
);

AOI21x1_ASAP7_75t_L g12146 ( 
.A1(n_9643),
.A2(n_9266),
.B(n_9190),
.Y(n_12146)
);

BUFx2_ASAP7_75t_L g12147 ( 
.A(n_9828),
.Y(n_12147)
);

INVx1_ASAP7_75t_L g12148 ( 
.A(n_10431),
.Y(n_12148)
);

OAI21x1_ASAP7_75t_L g12149 ( 
.A1(n_10717),
.A2(n_9528),
.B(n_9526),
.Y(n_12149)
);

INVx2_ASAP7_75t_L g12150 ( 
.A(n_10413),
.Y(n_12150)
);

INVx2_ASAP7_75t_L g12151 ( 
.A(n_10413),
.Y(n_12151)
);

OAI21xp5_ASAP7_75t_L g12152 ( 
.A1(n_10033),
.A2(n_8987),
.B(n_8971),
.Y(n_12152)
);

BUFx6f_ASAP7_75t_L g12153 ( 
.A(n_9828),
.Y(n_12153)
);

OR2x6_ASAP7_75t_L g12154 ( 
.A(n_9856),
.B(n_9060),
.Y(n_12154)
);

INVx2_ASAP7_75t_SL g12155 ( 
.A(n_9828),
.Y(n_12155)
);

INVx2_ASAP7_75t_L g12156 ( 
.A(n_10415),
.Y(n_12156)
);

AOI21x1_ASAP7_75t_L g12157 ( 
.A1(n_9643),
.A2(n_9329),
.B(n_9318),
.Y(n_12157)
);

INVx2_ASAP7_75t_L g12158 ( 
.A(n_10415),
.Y(n_12158)
);

NAND2xp5_ASAP7_75t_L g12159 ( 
.A(n_10404),
.B(n_9301),
.Y(n_12159)
);

OR2x2_ASAP7_75t_L g12160 ( 
.A(n_10414),
.B(n_8861),
.Y(n_12160)
);

BUFx4f_ASAP7_75t_L g12161 ( 
.A(n_9856),
.Y(n_12161)
);

INVx1_ASAP7_75t_L g12162 ( 
.A(n_10436),
.Y(n_12162)
);

INVx1_ASAP7_75t_L g12163 ( 
.A(n_10436),
.Y(n_12163)
);

INVx1_ASAP7_75t_L g12164 ( 
.A(n_10437),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_10437),
.Y(n_12165)
);

BUFx6f_ASAP7_75t_L g12166 ( 
.A(n_9856),
.Y(n_12166)
);

INVx2_ASAP7_75t_L g12167 ( 
.A(n_10415),
.Y(n_12167)
);

CKINVDCx20_ASAP7_75t_R g12168 ( 
.A(n_9706),
.Y(n_12168)
);

HB1xp67_ASAP7_75t_L g12169 ( 
.A(n_10443),
.Y(n_12169)
);

INVx3_ASAP7_75t_L g12170 ( 
.A(n_11014),
.Y(n_12170)
);

AOI22xp33_ASAP7_75t_L g12171 ( 
.A1(n_10521),
.A2(n_8150),
.B1(n_8571),
.B2(n_8297),
.Y(n_12171)
);

INVx1_ASAP7_75t_L g12172 ( 
.A(n_10443),
.Y(n_12172)
);

AND2x2_ASAP7_75t_L g12173 ( 
.A(n_10733),
.B(n_8256),
.Y(n_12173)
);

INVxp33_ASAP7_75t_SL g12174 ( 
.A(n_10753),
.Y(n_12174)
);

AO21x2_ASAP7_75t_L g12175 ( 
.A1(n_10004),
.A2(n_9027),
.B(n_9019),
.Y(n_12175)
);

INVx2_ASAP7_75t_SL g12176 ( 
.A(n_10233),
.Y(n_12176)
);

OAI21x1_ASAP7_75t_L g12177 ( 
.A1(n_10717),
.A2(n_9528),
.B(n_9526),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_10444),
.Y(n_12178)
);

INVx1_ASAP7_75t_L g12179 ( 
.A(n_10444),
.Y(n_12179)
);

INVx2_ASAP7_75t_L g12180 ( 
.A(n_10417),
.Y(n_12180)
);

BUFx4f_ASAP7_75t_SL g12181 ( 
.A(n_10493),
.Y(n_12181)
);

OR2x6_ASAP7_75t_L g12182 ( 
.A(n_9894),
.B(n_9060),
.Y(n_12182)
);

INVx1_ASAP7_75t_L g12183 ( 
.A(n_10451),
.Y(n_12183)
);

INVx1_ASAP7_75t_L g12184 ( 
.A(n_10451),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_10033),
.B(n_9258),
.Y(n_12185)
);

INVx1_ASAP7_75t_SL g12186 ( 
.A(n_9859),
.Y(n_12186)
);

INVx1_ASAP7_75t_L g12187 ( 
.A(n_10452),
.Y(n_12187)
);

BUFx6f_ASAP7_75t_L g12188 ( 
.A(n_9894),
.Y(n_12188)
);

INVx2_ASAP7_75t_L g12189 ( 
.A(n_10417),
.Y(n_12189)
);

BUFx2_ASAP7_75t_SL g12190 ( 
.A(n_9767),
.Y(n_12190)
);

INVx3_ASAP7_75t_L g12191 ( 
.A(n_11014),
.Y(n_12191)
);

INVx2_ASAP7_75t_L g12192 ( 
.A(n_10417),
.Y(n_12192)
);

INVx1_ASAP7_75t_L g12193 ( 
.A(n_10452),
.Y(n_12193)
);

INVx1_ASAP7_75t_L g12194 ( 
.A(n_10456),
.Y(n_12194)
);

INVx2_ASAP7_75t_L g12195 ( 
.A(n_10419),
.Y(n_12195)
);

INVx1_ASAP7_75t_L g12196 ( 
.A(n_10456),
.Y(n_12196)
);

INVxp67_ASAP7_75t_R g12197 ( 
.A(n_10933),
.Y(n_12197)
);

HB1xp67_ASAP7_75t_L g12198 ( 
.A(n_10463),
.Y(n_12198)
);

BUFx6f_ASAP7_75t_L g12199 ( 
.A(n_9894),
.Y(n_12199)
);

AO21x2_ASAP7_75t_L g12200 ( 
.A1(n_10004),
.A2(n_9019),
.B(n_8855),
.Y(n_12200)
);

INVx2_ASAP7_75t_L g12201 ( 
.A(n_10419),
.Y(n_12201)
);

OR2x2_ASAP7_75t_L g12202 ( 
.A(n_10607),
.B(n_8861),
.Y(n_12202)
);

INVx1_ASAP7_75t_L g12203 ( 
.A(n_10463),
.Y(n_12203)
);

NOR2x1_ASAP7_75t_R g12204 ( 
.A(n_9697),
.B(n_7326),
.Y(n_12204)
);

INVx2_ASAP7_75t_L g12205 ( 
.A(n_10419),
.Y(n_12205)
);

OAI22xp5_ASAP7_75t_L g12206 ( 
.A1(n_9760),
.A2(n_9076),
.B1(n_9081),
.B2(n_9037),
.Y(n_12206)
);

AOI22xp33_ASAP7_75t_L g12207 ( 
.A1(n_10536),
.A2(n_10535),
.B1(n_10562),
.B2(n_10537),
.Y(n_12207)
);

A2O1A1Ixp33_ASAP7_75t_L g12208 ( 
.A1(n_9699),
.A2(n_8873),
.B(n_8994),
.C(n_8859),
.Y(n_12208)
);

BUFx6f_ASAP7_75t_L g12209 ( 
.A(n_9894),
.Y(n_12209)
);

AND2x2_ASAP7_75t_L g12210 ( 
.A(n_10793),
.B(n_8256),
.Y(n_12210)
);

BUFx2_ASAP7_75t_L g12211 ( 
.A(n_10371),
.Y(n_12211)
);

INVx1_ASAP7_75t_L g12212 ( 
.A(n_10466),
.Y(n_12212)
);

INVx2_ASAP7_75t_L g12213 ( 
.A(n_10421),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_10466),
.Y(n_12214)
);

BUFx2_ASAP7_75t_SL g12215 ( 
.A(n_9804),
.Y(n_12215)
);

INVx1_ASAP7_75t_L g12216 ( 
.A(n_10478),
.Y(n_12216)
);

INVx1_ASAP7_75t_L g12217 ( 
.A(n_10478),
.Y(n_12217)
);

OAI21x1_ASAP7_75t_L g12218 ( 
.A1(n_10768),
.A2(n_9533),
.B(n_9528),
.Y(n_12218)
);

INVx1_ASAP7_75t_L g12219 ( 
.A(n_10480),
.Y(n_12219)
);

INVx1_ASAP7_75t_L g12220 ( 
.A(n_10480),
.Y(n_12220)
);

INVx3_ASAP7_75t_L g12221 ( 
.A(n_10011),
.Y(n_12221)
);

AOI22xp33_ASAP7_75t_L g12222 ( 
.A1(n_10535),
.A2(n_8150),
.B1(n_8571),
.B2(n_8297),
.Y(n_12222)
);

INVx2_ASAP7_75t_SL g12223 ( 
.A(n_10233),
.Y(n_12223)
);

AND2x2_ASAP7_75t_L g12224 ( 
.A(n_10793),
.B(n_8256),
.Y(n_12224)
);

INVx2_ASAP7_75t_SL g12225 ( 
.A(n_9588),
.Y(n_12225)
);

INVx1_ASAP7_75t_L g12226 ( 
.A(n_10490),
.Y(n_12226)
);

INVxp33_ASAP7_75t_L g12227 ( 
.A(n_9776),
.Y(n_12227)
);

INVx1_ASAP7_75t_L g12228 ( 
.A(n_10490),
.Y(n_12228)
);

INVx1_ASAP7_75t_L g12229 ( 
.A(n_10494),
.Y(n_12229)
);

AOI22xp33_ASAP7_75t_L g12230 ( 
.A1(n_10537),
.A2(n_8571),
.B1(n_8297),
.B2(n_8391),
.Y(n_12230)
);

INVx2_ASAP7_75t_L g12231 ( 
.A(n_10421),
.Y(n_12231)
);

INVx3_ASAP7_75t_L g12232 ( 
.A(n_10011),
.Y(n_12232)
);

INVx2_ASAP7_75t_L g12233 ( 
.A(n_10421),
.Y(n_12233)
);

INVx1_ASAP7_75t_L g12234 ( 
.A(n_10494),
.Y(n_12234)
);

NOR2xp33_ASAP7_75t_L g12235 ( 
.A(n_10357),
.B(n_9339),
.Y(n_12235)
);

BUFx3_ASAP7_75t_L g12236 ( 
.A(n_9710),
.Y(n_12236)
);

AOI22xp33_ASAP7_75t_L g12237 ( 
.A1(n_10536),
.A2(n_8571),
.B1(n_8391),
.B2(n_8991),
.Y(n_12237)
);

INVx3_ASAP7_75t_SL g12238 ( 
.A(n_10722),
.Y(n_12238)
);

INVx1_ASAP7_75t_L g12239 ( 
.A(n_10496),
.Y(n_12239)
);

INVx2_ASAP7_75t_L g12240 ( 
.A(n_10428),
.Y(n_12240)
);

OR2x2_ASAP7_75t_L g12241 ( 
.A(n_10607),
.B(n_8861),
.Y(n_12241)
);

INVx1_ASAP7_75t_SL g12242 ( 
.A(n_9859),
.Y(n_12242)
);

INVx1_ASAP7_75t_L g12243 ( 
.A(n_10496),
.Y(n_12243)
);

INVx1_ASAP7_75t_L g12244 ( 
.A(n_10499),
.Y(n_12244)
);

INVx2_ASAP7_75t_L g12245 ( 
.A(n_10428),
.Y(n_12245)
);

AOI22xp33_ASAP7_75t_SL g12246 ( 
.A1(n_10518),
.A2(n_10440),
.B1(n_10537),
.B2(n_10536),
.Y(n_12246)
);

AOI21xp5_ASAP7_75t_L g12247 ( 
.A1(n_10447),
.A2(n_9003),
.B(n_8930),
.Y(n_12247)
);

AND2x2_ASAP7_75t_L g12248 ( 
.A(n_10769),
.B(n_8317),
.Y(n_12248)
);

BUFx2_ASAP7_75t_L g12249 ( 
.A(n_10371),
.Y(n_12249)
);

AO21x2_ASAP7_75t_L g12250 ( 
.A1(n_10206),
.A2(n_8855),
.B(n_8820),
.Y(n_12250)
);

OAI21x1_ASAP7_75t_L g12251 ( 
.A1(n_10768),
.A2(n_9541),
.B(n_9533),
.Y(n_12251)
);

BUFx2_ASAP7_75t_L g12252 ( 
.A(n_10371),
.Y(n_12252)
);

INVx2_ASAP7_75t_SL g12253 ( 
.A(n_10233),
.Y(n_12253)
);

NAND2xp5_ASAP7_75t_L g12254 ( 
.A(n_10447),
.B(n_9258),
.Y(n_12254)
);

INVx2_ASAP7_75t_L g12255 ( 
.A(n_10428),
.Y(n_12255)
);

BUFx2_ASAP7_75t_L g12256 ( 
.A(n_10371),
.Y(n_12256)
);

INVx1_ASAP7_75t_L g12257 ( 
.A(n_10499),
.Y(n_12257)
);

INVx1_ASAP7_75t_L g12258 ( 
.A(n_10508),
.Y(n_12258)
);

INVx2_ASAP7_75t_L g12259 ( 
.A(n_10433),
.Y(n_12259)
);

INVx1_ASAP7_75t_L g12260 ( 
.A(n_10508),
.Y(n_12260)
);

AO21x2_ASAP7_75t_L g12261 ( 
.A1(n_10206),
.A2(n_8820),
.B(n_9154),
.Y(n_12261)
);

AND2x2_ASAP7_75t_L g12262 ( 
.A(n_11062),
.B(n_10722),
.Y(n_12262)
);

AOI22xp33_ASAP7_75t_L g12263 ( 
.A1(n_11025),
.A2(n_10518),
.B1(n_9605),
.B2(n_10001),
.Y(n_12263)
);

AOI211xp5_ASAP7_75t_L g12264 ( 
.A1(n_11025),
.A2(n_10681),
.B(n_10532),
.C(n_10747),
.Y(n_12264)
);

OR2x2_ASAP7_75t_L g12265 ( 
.A(n_11226),
.B(n_10792),
.Y(n_12265)
);

AND2x2_ASAP7_75t_L g12266 ( 
.A(n_11090),
.B(n_10754),
.Y(n_12266)
);

AOI22xp33_ASAP7_75t_SL g12267 ( 
.A1(n_11289),
.A2(n_10573),
.B1(n_10579),
.B2(n_10562),
.Y(n_12267)
);

OAI21x1_ASAP7_75t_L g12268 ( 
.A1(n_11548),
.A2(n_11819),
.B(n_11810),
.Y(n_12268)
);

CKINVDCx5p33_ASAP7_75t_R g12269 ( 
.A(n_12043),
.Y(n_12269)
);

OAI21x1_ASAP7_75t_L g12270 ( 
.A1(n_11664),
.A2(n_9616),
.B(n_9587),
.Y(n_12270)
);

INVx4_ASAP7_75t_L g12271 ( 
.A(n_12043),
.Y(n_12271)
);

INVx5_ASAP7_75t_SL g12272 ( 
.A(n_11325),
.Y(n_12272)
);

NAND2xp5_ASAP7_75t_L g12273 ( 
.A(n_11045),
.B(n_10390),
.Y(n_12273)
);

OR2x6_ASAP7_75t_L g12274 ( 
.A(n_11355),
.B(n_9894),
.Y(n_12274)
);

AND2x4_ASAP7_75t_L g12275 ( 
.A(n_11755),
.B(n_9972),
.Y(n_12275)
);

INVx1_ASAP7_75t_L g12276 ( 
.A(n_11822),
.Y(n_12276)
);

AND2x4_ASAP7_75t_L g12277 ( 
.A(n_11789),
.B(n_9972),
.Y(n_12277)
);

AOI221x1_ASAP7_75t_SL g12278 ( 
.A1(n_12004),
.A2(n_10322),
.B1(n_10747),
.B2(n_10532),
.C(n_10370),
.Y(n_12278)
);

INVx1_ASAP7_75t_L g12279 ( 
.A(n_11822),
.Y(n_12279)
);

AOI22xp33_ASAP7_75t_L g12280 ( 
.A1(n_11034),
.A2(n_9605),
.B1(n_10001),
.B2(n_10020),
.Y(n_12280)
);

OAI22xp5_ASAP7_75t_L g12281 ( 
.A1(n_11217),
.A2(n_10754),
.B1(n_9781),
.B2(n_10117),
.Y(n_12281)
);

INVx2_ASAP7_75t_L g12282 ( 
.A(n_12059),
.Y(n_12282)
);

AOI22xp33_ASAP7_75t_L g12283 ( 
.A1(n_11289),
.A2(n_9605),
.B1(n_10001),
.B2(n_10020),
.Y(n_12283)
);

AOI221xp5_ASAP7_75t_L g12284 ( 
.A1(n_11256),
.A2(n_10579),
.B1(n_10581),
.B2(n_10573),
.C(n_10562),
.Y(n_12284)
);

AOI22xp33_ASAP7_75t_L g12285 ( 
.A1(n_11590),
.A2(n_11946),
.B1(n_11962),
.B2(n_11204),
.Y(n_12285)
);

AOI22xp33_ASAP7_75t_L g12286 ( 
.A1(n_11775),
.A2(n_12021),
.B1(n_11371),
.B2(n_11541),
.Y(n_12286)
);

NAND2xp5_ASAP7_75t_L g12287 ( 
.A(n_11179),
.B(n_10567),
.Y(n_12287)
);

AOI22xp33_ASAP7_75t_L g12288 ( 
.A1(n_11541),
.A2(n_9605),
.B1(n_10001),
.B2(n_10020),
.Y(n_12288)
);

AOI211x1_ASAP7_75t_L g12289 ( 
.A1(n_11123),
.A2(n_10322),
.B(n_10370),
.C(n_10285),
.Y(n_12289)
);

AOI22xp33_ASAP7_75t_L g12290 ( 
.A1(n_12246),
.A2(n_9605),
.B1(n_10001),
.B2(n_10020),
.Y(n_12290)
);

NAND2xp5_ASAP7_75t_L g12291 ( 
.A(n_11183),
.B(n_10296),
.Y(n_12291)
);

INVx6_ASAP7_75t_L g12292 ( 
.A(n_11598),
.Y(n_12292)
);

INVx2_ASAP7_75t_SL g12293 ( 
.A(n_12128),
.Y(n_12293)
);

AOI22xp33_ASAP7_75t_L g12294 ( 
.A1(n_11882),
.A2(n_9585),
.B1(n_9615),
.B2(n_10573),
.Y(n_12294)
);

AOI222xp33_ASAP7_75t_L g12295 ( 
.A1(n_12005),
.A2(n_10579),
.B1(n_10581),
.B2(n_10587),
.C1(n_10586),
.C2(n_10585),
.Y(n_12295)
);

AOI221xp5_ASAP7_75t_L g12296 ( 
.A1(n_11256),
.A2(n_10586),
.B1(n_10587),
.B2(n_10585),
.C(n_10581),
.Y(n_12296)
);

AOI21xp5_ASAP7_75t_L g12297 ( 
.A1(n_11186),
.A2(n_11579),
.B(n_12152),
.Y(n_12297)
);

INVx2_ASAP7_75t_L g12298 ( 
.A(n_12225),
.Y(n_12298)
);

AND2x2_ASAP7_75t_L g12299 ( 
.A(n_11101),
.B(n_11135),
.Y(n_12299)
);

INVx1_ASAP7_75t_L g12300 ( 
.A(n_11896),
.Y(n_12300)
);

NAND2xp5_ASAP7_75t_L g12301 ( 
.A(n_11138),
.B(n_10296),
.Y(n_12301)
);

AOI211x1_ASAP7_75t_L g12302 ( 
.A1(n_11227),
.A2(n_10285),
.B(n_10904),
.C(n_10903),
.Y(n_12302)
);

AOI21xp33_ASAP7_75t_L g12303 ( 
.A1(n_11980),
.A2(n_11933),
.B(n_11757),
.Y(n_12303)
);

OAI211xp5_ASAP7_75t_SL g12304 ( 
.A1(n_11446),
.A2(n_11202),
.B(n_11044),
.C(n_11120),
.Y(n_12304)
);

NAND3xp33_ASAP7_75t_L g12305 ( 
.A(n_11866),
.B(n_10966),
.C(n_10085),
.Y(n_12305)
);

AOI22xp33_ASAP7_75t_SL g12306 ( 
.A1(n_11033),
.A2(n_10586),
.B1(n_10587),
.B2(n_10585),
.Y(n_12306)
);

AOI22xp33_ASAP7_75t_L g12307 ( 
.A1(n_11476),
.A2(n_10596),
.B1(n_10646),
.B2(n_10595),
.Y(n_12307)
);

AOI22xp33_ASAP7_75t_L g12308 ( 
.A1(n_11343),
.A2(n_11911),
.B1(n_11900),
.B2(n_11323),
.Y(n_12308)
);

NAND2xp5_ASAP7_75t_L g12309 ( 
.A(n_11160),
.B(n_10409),
.Y(n_12309)
);

OA21x2_ASAP7_75t_L g12310 ( 
.A1(n_11115),
.A2(n_10795),
.B(n_10781),
.Y(n_12310)
);

AOI22xp5_ASAP7_75t_L g12311 ( 
.A1(n_11033),
.A2(n_10440),
.B1(n_10811),
.B2(n_10273),
.Y(n_12311)
);

AND2x2_ASAP7_75t_L g12312 ( 
.A(n_11694),
.B(n_10321),
.Y(n_12312)
);

OAI211xp5_ASAP7_75t_L g12313 ( 
.A1(n_11980),
.A2(n_11004),
.B(n_9922),
.C(n_9822),
.Y(n_12313)
);

INVx2_ASAP7_75t_L g12314 ( 
.A(n_11599),
.Y(n_12314)
);

AND2x2_ASAP7_75t_L g12315 ( 
.A(n_11718),
.B(n_10321),
.Y(n_12315)
);

AND2x2_ASAP7_75t_L g12316 ( 
.A(n_11771),
.B(n_10258),
.Y(n_12316)
);

AOI222xp33_ASAP7_75t_L g12317 ( 
.A1(n_11858),
.A2(n_10595),
.B1(n_10596),
.B2(n_10647),
.C1(n_10646),
.C2(n_10148),
.Y(n_12317)
);

OAI22xp5_ASAP7_75t_L g12318 ( 
.A1(n_11238),
.A2(n_11329),
.B1(n_11933),
.B2(n_12247),
.Y(n_12318)
);

AOI221xp5_ASAP7_75t_L g12319 ( 
.A1(n_11713),
.A2(n_10596),
.B1(n_10647),
.B2(n_10646),
.C(n_10595),
.Y(n_12319)
);

AOI22xp33_ASAP7_75t_L g12320 ( 
.A1(n_11343),
.A2(n_10647),
.B1(n_9928),
.B2(n_10055),
.Y(n_12320)
);

NOR2xp33_ASAP7_75t_L g12321 ( 
.A(n_11637),
.B(n_9765),
.Y(n_12321)
);

OAI22xp5_ASAP7_75t_L g12322 ( 
.A1(n_11861),
.A2(n_10679),
.B1(n_10374),
.B2(n_10903),
.Y(n_12322)
);

NAND2xp5_ASAP7_75t_L g12323 ( 
.A(n_11269),
.B(n_10409),
.Y(n_12323)
);

AOI21xp5_ASAP7_75t_SL g12324 ( 
.A1(n_11115),
.A2(n_10293),
.B(n_10346),
.Y(n_12324)
);

AOI22xp33_ASAP7_75t_SL g12325 ( 
.A1(n_11757),
.A2(n_10374),
.B1(n_10695),
.B2(n_9705),
.Y(n_12325)
);

OAI22xp33_ASAP7_75t_L g12326 ( 
.A1(n_11801),
.A2(n_10679),
.B1(n_10273),
.B2(n_10811),
.Y(n_12326)
);

OR2x6_ASAP7_75t_L g12327 ( 
.A(n_11355),
.B(n_11039),
.Y(n_12327)
);

OAI22xp5_ASAP7_75t_L g12328 ( 
.A1(n_11332),
.A2(n_9897),
.B1(n_9674),
.B2(n_9705),
.Y(n_12328)
);

AOI22xp33_ASAP7_75t_L g12329 ( 
.A1(n_11323),
.A2(n_9930),
.B1(n_10003),
.B2(n_10024),
.Y(n_12329)
);

AOI22xp33_ASAP7_75t_L g12330 ( 
.A1(n_11805),
.A2(n_10024),
.B1(n_9966),
.B2(n_10288),
.Y(n_12330)
);

INVx4_ASAP7_75t_L g12331 ( 
.A(n_11355),
.Y(n_12331)
);

AOI221xp5_ASAP7_75t_L g12332 ( 
.A1(n_11713),
.A2(n_9939),
.B1(n_9968),
.B2(n_9733),
.C(n_9770),
.Y(n_12332)
);

A2O1A1Ixp33_ASAP7_75t_L g12333 ( 
.A1(n_11381),
.A2(n_9822),
.B(n_9968),
.C(n_9648),
.Y(n_12333)
);

AND2x2_ASAP7_75t_L g12334 ( 
.A(n_11778),
.B(n_11093),
.Y(n_12334)
);

INVx2_ASAP7_75t_L g12335 ( 
.A(n_11617),
.Y(n_12335)
);

OAI22xp5_ASAP7_75t_SL g12336 ( 
.A1(n_12238),
.A2(n_10357),
.B1(n_9867),
.B2(n_9997),
.Y(n_12336)
);

OAI332xp33_ASAP7_75t_L g12337 ( 
.A1(n_12105),
.A2(n_10100),
.A3(n_9939),
.B1(n_10904),
.B2(n_9840),
.B3(n_9873),
.C1(n_9870),
.C2(n_9844),
.Y(n_12337)
);

AOI22xp33_ASAP7_75t_L g12338 ( 
.A1(n_11813),
.A2(n_10288),
.B1(n_9985),
.B2(n_9937),
.Y(n_12338)
);

NAND2xp5_ASAP7_75t_L g12339 ( 
.A(n_11437),
.B(n_10426),
.Y(n_12339)
);

INVx2_ASAP7_75t_L g12340 ( 
.A(n_11623),
.Y(n_12340)
);

AOI22xp33_ASAP7_75t_L g12341 ( 
.A1(n_11856),
.A2(n_10288),
.B1(n_9638),
.B2(n_9659),
.Y(n_12341)
);

OR2x2_ASAP7_75t_L g12342 ( 
.A(n_11026),
.B(n_10792),
.Y(n_12342)
);

AND2x2_ASAP7_75t_L g12343 ( 
.A(n_11094),
.B(n_10258),
.Y(n_12343)
);

OR2x2_ASAP7_75t_L g12344 ( 
.A(n_11632),
.B(n_11636),
.Y(n_12344)
);

CKINVDCx5p33_ASAP7_75t_R g12345 ( 
.A(n_11038),
.Y(n_12345)
);

OAI22xp5_ASAP7_75t_L g12346 ( 
.A1(n_11829),
.A2(n_9897),
.B1(n_9674),
.B2(n_10204),
.Y(n_12346)
);

AOI22xp33_ASAP7_75t_L g12347 ( 
.A1(n_11826),
.A2(n_10288),
.B1(n_9692),
.B2(n_9683),
.Y(n_12347)
);

INVx1_ASAP7_75t_L g12348 ( 
.A(n_11896),
.Y(n_12348)
);

AOI22xp33_ASAP7_75t_L g12349 ( 
.A1(n_11869),
.A2(n_10288),
.B1(n_9931),
.B2(n_10068),
.Y(n_12349)
);

INVx2_ASAP7_75t_SL g12350 ( 
.A(n_12128),
.Y(n_12350)
);

OA21x2_ASAP7_75t_L g12351 ( 
.A1(n_11664),
.A2(n_10795),
.B(n_10781),
.Y(n_12351)
);

NAND2xp5_ASAP7_75t_L g12352 ( 
.A(n_11437),
.B(n_10426),
.Y(n_12352)
);

INVx2_ASAP7_75t_L g12353 ( 
.A(n_11627),
.Y(n_12353)
);

CKINVDCx5p33_ASAP7_75t_R g12354 ( 
.A(n_11038),
.Y(n_12354)
);

AOI22xp33_ASAP7_75t_L g12355 ( 
.A1(n_11783),
.A2(n_10106),
.B1(n_10727),
.B2(n_10540),
.Y(n_12355)
);

OAI211xp5_ASAP7_75t_L g12356 ( 
.A1(n_11897),
.A2(n_11004),
.B(n_10100),
.C(n_9648),
.Y(n_12356)
);

OAI221xp5_ASAP7_75t_L g12357 ( 
.A1(n_11048),
.A2(n_9748),
.B1(n_10468),
.B2(n_10461),
.C(n_10460),
.Y(n_12357)
);

AOI22xp33_ASAP7_75t_L g12358 ( 
.A1(n_11783),
.A2(n_10727),
.B1(n_10464),
.B2(n_10696),
.Y(n_12358)
);

OAI22xp33_ASAP7_75t_L g12359 ( 
.A1(n_12185),
.A2(n_10090),
.B1(n_10204),
.B2(n_10283),
.Y(n_12359)
);

INVx1_ASAP7_75t_L g12360 ( 
.A(n_11904),
.Y(n_12360)
);

AOI22xp33_ASAP7_75t_SL g12361 ( 
.A1(n_11689),
.A2(n_10695),
.B1(n_10533),
.B2(n_10332),
.Y(n_12361)
);

INVx1_ASAP7_75t_L g12362 ( 
.A(n_11904),
.Y(n_12362)
);

OAI22xp5_ASAP7_75t_L g12363 ( 
.A1(n_11642),
.A2(n_9817),
.B1(n_10090),
.B2(n_9984),
.Y(n_12363)
);

INVx6_ASAP7_75t_L g12364 ( 
.A(n_11598),
.Y(n_12364)
);

AOI222xp33_ASAP7_75t_L g12365 ( 
.A1(n_11720),
.A2(n_9898),
.B1(n_9742),
.B2(n_9660),
.C1(n_9680),
.C2(n_9730),
.Y(n_12365)
);

AND2x4_ASAP7_75t_SL g12366 ( 
.A(n_11251),
.B(n_9869),
.Y(n_12366)
);

OR2x2_ASAP7_75t_L g12367 ( 
.A(n_11715),
.B(n_10797),
.Y(n_12367)
);

AND2x2_ASAP7_75t_L g12368 ( 
.A(n_11099),
.B(n_10850),
.Y(n_12368)
);

INVx1_ASAP7_75t_L g12369 ( 
.A(n_11914),
.Y(n_12369)
);

AOI22xp33_ASAP7_75t_L g12370 ( 
.A1(n_11853),
.A2(n_11689),
.B1(n_11779),
.B2(n_11402),
.Y(n_12370)
);

OAI21xp5_ASAP7_75t_L g12371 ( 
.A1(n_11389),
.A2(n_10210),
.B(n_9817),
.Y(n_12371)
);

AOI22xp33_ASAP7_75t_L g12372 ( 
.A1(n_11779),
.A2(n_11048),
.B1(n_11848),
.B2(n_11389),
.Y(n_12372)
);

OAI22xp33_ASAP7_75t_L g12373 ( 
.A1(n_11666),
.A2(n_10283),
.B1(n_10430),
.B2(n_10464),
.Y(n_12373)
);

AND2x2_ASAP7_75t_L g12374 ( 
.A(n_11325),
.B(n_10850),
.Y(n_12374)
);

INVx6_ASAP7_75t_L g12375 ( 
.A(n_11598),
.Y(n_12375)
);

OAI221xp5_ASAP7_75t_L g12376 ( 
.A1(n_11722),
.A2(n_10617),
.B1(n_10653),
.B2(n_10491),
.C(n_9848),
.Y(n_12376)
);

AND2x2_ASAP7_75t_L g12377 ( 
.A(n_12017),
.B(n_10850),
.Y(n_12377)
);

INVx1_ASAP7_75t_L g12378 ( 
.A(n_11914),
.Y(n_12378)
);

AND2x2_ASAP7_75t_L g12379 ( 
.A(n_12017),
.B(n_10870),
.Y(n_12379)
);

AOI22xp33_ASAP7_75t_L g12380 ( 
.A1(n_11848),
.A2(n_10464),
.B1(n_10696),
.B2(n_10639),
.Y(n_12380)
);

INVx1_ASAP7_75t_L g12381 ( 
.A(n_11931),
.Y(n_12381)
);

CKINVDCx5p33_ASAP7_75t_R g12382 ( 
.A(n_11168),
.Y(n_12382)
);

OAI21x1_ASAP7_75t_L g12383 ( 
.A1(n_11955),
.A2(n_9616),
.B(n_9587),
.Y(n_12383)
);

BUFx3_ASAP7_75t_L g12384 ( 
.A(n_11251),
.Y(n_12384)
);

OAI22xp5_ASAP7_75t_L g12385 ( 
.A1(n_11642),
.A2(n_9979),
.B1(n_10860),
.B2(n_10475),
.Y(n_12385)
);

OAI211xp5_ASAP7_75t_SL g12386 ( 
.A1(n_11839),
.A2(n_10788),
.B(n_10962),
.C(n_10755),
.Y(n_12386)
);

BUFx2_ASAP7_75t_L g12387 ( 
.A(n_11486),
.Y(n_12387)
);

OAI21x1_ASAP7_75t_L g12388 ( 
.A1(n_12146),
.A2(n_9616),
.B(n_9587),
.Y(n_12388)
);

NAND3xp33_ASAP7_75t_L g12389 ( 
.A(n_11839),
.B(n_9644),
.C(n_10533),
.Y(n_12389)
);

NAND2xp5_ASAP7_75t_L g12390 ( 
.A(n_11443),
.B(n_10483),
.Y(n_12390)
);

OAI211xp5_ASAP7_75t_L g12391 ( 
.A1(n_11897),
.A2(n_10533),
.B(n_9644),
.C(n_9844),
.Y(n_12391)
);

OAI211xp5_ASAP7_75t_L g12392 ( 
.A1(n_11394),
.A2(n_10533),
.B(n_9844),
.C(n_9861),
.Y(n_12392)
);

NAND3xp33_ASAP7_75t_L g12393 ( 
.A(n_11147),
.B(n_10735),
.C(n_10448),
.Y(n_12393)
);

OAI22xp5_ASAP7_75t_L g12394 ( 
.A1(n_12031),
.A2(n_10860),
.B1(n_10208),
.B2(n_10481),
.Y(n_12394)
);

OAI22xp5_ASAP7_75t_L g12395 ( 
.A1(n_11745),
.A2(n_10208),
.B1(n_10481),
.B2(n_10475),
.Y(n_12395)
);

AOI221xp5_ASAP7_75t_L g12396 ( 
.A1(n_11722),
.A2(n_10450),
.B1(n_10462),
.B2(n_10446),
.C(n_10433),
.Y(n_12396)
);

INVx2_ASAP7_75t_SL g12397 ( 
.A(n_11168),
.Y(n_12397)
);

OAI221xp5_ASAP7_75t_L g12398 ( 
.A1(n_11613),
.A2(n_9720),
.B1(n_9814),
.B2(n_9813),
.C(n_10862),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_11714),
.A2(n_10464),
.B1(n_10639),
.B2(n_9883),
.Y(n_12399)
);

AND2x2_ASAP7_75t_L g12400 ( 
.A(n_12235),
.B(n_10870),
.Y(n_12400)
);

AOI22xp33_ASAP7_75t_L g12401 ( 
.A1(n_11714),
.A2(n_10464),
.B1(n_9898),
.B2(n_10250),
.Y(n_12401)
);

INVx2_ASAP7_75t_SL g12402 ( 
.A(n_11333),
.Y(n_12402)
);

AO31x2_ASAP7_75t_L g12403 ( 
.A1(n_11218),
.A2(n_10795),
.A3(n_10824),
.B(n_10781),
.Y(n_12403)
);

AOI22xp33_ASAP7_75t_L g12404 ( 
.A1(n_11146),
.A2(n_11297),
.B1(n_11326),
.B2(n_11199),
.Y(n_12404)
);

OAI21xp33_ASAP7_75t_L g12405 ( 
.A1(n_11711),
.A2(n_10782),
.B(n_9967),
.Y(n_12405)
);

AOI21xp33_ASAP7_75t_L g12406 ( 
.A1(n_11146),
.A2(n_10221),
.B(n_9235),
.Y(n_12406)
);

AO21x2_ASAP7_75t_L g12407 ( 
.A1(n_12133),
.A2(n_10210),
.B(n_10824),
.Y(n_12407)
);

OAI22xp5_ASAP7_75t_L g12408 ( 
.A1(n_11711),
.A2(n_10208),
.B1(n_10481),
.B2(n_10475),
.Y(n_12408)
);

AOI22xp33_ASAP7_75t_L g12409 ( 
.A1(n_11354),
.A2(n_10231),
.B1(n_10839),
.B2(n_10764),
.Y(n_12409)
);

AOI222xp33_ASAP7_75t_L g12410 ( 
.A1(n_11613),
.A2(n_9742),
.B1(n_10008),
.B2(n_10450),
.C1(n_10446),
.C2(n_10433),
.Y(n_12410)
);

INVx5_ASAP7_75t_L g12411 ( 
.A(n_11039),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_11931),
.Y(n_12412)
);

OAI211xp5_ASAP7_75t_L g12413 ( 
.A1(n_11443),
.A2(n_9861),
.B(n_9870),
.C(n_9840),
.Y(n_12413)
);

OAI22xp5_ASAP7_75t_L g12414 ( 
.A1(n_11750),
.A2(n_10430),
.B1(n_9993),
.B2(n_10556),
.Y(n_12414)
);

AOI221xp5_ASAP7_75t_L g12415 ( 
.A1(n_11203),
.A2(n_10462),
.B1(n_10472),
.B2(n_10450),
.C(n_10446),
.Y(n_12415)
);

OAI21xp33_ASAP7_75t_L g12416 ( 
.A1(n_12254),
.A2(n_10782),
.B(n_9967),
.Y(n_12416)
);

INVx4_ASAP7_75t_L g12417 ( 
.A(n_11519),
.Y(n_12417)
);

INVx1_ASAP7_75t_L g12418 ( 
.A(n_11943),
.Y(n_12418)
);

NAND2xp5_ASAP7_75t_L g12419 ( 
.A(n_11453),
.B(n_10483),
.Y(n_12419)
);

NOR2xp33_ASAP7_75t_L g12420 ( 
.A(n_11637),
.B(n_12174),
.Y(n_12420)
);

OAI221xp5_ASAP7_75t_L g12421 ( 
.A1(n_11890),
.A2(n_10934),
.B1(n_10911),
.B2(n_10608),
.C(n_10604),
.Y(n_12421)
);

AND2x2_ASAP7_75t_L g12422 ( 
.A(n_12235),
.B(n_10870),
.Y(n_12422)
);

AOI21xp5_ASAP7_75t_L g12423 ( 
.A1(n_11890),
.A2(n_10837),
.B(n_10427),
.Y(n_12423)
);

AO22x1_ASAP7_75t_L g12424 ( 
.A1(n_11790),
.A2(n_10448),
.B1(n_10735),
.B2(n_10847),
.Y(n_12424)
);

NOR2xp33_ASAP7_75t_SL g12425 ( 
.A(n_12103),
.B(n_9765),
.Y(n_12425)
);

CKINVDCx20_ASAP7_75t_R g12426 ( 
.A(n_11982),
.Y(n_12426)
);

AOI22xp5_ASAP7_75t_L g12427 ( 
.A1(n_11704),
.A2(n_9995),
.B1(n_10158),
.B2(n_10786),
.Y(n_12427)
);

AOI22xp33_ASAP7_75t_L g12428 ( 
.A1(n_11203),
.A2(n_10764),
.B1(n_10839),
.B2(n_10105),
.Y(n_12428)
);

AOI22xp33_ASAP7_75t_L g12429 ( 
.A1(n_11254),
.A2(n_10126),
.B1(n_9874),
.B2(n_10275),
.Y(n_12429)
);

AOI222xp33_ASAP7_75t_L g12430 ( 
.A1(n_11254),
.A2(n_10472),
.B1(n_10484),
.B2(n_10462),
.C1(n_9861),
.C2(n_9870),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_11943),
.Y(n_12431)
);

INVx1_ASAP7_75t_L g12432 ( 
.A(n_11949),
.Y(n_12432)
);

INVx1_ASAP7_75t_SL g12433 ( 
.A(n_12054),
.Y(n_12433)
);

OAI211xp5_ASAP7_75t_L g12434 ( 
.A1(n_11453),
.A2(n_9875),
.B(n_9895),
.C(n_9873),
.Y(n_12434)
);

AND2x2_ASAP7_75t_L g12435 ( 
.A(n_11816),
.B(n_10948),
.Y(n_12435)
);

AOI222xp33_ASAP7_75t_L g12436 ( 
.A1(n_11556),
.A2(n_10484),
.B1(n_10472),
.B2(n_9873),
.C1(n_9875),
.C2(n_9895),
.Y(n_12436)
);

INVx2_ASAP7_75t_L g12437 ( 
.A(n_11638),
.Y(n_12437)
);

AOI211xp5_ASAP7_75t_L g12438 ( 
.A1(n_11245),
.A2(n_9895),
.B(n_9875),
.C(n_9993),
.Y(n_12438)
);

AOI22xp33_ASAP7_75t_SL g12439 ( 
.A1(n_11376),
.A2(n_10378),
.B1(n_10332),
.B2(n_10394),
.Y(n_12439)
);

AOI21xp33_ASAP7_75t_L g12440 ( 
.A1(n_11803),
.A2(n_10221),
.B(n_10332),
.Y(n_12440)
);

AOI22xp5_ASAP7_75t_L g12441 ( 
.A1(n_11606),
.A2(n_10467),
.B1(n_10780),
.B2(n_10842),
.Y(n_12441)
);

INVx11_ASAP7_75t_L g12442 ( 
.A(n_12054),
.Y(n_12442)
);

INVx1_ASAP7_75t_L g12443 ( 
.A(n_11949),
.Y(n_12443)
);

AOI21xp33_ASAP7_75t_L g12444 ( 
.A1(n_11046),
.A2(n_10221),
.B(n_10332),
.Y(n_12444)
);

OAI22xp5_ASAP7_75t_L g12445 ( 
.A1(n_11750),
.A2(n_10556),
.B1(n_9913),
.B2(n_9925),
.Y(n_12445)
);

NOR2xp33_ASAP7_75t_L g12446 ( 
.A(n_12174),
.B(n_10113),
.Y(n_12446)
);

OR2x2_ASAP7_75t_L g12447 ( 
.A(n_11129),
.B(n_10797),
.Y(n_12447)
);

OAI221xp5_ASAP7_75t_L g12448 ( 
.A1(n_11379),
.A2(n_11556),
.B1(n_11705),
.B2(n_12208),
.C(n_11948),
.Y(n_12448)
);

OR2x2_ASAP7_75t_L g12449 ( 
.A(n_11148),
.B(n_10807),
.Y(n_12449)
);

CKINVDCx5p33_ASAP7_75t_R g12450 ( 
.A(n_11333),
.Y(n_12450)
);

INVx1_ASAP7_75t_L g12451 ( 
.A(n_11981),
.Y(n_12451)
);

NOR2xp33_ASAP7_75t_L g12452 ( 
.A(n_11331),
.B(n_10113),
.Y(n_12452)
);

AND2x2_ASAP7_75t_L g12453 ( 
.A(n_11844),
.B(n_10948),
.Y(n_12453)
);

AND2x2_ASAP7_75t_L g12454 ( 
.A(n_11847),
.B(n_10948),
.Y(n_12454)
);

AOI221xp5_ASAP7_75t_L g12455 ( 
.A1(n_11379),
.A2(n_11705),
.B1(n_12237),
.B2(n_12230),
.C(n_12089),
.Y(n_12455)
);

AOI22xp5_ASAP7_75t_L g12456 ( 
.A1(n_11346),
.A2(n_10363),
.B1(n_10640),
.B2(n_10378),
.Y(n_12456)
);

AND2x2_ASAP7_75t_L g12457 ( 
.A(n_11873),
.B(n_9842),
.Y(n_12457)
);

AOI31xp33_ASAP7_75t_L g12458 ( 
.A1(n_11486),
.A2(n_10453),
.A3(n_10346),
.B(n_9891),
.Y(n_12458)
);

AOI221xp5_ASAP7_75t_L g12459 ( 
.A1(n_12237),
.A2(n_10484),
.B1(n_9983),
.B2(n_10135),
.C(n_10097),
.Y(n_12459)
);

INVx8_ASAP7_75t_L g12460 ( 
.A(n_11039),
.Y(n_12460)
);

AOI22xp33_ASAP7_75t_SL g12461 ( 
.A1(n_11760),
.A2(n_10378),
.B1(n_10394),
.B2(n_8621),
.Y(n_12461)
);

OAI211xp5_ASAP7_75t_L g12462 ( 
.A1(n_11461),
.A2(n_10221),
.B(n_10110),
.C(n_9616),
.Y(n_12462)
);

BUFx2_ASAP7_75t_L g12463 ( 
.A(n_12072),
.Y(n_12463)
);

AOI22xp33_ASAP7_75t_L g12464 ( 
.A1(n_11305),
.A2(n_10281),
.B1(n_10378),
.B2(n_9560),
.Y(n_12464)
);

OAI22xp5_ASAP7_75t_L g12465 ( 
.A1(n_12206),
.A2(n_10556),
.B1(n_9913),
.B2(n_9925),
.Y(n_12465)
);

HB1xp67_ASAP7_75t_L g12466 ( 
.A(n_11468),
.Y(n_12466)
);

CKINVDCx5p33_ASAP7_75t_R g12467 ( 
.A(n_11524),
.Y(n_12467)
);

AND2x2_ASAP7_75t_L g12468 ( 
.A(n_11907),
.B(n_9842),
.Y(n_12468)
);

OAI22xp5_ASAP7_75t_L g12469 ( 
.A1(n_11948),
.A2(n_12208),
.B1(n_11781),
.B2(n_11635),
.Y(n_12469)
);

AO221x2_ASAP7_75t_L g12470 ( 
.A1(n_12120),
.A2(n_10837),
.B1(n_7669),
.B2(n_8918),
.C(n_9013),
.Y(n_12470)
);

OA21x2_ASAP7_75t_L g12471 ( 
.A1(n_11831),
.A2(n_10826),
.B(n_10824),
.Y(n_12471)
);

AOI22xp33_ASAP7_75t_L g12472 ( 
.A1(n_11546),
.A2(n_9560),
.B1(n_10071),
.B2(n_10069),
.Y(n_12472)
);

INVx1_ASAP7_75t_L g12473 ( 
.A(n_11981),
.Y(n_12473)
);

OAI22xp5_ASAP7_75t_L g12474 ( 
.A1(n_11086),
.A2(n_9913),
.B1(n_9925),
.B2(n_9798),
.Y(n_12474)
);

AOI33xp33_ASAP7_75t_L g12475 ( 
.A1(n_12230),
.A2(n_10728),
.A3(n_10553),
.B1(n_10744),
.B2(n_10658),
.B3(n_10548),
.Y(n_12475)
);

INVx1_ASAP7_75t_SL g12476 ( 
.A(n_11395),
.Y(n_12476)
);

INVx2_ASAP7_75t_SL g12477 ( 
.A(n_11524),
.Y(n_12477)
);

OAI22xp5_ASAP7_75t_L g12478 ( 
.A1(n_11121),
.A2(n_9988),
.B1(n_10037),
.B2(n_9798),
.Y(n_12478)
);

AOI22xp33_ASAP7_75t_L g12479 ( 
.A1(n_11046),
.A2(n_11124),
.B1(n_11703),
.B2(n_11221),
.Y(n_12479)
);

AND2x2_ASAP7_75t_L g12480 ( 
.A(n_11457),
.B(n_9849),
.Y(n_12480)
);

NAND3xp33_ASAP7_75t_L g12481 ( 
.A(n_11461),
.B(n_10735),
.C(n_10448),
.Y(n_12481)
);

AOI21xp5_ASAP7_75t_L g12482 ( 
.A1(n_11480),
.A2(n_9973),
.B(n_9986),
.Y(n_12482)
);

INVx3_ASAP7_75t_L g12483 ( 
.A(n_11491),
.Y(n_12483)
);

A2O1A1Ixp33_ASAP7_75t_L g12484 ( 
.A1(n_11082),
.A2(n_10134),
.B(n_10167),
.C(n_10131),
.Y(n_12484)
);

OAI221xp5_ASAP7_75t_L g12485 ( 
.A1(n_12041),
.A2(n_10603),
.B1(n_10294),
.B2(n_10300),
.C(n_10299),
.Y(n_12485)
);

INVx1_ASAP7_75t_L g12486 ( 
.A(n_12082),
.Y(n_12486)
);

INVx1_ASAP7_75t_L g12487 ( 
.A(n_12082),
.Y(n_12487)
);

AOI22xp33_ASAP7_75t_L g12488 ( 
.A1(n_11124),
.A2(n_9560),
.B1(n_9775),
.B2(n_9771),
.Y(n_12488)
);

AOI22xp33_ASAP7_75t_L g12489 ( 
.A1(n_11218),
.A2(n_9560),
.B1(n_10265),
.B2(n_10394),
.Y(n_12489)
);

OR2x2_ASAP7_75t_L g12490 ( 
.A(n_11173),
.B(n_10807),
.Y(n_12490)
);

AOI22xp33_ASAP7_75t_L g12491 ( 
.A1(n_11221),
.A2(n_9560),
.B1(n_10394),
.B2(n_10181),
.Y(n_12491)
);

OAI33xp33_ASAP7_75t_L g12492 ( 
.A1(n_12132),
.A2(n_9973),
.A3(n_9986),
.B1(n_9013),
.B2(n_8918),
.B3(n_8974),
.Y(n_12492)
);

AOI22xp33_ASAP7_75t_L g12493 ( 
.A1(n_11225),
.A2(n_9871),
.B1(n_10895),
.B2(n_10479),
.Y(n_12493)
);

AOI22xp33_ASAP7_75t_SL g12494 ( 
.A1(n_12046),
.A2(n_8621),
.B1(n_8640),
.B2(n_10832),
.Y(n_12494)
);

NAND2xp5_ASAP7_75t_L g12495 ( 
.A(n_11407),
.B(n_10548),
.Y(n_12495)
);

BUFx12f_ASAP7_75t_L g12496 ( 
.A(n_11655),
.Y(n_12496)
);

INVx6_ASAP7_75t_L g12497 ( 
.A(n_11054),
.Y(n_12497)
);

OAI211xp5_ASAP7_75t_SL g12498 ( 
.A1(n_12222),
.A2(n_10788),
.B(n_10962),
.C(n_10755),
.Y(n_12498)
);

BUFx6f_ASAP7_75t_L g12499 ( 
.A(n_11039),
.Y(n_12499)
);

OAI211xp5_ASAP7_75t_L g12500 ( 
.A1(n_11287),
.A2(n_10110),
.B(n_9587),
.C(n_10298),
.Y(n_12500)
);

AOI22xp33_ASAP7_75t_L g12501 ( 
.A1(n_11225),
.A2(n_9871),
.B1(n_10623),
.B2(n_9159),
.Y(n_12501)
);

INVx1_ASAP7_75t_L g12502 ( 
.A(n_12088),
.Y(n_12502)
);

AOI22xp5_ASAP7_75t_L g12503 ( 
.A1(n_11346),
.A2(n_11868),
.B1(n_11922),
.B2(n_11842),
.Y(n_12503)
);

AOI22xp33_ASAP7_75t_L g12504 ( 
.A1(n_11248),
.A2(n_9871),
.B1(n_9159),
.B2(n_9024),
.Y(n_12504)
);

OAI22xp33_ASAP7_75t_L g12505 ( 
.A1(n_11665),
.A2(n_10449),
.B1(n_8488),
.B2(n_8481),
.Y(n_12505)
);

OAI22xp5_ASAP7_75t_L g12506 ( 
.A1(n_12041),
.A2(n_9988),
.B1(n_10037),
.B2(n_9798),
.Y(n_12506)
);

AND2x4_ASAP7_75t_L g12507 ( 
.A(n_11087),
.B(n_9972),
.Y(n_12507)
);

INVx1_ASAP7_75t_L g12508 ( 
.A(n_12088),
.Y(n_12508)
);

AOI221xp5_ASAP7_75t_L g12509 ( 
.A1(n_12085),
.A2(n_10165),
.B1(n_10197),
.B2(n_10196),
.C(n_10046),
.Y(n_12509)
);

INVx1_ASAP7_75t_SL g12510 ( 
.A(n_12181),
.Y(n_12510)
);

OAI221xp5_ASAP7_75t_SL g12511 ( 
.A1(n_12044),
.A2(n_9864),
.B1(n_10848),
.B2(n_10836),
.C(n_10832),
.Y(n_12511)
);

OAI21xp33_ASAP7_75t_L g12512 ( 
.A1(n_12159),
.A2(n_10154),
.B(n_10114),
.Y(n_12512)
);

AOI221xp5_ASAP7_75t_L g12513 ( 
.A1(n_12085),
.A2(n_10225),
.B1(n_10340),
.B2(n_10295),
.C(n_10223),
.Y(n_12513)
);

OAI22xp5_ASAP7_75t_L g12514 ( 
.A1(n_12044),
.A2(n_10037),
.B1(n_9988),
.B2(n_10180),
.Y(n_12514)
);

AND2x4_ASAP7_75t_L g12515 ( 
.A(n_11493),
.B(n_9990),
.Y(n_12515)
);

NAND2xp5_ASAP7_75t_L g12516 ( 
.A(n_11407),
.B(n_10553),
.Y(n_12516)
);

INVx2_ASAP7_75t_L g12517 ( 
.A(n_11688),
.Y(n_12517)
);

OAI22xp5_ASAP7_75t_L g12518 ( 
.A1(n_12171),
.A2(n_10219),
.B1(n_10180),
.B2(n_10174),
.Y(n_12518)
);

AOI21xp5_ASAP7_75t_L g12519 ( 
.A1(n_11746),
.A2(n_10912),
.B(n_10820),
.Y(n_12519)
);

AOI22xp33_ASAP7_75t_SL g12520 ( 
.A1(n_11842),
.A2(n_8621),
.B1(n_8640),
.B2(n_10832),
.Y(n_12520)
);

AOI22xp33_ASAP7_75t_L g12521 ( 
.A1(n_11248),
.A2(n_9871),
.B1(n_9024),
.B2(n_9794),
.Y(n_12521)
);

AOI22xp5_ASAP7_75t_L g12522 ( 
.A1(n_11868),
.A2(n_11922),
.B1(n_11501),
.B2(n_12250),
.Y(n_12522)
);

BUFx3_ASAP7_75t_L g12523 ( 
.A(n_11982),
.Y(n_12523)
);

OAI21xp5_ASAP7_75t_L g12524 ( 
.A1(n_11276),
.A2(n_8528),
.B(n_8534),
.Y(n_12524)
);

AOI22xp33_ASAP7_75t_L g12525 ( 
.A1(n_11501),
.A2(n_10248),
.B1(n_10991),
.B2(n_8391),
.Y(n_12525)
);

INVx1_ASAP7_75t_L g12526 ( 
.A(n_12096),
.Y(n_12526)
);

AOI33xp33_ASAP7_75t_L g12527 ( 
.A1(n_12171),
.A2(n_10876),
.A3(n_10728),
.B1(n_10970),
.B2(n_10744),
.B3(n_10658),
.Y(n_12527)
);

INVx2_ASAP7_75t_SL g12528 ( 
.A(n_11655),
.Y(n_12528)
);

INVx4_ASAP7_75t_L g12529 ( 
.A(n_11519),
.Y(n_12529)
);

AND2x2_ASAP7_75t_L g12530 ( 
.A(n_11458),
.B(n_9849),
.Y(n_12530)
);

CKINVDCx5p33_ASAP7_75t_R g12531 ( 
.A(n_11656),
.Y(n_12531)
);

AOI22xp33_ASAP7_75t_L g12532 ( 
.A1(n_11069),
.A2(n_8391),
.B1(n_9503),
.B2(n_10836),
.Y(n_12532)
);

AOI222xp33_ASAP7_75t_L g12533 ( 
.A1(n_11862),
.A2(n_10470),
.B1(n_10384),
.B2(n_10505),
.C1(n_10435),
.C2(n_10354),
.Y(n_12533)
);

AOI22xp33_ASAP7_75t_SL g12534 ( 
.A1(n_11743),
.A2(n_8640),
.B1(n_10848),
.B2(n_10836),
.Y(n_12534)
);

AND2x2_ASAP7_75t_L g12535 ( 
.A(n_11471),
.B(n_9853),
.Y(n_12535)
);

O2A1O1Ixp33_ASAP7_75t_L g12536 ( 
.A1(n_11412),
.A2(n_10515),
.B(n_10563),
.C(n_10513),
.Y(n_12536)
);

INVx1_ASAP7_75t_L g12537 ( 
.A(n_12096),
.Y(n_12537)
);

OA21x2_ASAP7_75t_L g12538 ( 
.A1(n_11753),
.A2(n_10827),
.B(n_10826),
.Y(n_12538)
);

INVx1_ASAP7_75t_L g12539 ( 
.A(n_12113),
.Y(n_12539)
);

INVx1_ASAP7_75t_L g12540 ( 
.A(n_12113),
.Y(n_12540)
);

AOI22xp33_ASAP7_75t_SL g12541 ( 
.A1(n_12250),
.A2(n_10869),
.B1(n_10880),
.B2(n_10848),
.Y(n_12541)
);

AOI22xp33_ASAP7_75t_L g12542 ( 
.A1(n_11069),
.A2(n_8391),
.B1(n_9503),
.B2(n_10869),
.Y(n_12542)
);

AOI221xp5_ASAP7_75t_L g12543 ( 
.A1(n_12089),
.A2(n_10654),
.B1(n_10670),
.B2(n_10626),
.C(n_10612),
.Y(n_12543)
);

OAI221xp5_ASAP7_75t_L g12544 ( 
.A1(n_12222),
.A2(n_10818),
.B1(n_10825),
.B2(n_10816),
.C(n_10800),
.Y(n_12544)
);

AND2x4_ASAP7_75t_L g12545 ( 
.A(n_11644),
.B(n_9990),
.Y(n_12545)
);

OR2x2_ASAP7_75t_L g12546 ( 
.A(n_11416),
.B(n_10114),
.Y(n_12546)
);

AOI22xp33_ASAP7_75t_SL g12547 ( 
.A1(n_12261),
.A2(n_10869),
.B1(n_10884),
.B2(n_10880),
.Y(n_12547)
);

AOI22xp33_ASAP7_75t_L g12548 ( 
.A1(n_11069),
.A2(n_9503),
.B1(n_10884),
.B2(n_10880),
.Y(n_12548)
);

BUFx4f_ASAP7_75t_SL g12549 ( 
.A(n_12168),
.Y(n_12549)
);

HB1xp67_ASAP7_75t_L g12550 ( 
.A(n_11468),
.Y(n_12550)
);

AOI22xp33_ASAP7_75t_L g12551 ( 
.A1(n_11070),
.A2(n_9503),
.B1(n_10887),
.B2(n_10884),
.Y(n_12551)
);

INVx1_ASAP7_75t_L g12552 ( 
.A(n_12129),
.Y(n_12552)
);

AOI22xp33_ASAP7_75t_L g12553 ( 
.A1(n_11070),
.A2(n_9503),
.B1(n_10888),
.B2(n_10887),
.Y(n_12553)
);

AND2x2_ASAP7_75t_L g12554 ( 
.A(n_11472),
.B(n_9853),
.Y(n_12554)
);

AOI221xp5_ASAP7_75t_L g12555 ( 
.A1(n_11231),
.A2(n_10703),
.B1(n_10888),
.B2(n_10920),
.C(n_10887),
.Y(n_12555)
);

OAI22xp33_ASAP7_75t_L g12556 ( 
.A1(n_11672),
.A2(n_10449),
.B1(n_8488),
.B2(n_8481),
.Y(n_12556)
);

INVx1_ASAP7_75t_L g12557 ( 
.A(n_12129),
.Y(n_12557)
);

AND2x4_ASAP7_75t_L g12558 ( 
.A(n_11686),
.B(n_9990),
.Y(n_12558)
);

AOI22xp33_ASAP7_75t_L g12559 ( 
.A1(n_11070),
.A2(n_10920),
.B1(n_10888),
.B2(n_10549),
.Y(n_12559)
);

INVx2_ASAP7_75t_L g12560 ( 
.A(n_11477),
.Y(n_12560)
);

AND2x2_ASAP7_75t_L g12561 ( 
.A(n_11507),
.B(n_11512),
.Y(n_12561)
);

AOI22xp33_ASAP7_75t_L g12562 ( 
.A1(n_12261),
.A2(n_10920),
.B1(n_10488),
.B2(n_10599),
.Y(n_12562)
);

OAI211xp5_ASAP7_75t_L g12563 ( 
.A1(n_11181),
.A2(n_10110),
.B(n_10304),
.C(n_10298),
.Y(n_12563)
);

AOI22xp33_ASAP7_75t_L g12564 ( 
.A1(n_11542),
.A2(n_10574),
.B1(n_9810),
.B2(n_9726),
.Y(n_12564)
);

INVx1_ASAP7_75t_L g12565 ( 
.A(n_12169),
.Y(n_12565)
);

OAI22xp5_ASAP7_75t_L g12566 ( 
.A1(n_11077),
.A2(n_10219),
.B1(n_10174),
.B2(n_10161),
.Y(n_12566)
);

AOI22xp33_ASAP7_75t_L g12567 ( 
.A1(n_11542),
.A2(n_9810),
.B1(n_9726),
.B2(n_8991),
.Y(n_12567)
);

AO21x2_ASAP7_75t_L g12568 ( 
.A1(n_11281),
.A2(n_10827),
.B(n_10826),
.Y(n_12568)
);

CKINVDCx11_ASAP7_75t_R g12569 ( 
.A(n_11582),
.Y(n_12569)
);

INVx2_ASAP7_75t_SL g12570 ( 
.A(n_11656),
.Y(n_12570)
);

A2O1A1Ixp33_ASAP7_75t_L g12571 ( 
.A1(n_11276),
.A2(n_8488),
.B(n_8481),
.C(n_10237),
.Y(n_12571)
);

AOI22xp33_ASAP7_75t_L g12572 ( 
.A1(n_11031),
.A2(n_9810),
.B1(n_9726),
.B2(n_8991),
.Y(n_12572)
);

NAND3xp33_ASAP7_75t_L g12573 ( 
.A(n_11031),
.B(n_10735),
.C(n_10448),
.Y(n_12573)
);

AOI22xp33_ASAP7_75t_L g12574 ( 
.A1(n_11031),
.A2(n_9810),
.B1(n_9726),
.B2(n_8991),
.Y(n_12574)
);

INVx1_ASAP7_75t_L g12575 ( 
.A(n_12169),
.Y(n_12575)
);

INVx1_ASAP7_75t_L g12576 ( 
.A(n_12198),
.Y(n_12576)
);

INVx1_ASAP7_75t_L g12577 ( 
.A(n_12198),
.Y(n_12577)
);

OAI22xp5_ASAP7_75t_L g12578 ( 
.A1(n_11083),
.A2(n_10174),
.B1(n_10161),
.B2(n_8586),
.Y(n_12578)
);

NAND2xp5_ASAP7_75t_L g12579 ( 
.A(n_11412),
.B(n_10876),
.Y(n_12579)
);

OAI22xp5_ASAP7_75t_L g12580 ( 
.A1(n_11791),
.A2(n_10161),
.B1(n_8586),
.B2(n_8632),
.Y(n_12580)
);

INVx2_ASAP7_75t_L g12581 ( 
.A(n_11550),
.Y(n_12581)
);

AOI22xp5_ASAP7_75t_L g12582 ( 
.A1(n_11640),
.A2(n_8668),
.B1(n_8913),
.B2(n_10284),
.Y(n_12582)
);

INVx2_ASAP7_75t_L g12583 ( 
.A(n_11570),
.Y(n_12583)
);

AND2x2_ASAP7_75t_L g12584 ( 
.A(n_11283),
.B(n_10232),
.Y(n_12584)
);

INVx2_ASAP7_75t_L g12585 ( 
.A(n_11050),
.Y(n_12585)
);

OR2x2_ASAP7_75t_L g12586 ( 
.A(n_11999),
.B(n_10154),
.Y(n_12586)
);

BUFx2_ASAP7_75t_L g12587 ( 
.A(n_11974),
.Y(n_12587)
);

AND2x2_ASAP7_75t_L g12588 ( 
.A(n_11283),
.B(n_10232),
.Y(n_12588)
);

AOI22xp33_ASAP7_75t_L g12589 ( 
.A1(n_11983),
.A2(n_8991),
.B1(n_9015),
.B2(n_9005),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_11406),
.Y(n_12590)
);

AOI22xp33_ASAP7_75t_L g12591 ( 
.A1(n_11983),
.A2(n_9005),
.B1(n_9015),
.B2(n_10973),
.Y(n_12591)
);

AND2x2_ASAP7_75t_L g12592 ( 
.A(n_11438),
.B(n_10858),
.Y(n_12592)
);

BUFx4f_ASAP7_75t_L g12593 ( 
.A(n_11041),
.Y(n_12593)
);

BUFx6f_ASAP7_75t_L g12594 ( 
.A(n_11041),
.Y(n_12594)
);

OAI22xp5_ASAP7_75t_L g12595 ( 
.A1(n_11408),
.A2(n_8586),
.B1(n_8632),
.B2(n_8468),
.Y(n_12595)
);

AND2x4_ASAP7_75t_L g12596 ( 
.A(n_11794),
.B(n_10009),
.Y(n_12596)
);

NOR3xp33_ASAP7_75t_L g12597 ( 
.A(n_11794),
.B(n_10095),
.C(n_9601),
.Y(n_12597)
);

AOI22xp5_ASAP7_75t_L g12598 ( 
.A1(n_11640),
.A2(n_8668),
.B1(n_8913),
.B2(n_8716),
.Y(n_12598)
);

OAI22xp5_ASAP7_75t_L g12599 ( 
.A1(n_11442),
.A2(n_8632),
.B1(n_8468),
.B2(n_8974),
.Y(n_12599)
);

INVx1_ASAP7_75t_L g12600 ( 
.A(n_11406),
.Y(n_12600)
);

OAI22xp33_ASAP7_75t_L g12601 ( 
.A1(n_11231),
.A2(n_10449),
.B1(n_8488),
.B2(n_8481),
.Y(n_12601)
);

AOI22xp33_ASAP7_75t_L g12602 ( 
.A1(n_11081),
.A2(n_12012),
.B1(n_11284),
.B2(n_11339),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_11800),
.Y(n_12603)
);

AOI22xp33_ASAP7_75t_L g12604 ( 
.A1(n_11081),
.A2(n_9005),
.B1(n_9015),
.B2(n_8322),
.Y(n_12604)
);

AOI22xp33_ASAP7_75t_L g12605 ( 
.A1(n_11081),
.A2(n_9005),
.B1(n_9015),
.B2(n_8322),
.Y(n_12605)
);

NAND2xp5_ASAP7_75t_L g12606 ( 
.A(n_12073),
.B(n_10970),
.Y(n_12606)
);

AND2x2_ASAP7_75t_L g12607 ( 
.A(n_11438),
.B(n_10858),
.Y(n_12607)
);

AOI22xp33_ASAP7_75t_L g12608 ( 
.A1(n_12012),
.A2(n_9005),
.B1(n_9015),
.B2(n_8322),
.Y(n_12608)
);

AND2x2_ASAP7_75t_L g12609 ( 
.A(n_11678),
.B(n_10858),
.Y(n_12609)
);

AOI22xp33_ASAP7_75t_L g12610 ( 
.A1(n_11244),
.A2(n_8322),
.B1(n_10631),
.B2(n_10110),
.Y(n_12610)
);

OAI221xp5_ASAP7_75t_L g12611 ( 
.A1(n_11539),
.A2(n_10882),
.B1(n_10892),
.B2(n_10846),
.C(n_10843),
.Y(n_12611)
);

HB1xp67_ASAP7_75t_L g12612 ( 
.A(n_11481),
.Y(n_12612)
);

AOI22xp33_ASAP7_75t_L g12613 ( 
.A1(n_11244),
.A2(n_8322),
.B1(n_8733),
.B2(n_8662),
.Y(n_12613)
);

BUFx6f_ASAP7_75t_L g12614 ( 
.A(n_11041),
.Y(n_12614)
);

AOI22xp33_ASAP7_75t_L g12615 ( 
.A1(n_11284),
.A2(n_8733),
.B1(n_8662),
.B2(n_10449),
.Y(n_12615)
);

NOR2xp33_ASAP7_75t_L g12616 ( 
.A(n_11663),
.B(n_10168),
.Y(n_12616)
);

NAND3xp33_ASAP7_75t_L g12617 ( 
.A(n_11339),
.B(n_11377),
.C(n_11366),
.Y(n_12617)
);

OAI22xp5_ASAP7_75t_L g12618 ( 
.A1(n_11679),
.A2(n_8468),
.B1(n_9081),
.B2(n_9037),
.Y(n_12618)
);

BUFx2_ASAP7_75t_L g12619 ( 
.A(n_11990),
.Y(n_12619)
);

OAI221xp5_ASAP7_75t_L g12620 ( 
.A1(n_11561),
.A2(n_10913),
.B1(n_10910),
.B2(n_10385),
.C(n_10386),
.Y(n_12620)
);

OA21x2_ASAP7_75t_L g12621 ( 
.A1(n_11753),
.A2(n_10827),
.B(n_9669),
.Y(n_12621)
);

AOI22xp33_ASAP7_75t_L g12622 ( 
.A1(n_11366),
.A2(n_10449),
.B1(n_10715),
.B2(n_8764),
.Y(n_12622)
);

BUFx3_ASAP7_75t_L g12623 ( 
.A(n_12168),
.Y(n_12623)
);

AOI22xp33_ASAP7_75t_SL g12624 ( 
.A1(n_12175),
.A2(n_8663),
.B1(n_8703),
.B2(n_8659),
.Y(n_12624)
);

AOI22xp33_ASAP7_75t_L g12625 ( 
.A1(n_11377),
.A2(n_8764),
.B1(n_8735),
.B2(n_8295),
.Y(n_12625)
);

AND2x2_ASAP7_75t_L g12626 ( 
.A(n_11678),
.B(n_10858),
.Y(n_12626)
);

AOI22xp33_ASAP7_75t_L g12627 ( 
.A1(n_11561),
.A2(n_8735),
.B1(n_8295),
.B2(n_10751),
.Y(n_12627)
);

AOI22xp33_ASAP7_75t_L g12628 ( 
.A1(n_11562),
.A2(n_8295),
.B1(n_10774),
.B2(n_10757),
.Y(n_12628)
);

CKINVDCx5p33_ASAP7_75t_R g12629 ( 
.A(n_11663),
.Y(n_12629)
);

OAI22xp5_ASAP7_75t_L g12630 ( 
.A1(n_11608),
.A2(n_11023),
.B1(n_10971),
.B2(n_9056),
.Y(n_12630)
);

INVx1_ASAP7_75t_L g12631 ( 
.A(n_11800),
.Y(n_12631)
);

HB1xp67_ASAP7_75t_L g12632 ( 
.A(n_11481),
.Y(n_12632)
);

OAI22xp5_ASAP7_75t_SL g12633 ( 
.A1(n_12238),
.A2(n_9830),
.B1(n_10002),
.B2(n_9910),
.Y(n_12633)
);

HB1xp67_ASAP7_75t_L g12634 ( 
.A(n_11428),
.Y(n_12634)
);

AND2x4_ASAP7_75t_L g12635 ( 
.A(n_11857),
.B(n_10009),
.Y(n_12635)
);

INVx1_ASAP7_75t_L g12636 ( 
.A(n_11802),
.Y(n_12636)
);

AOI22xp5_ASAP7_75t_L g12637 ( 
.A1(n_12200),
.A2(n_10207),
.B1(n_9348),
.B2(n_9354),
.Y(n_12637)
);

AOI221xp5_ASAP7_75t_L g12638 ( 
.A1(n_11562),
.A2(n_10244),
.B1(n_10257),
.B2(n_10240),
.C(n_10237),
.Y(n_12638)
);

OAI22xp5_ASAP7_75t_L g12639 ( 
.A1(n_11608),
.A2(n_11023),
.B1(n_10971),
.B2(n_9056),
.Y(n_12639)
);

INVx1_ASAP7_75t_L g12640 ( 
.A(n_11802),
.Y(n_12640)
);

AND2x2_ASAP7_75t_L g12641 ( 
.A(n_11761),
.B(n_10889),
.Y(n_12641)
);

AND2x4_ASAP7_75t_L g12642 ( 
.A(n_11857),
.B(n_11880),
.Y(n_12642)
);

CKINVDCx5p33_ASAP7_75t_R g12643 ( 
.A(n_11719),
.Y(n_12643)
);

AOI221xp5_ASAP7_75t_L g12644 ( 
.A1(n_11577),
.A2(n_11578),
.B1(n_11063),
.B2(n_11066),
.C(n_11057),
.Y(n_12644)
);

AOI21xp33_ASAP7_75t_L g12645 ( 
.A1(n_11140),
.A2(n_10304),
.B(n_10298),
.Y(n_12645)
);

OAI21xp33_ASAP7_75t_L g12646 ( 
.A1(n_11140),
.A2(n_10194),
.B(n_10185),
.Y(n_12646)
);

INVx1_ASAP7_75t_SL g12647 ( 
.A(n_12181),
.Y(n_12647)
);

AOI22xp33_ASAP7_75t_L g12648 ( 
.A1(n_11577),
.A2(n_8295),
.B1(n_10775),
.B2(n_8841),
.Y(n_12648)
);

AOI22xp33_ASAP7_75t_SL g12649 ( 
.A1(n_12175),
.A2(n_8663),
.B1(n_8703),
.B2(n_8659),
.Y(n_12649)
);

BUFx4f_ASAP7_75t_L g12650 ( 
.A(n_11041),
.Y(n_12650)
);

AOI22xp5_ASAP7_75t_L g12651 ( 
.A1(n_12200),
.A2(n_10207),
.B1(n_9348),
.B2(n_9354),
.Y(n_12651)
);

CKINVDCx5p33_ASAP7_75t_R g12652 ( 
.A(n_11719),
.Y(n_12652)
);

AOI22xp33_ASAP7_75t_L g12653 ( 
.A1(n_11578),
.A2(n_8295),
.B1(n_8841),
.B2(n_8470),
.Y(n_12653)
);

AOI22xp33_ASAP7_75t_L g12654 ( 
.A1(n_11768),
.A2(n_11782),
.B1(n_11804),
.B2(n_11786),
.Y(n_12654)
);

AND2x2_ASAP7_75t_L g12655 ( 
.A(n_11761),
.B(n_10889),
.Y(n_12655)
);

BUFx8_ASAP7_75t_L g12656 ( 
.A(n_11078),
.Y(n_12656)
);

AOI22xp5_ASAP7_75t_L g12657 ( 
.A1(n_11072),
.A2(n_8448),
.B1(n_8750),
.B2(n_8290),
.Y(n_12657)
);

OR2x2_ASAP7_75t_L g12658 ( 
.A(n_12028),
.B(n_10185),
.Y(n_12658)
);

NAND2xp5_ASAP7_75t_L g12659 ( 
.A(n_11508),
.B(n_10194),
.Y(n_12659)
);

AOI22xp33_ASAP7_75t_L g12660 ( 
.A1(n_11768),
.A2(n_11782),
.B1(n_11804),
.B2(n_11786),
.Y(n_12660)
);

BUFx2_ASAP7_75t_L g12661 ( 
.A(n_11380),
.Y(n_12661)
);

NOR2xp33_ASAP7_75t_L g12662 ( 
.A(n_12227),
.B(n_10168),
.Y(n_12662)
);

INVx3_ASAP7_75t_L g12663 ( 
.A(n_11491),
.Y(n_12663)
);

AOI22xp33_ASAP7_75t_L g12664 ( 
.A1(n_11808),
.A2(n_8470),
.B1(n_8167),
.B2(n_10361),
.Y(n_12664)
);

AOI22xp33_ASAP7_75t_L g12665 ( 
.A1(n_11808),
.A2(n_8167),
.B1(n_10375),
.B2(n_9649),
.Y(n_12665)
);

INVx1_ASAP7_75t_L g12666 ( 
.A(n_11806),
.Y(n_12666)
);

AND2x2_ASAP7_75t_L g12667 ( 
.A(n_12095),
.B(n_10889),
.Y(n_12667)
);

AND2x2_ASAP7_75t_L g12668 ( 
.A(n_11652),
.B(n_10889),
.Y(n_12668)
);

HB1xp67_ASAP7_75t_L g12669 ( 
.A(n_11428),
.Y(n_12669)
);

INVx1_ASAP7_75t_L g12670 ( 
.A(n_11806),
.Y(n_12670)
);

AO31x2_ASAP7_75t_L g12671 ( 
.A1(n_11708),
.A2(n_10886),
.A3(n_10763),
.B(n_10555),
.Y(n_12671)
);

OAI221xp5_ASAP7_75t_L g12672 ( 
.A1(n_12207),
.A2(n_9744),
.B1(n_9761),
.B2(n_9691),
.C(n_9613),
.Y(n_12672)
);

OAI221xp5_ASAP7_75t_L g12673 ( 
.A1(n_12207),
.A2(n_9795),
.B1(n_9941),
.B2(n_9863),
.C(n_9847),
.Y(n_12673)
);

AOI22xp5_ASAP7_75t_L g12674 ( 
.A1(n_11113),
.A2(n_8448),
.B1(n_8750),
.B2(n_8290),
.Y(n_12674)
);

INVx1_ASAP7_75t_L g12675 ( 
.A(n_11027),
.Y(n_12675)
);

AOI21xp33_ASAP7_75t_L g12676 ( 
.A1(n_11161),
.A2(n_11243),
.B(n_11652),
.Y(n_12676)
);

NAND2xp5_ASAP7_75t_L g12677 ( 
.A(n_11508),
.B(n_10214),
.Y(n_12677)
);

BUFx3_ASAP7_75t_L g12678 ( 
.A(n_11103),
.Y(n_12678)
);

AOI22xp33_ASAP7_75t_L g12679 ( 
.A1(n_11809),
.A2(n_8167),
.B1(n_9649),
.B2(n_9646),
.Y(n_12679)
);

OAI21xp5_ASAP7_75t_SL g12680 ( 
.A1(n_11200),
.A2(n_10930),
.B(n_10909),
.Y(n_12680)
);

NAND2xp5_ASAP7_75t_L g12681 ( 
.A(n_11525),
.B(n_10214),
.Y(n_12681)
);

AOI22xp33_ASAP7_75t_SL g12682 ( 
.A1(n_11296),
.A2(n_8663),
.B1(n_8703),
.B2(n_8659),
.Y(n_12682)
);

AOI22xp33_ASAP7_75t_L g12683 ( 
.A1(n_11809),
.A2(n_8167),
.B1(n_9649),
.B2(n_9646),
.Y(n_12683)
);

OAI22xp5_ASAP7_75t_L g12684 ( 
.A1(n_11671),
.A2(n_9056),
.B1(n_9954),
.B2(n_9953),
.Y(n_12684)
);

OAI221xp5_ASAP7_75t_L g12685 ( 
.A1(n_11296),
.A2(n_10060),
.B1(n_10133),
.B2(n_10058),
.C(n_10005),
.Y(n_12685)
);

CKINVDCx20_ASAP7_75t_R g12686 ( 
.A(n_11582),
.Y(n_12686)
);

INVx2_ASAP7_75t_L g12687 ( 
.A(n_11050),
.Y(n_12687)
);

AOI21x1_ASAP7_75t_L g12688 ( 
.A1(n_11863),
.A2(n_9956),
.B(n_9916),
.Y(n_12688)
);

NAND2xp5_ASAP7_75t_L g12689 ( 
.A(n_11525),
.B(n_11670),
.Y(n_12689)
);

INVx2_ASAP7_75t_L g12690 ( 
.A(n_11071),
.Y(n_12690)
);

OAI33xp33_ASAP7_75t_L g12691 ( 
.A1(n_11934),
.A2(n_10280),
.A3(n_10783),
.B1(n_10711),
.B2(n_8824),
.B3(n_8582),
.Y(n_12691)
);

INVx1_ASAP7_75t_L g12692 ( 
.A(n_11030),
.Y(n_12692)
);

AOI222xp33_ASAP7_75t_L g12693 ( 
.A1(n_11040),
.A2(n_10240),
.B1(n_10244),
.B2(n_10268),
.C1(n_10257),
.C2(n_10237),
.Y(n_12693)
);

OR2x2_ASAP7_75t_L g12694 ( 
.A(n_12039),
.B(n_10280),
.Y(n_12694)
);

AND2x2_ASAP7_75t_L g12695 ( 
.A(n_11671),
.B(n_10957),
.Y(n_12695)
);

AOI22xp33_ASAP7_75t_SL g12696 ( 
.A1(n_11296),
.A2(n_8663),
.B1(n_8703),
.B2(n_8659),
.Y(n_12696)
);

INVxp33_ASAP7_75t_L g12697 ( 
.A(n_11777),
.Y(n_12697)
);

OAI22xp5_ASAP7_75t_L g12698 ( 
.A1(n_11723),
.A2(n_9056),
.B1(n_9954),
.B2(n_9953),
.Y(n_12698)
);

HB1xp67_ASAP7_75t_L g12699 ( 
.A(n_11670),
.Y(n_12699)
);

INVx4_ASAP7_75t_L g12700 ( 
.A(n_11078),
.Y(n_12700)
);

AND2x2_ASAP7_75t_L g12701 ( 
.A(n_11723),
.B(n_10957),
.Y(n_12701)
);

INVx1_ASAP7_75t_L g12702 ( 
.A(n_11037),
.Y(n_12702)
);

INVx2_ASAP7_75t_L g12703 ( 
.A(n_11071),
.Y(n_12703)
);

OR2x2_ASAP7_75t_L g12704 ( 
.A(n_11754),
.B(n_10711),
.Y(n_12704)
);

OAI221xp5_ASAP7_75t_L g12705 ( 
.A1(n_11040),
.A2(n_10162),
.B1(n_10179),
.B2(n_10149),
.C(n_10145),
.Y(n_12705)
);

NAND4xp25_ASAP7_75t_L g12706 ( 
.A(n_12047),
.B(n_10081),
.C(n_10086),
.D(n_10009),
.Y(n_12706)
);

AOI221xp5_ASAP7_75t_L g12707 ( 
.A1(n_11057),
.A2(n_10257),
.B1(n_10268),
.B2(n_10244),
.C(n_10240),
.Y(n_12707)
);

AND2x2_ASAP7_75t_L g12708 ( 
.A(n_12256),
.B(n_10957),
.Y(n_12708)
);

AOI222xp33_ASAP7_75t_L g12709 ( 
.A1(n_11063),
.A2(n_10287),
.B1(n_10297),
.B2(n_10308),
.C1(n_10305),
.C2(n_10268),
.Y(n_12709)
);

AND2x2_ASAP7_75t_L g12710 ( 
.A(n_12211),
.B(n_10957),
.Y(n_12710)
);

INVx1_ASAP7_75t_L g12711 ( 
.A(n_11049),
.Y(n_12711)
);

A2O1A1Ixp33_ASAP7_75t_L g12712 ( 
.A1(n_11334),
.A2(n_10297),
.B(n_10305),
.C(n_10287),
.Y(n_12712)
);

INVx2_ASAP7_75t_L g12713 ( 
.A(n_11085),
.Y(n_12713)
);

AOI22xp33_ASAP7_75t_L g12714 ( 
.A1(n_12259),
.A2(n_8167),
.B1(n_9649),
.B2(n_9646),
.Y(n_12714)
);

INVx2_ASAP7_75t_L g12715 ( 
.A(n_11085),
.Y(n_12715)
);

INVx1_ASAP7_75t_L g12716 ( 
.A(n_11053),
.Y(n_12716)
);

AOI22xp33_ASAP7_75t_L g12717 ( 
.A1(n_12090),
.A2(n_8167),
.B1(n_9646),
.B2(n_9048),
.Y(n_12717)
);

AOI211xp5_ASAP7_75t_L g12718 ( 
.A1(n_11139),
.A2(n_12197),
.B(n_11756),
.C(n_11334),
.Y(n_12718)
);

INVx2_ASAP7_75t_L g12719 ( 
.A(n_11196),
.Y(n_12719)
);

CKINVDCx5p33_ASAP7_75t_R g12720 ( 
.A(n_11132),
.Y(n_12720)
);

NOR2xp33_ASAP7_75t_L g12721 ( 
.A(n_12227),
.B(n_9811),
.Y(n_12721)
);

OAI21xp5_ASAP7_75t_L g12722 ( 
.A1(n_11139),
.A2(n_8528),
.B(n_8534),
.Y(n_12722)
);

OAI221xp5_ASAP7_75t_L g12723 ( 
.A1(n_11066),
.A2(n_10227),
.B1(n_10184),
.B2(n_10297),
.C(n_10287),
.Y(n_12723)
);

OR2x6_ASAP7_75t_L g12724 ( 
.A(n_11078),
.B(n_9894),
.Y(n_12724)
);

OAI22xp5_ASAP7_75t_L g12725 ( 
.A1(n_11879),
.A2(n_9954),
.B1(n_9970),
.B2(n_9953),
.Y(n_12725)
);

AOI22xp33_ASAP7_75t_L g12726 ( 
.A1(n_12255),
.A2(n_9048),
.B1(n_8663),
.B2(n_8703),
.Y(n_12726)
);

AOI22xp33_ASAP7_75t_L g12727 ( 
.A1(n_12255),
.A2(n_12098),
.B1(n_12099),
.B2(n_12090),
.Y(n_12727)
);

BUFx4f_ASAP7_75t_SL g12728 ( 
.A(n_12236),
.Y(n_12728)
);

AND2x2_ASAP7_75t_L g12729 ( 
.A(n_12249),
.B(n_12252),
.Y(n_12729)
);

AOI22xp33_ASAP7_75t_L g12730 ( 
.A1(n_12259),
.A2(n_9048),
.B1(n_8663),
.B2(n_8703),
.Y(n_12730)
);

A2O1A1Ixp33_ASAP7_75t_L g12731 ( 
.A1(n_11151),
.A2(n_10308),
.B(n_10311),
.C(n_10305),
.Y(n_12731)
);

AOI22xp33_ASAP7_75t_L g12732 ( 
.A1(n_12098),
.A2(n_9048),
.B1(n_8741),
.B2(n_8797),
.Y(n_12732)
);

AND2x4_ASAP7_75t_L g12733 ( 
.A(n_11880),
.B(n_10081),
.Y(n_12733)
);

AOI22xp5_ASAP7_75t_L g12734 ( 
.A1(n_11236),
.A2(n_8348),
.B1(n_10129),
.B2(n_10034),
.Y(n_12734)
);

AOI22x1_ASAP7_75t_L g12735 ( 
.A1(n_11877),
.A2(n_9845),
.B1(n_9934),
.B2(n_9774),
.Y(n_12735)
);

AND2x4_ASAP7_75t_L g12736 ( 
.A(n_11902),
.B(n_10081),
.Y(n_12736)
);

AOI22xp5_ASAP7_75t_L g12737 ( 
.A1(n_11255),
.A2(n_8348),
.B1(n_10129),
.B2(n_10034),
.Y(n_12737)
);

AOI221xp5_ASAP7_75t_L g12738 ( 
.A1(n_11073),
.A2(n_10316),
.B1(n_10335),
.B2(n_10311),
.C(n_10308),
.Y(n_12738)
);

INVxp33_ASAP7_75t_L g12739 ( 
.A(n_11777),
.Y(n_12739)
);

INVx1_ASAP7_75t_L g12740 ( 
.A(n_11058),
.Y(n_12740)
);

OAI211xp5_ASAP7_75t_L g12741 ( 
.A1(n_11042),
.A2(n_10298),
.B(n_10304),
.C(n_10755),
.Y(n_12741)
);

INVx2_ASAP7_75t_L g12742 ( 
.A(n_11196),
.Y(n_12742)
);

AOI22xp5_ASAP7_75t_L g12743 ( 
.A1(n_11288),
.A2(n_9800),
.B1(n_8374),
.B2(n_8493),
.Y(n_12743)
);

CKINVDCx20_ASAP7_75t_R g12744 ( 
.A(n_11817),
.Y(n_12744)
);

INVx2_ASAP7_75t_L g12745 ( 
.A(n_11237),
.Y(n_12745)
);

AND2x6_ASAP7_75t_L g12746 ( 
.A(n_11580),
.B(n_10086),
.Y(n_12746)
);

OAI332xp33_ASAP7_75t_L g12747 ( 
.A1(n_11314),
.A2(n_10316),
.A3(n_10335),
.B1(n_10311),
.B2(n_10939),
.B3(n_10946),
.C1(n_10942),
.C2(n_10935),
.Y(n_12747)
);

INVx2_ASAP7_75t_L g12748 ( 
.A(n_11237),
.Y(n_12748)
);

OAI221xp5_ASAP7_75t_L g12749 ( 
.A1(n_11073),
.A2(n_10335),
.B1(n_10316),
.B2(n_10927),
.C(n_10925),
.Y(n_12749)
);

INVx1_ASAP7_75t_L g12750 ( 
.A(n_11060),
.Y(n_12750)
);

INVxp67_ASAP7_75t_SL g12751 ( 
.A(n_11830),
.Y(n_12751)
);

HB1xp67_ASAP7_75t_L g12752 ( 
.A(n_11682),
.Y(n_12752)
);

BUFx12f_ASAP7_75t_L g12753 ( 
.A(n_11078),
.Y(n_12753)
);

INVx6_ASAP7_75t_SL g12754 ( 
.A(n_11249),
.Y(n_12754)
);

AOI22xp33_ASAP7_75t_L g12755 ( 
.A1(n_12245),
.A2(n_9048),
.B1(n_8741),
.B2(n_8797),
.Y(n_12755)
);

OAI22xp5_ASAP7_75t_L g12756 ( 
.A1(n_11879),
.A2(n_9954),
.B1(n_9970),
.B2(n_9953),
.Y(n_12756)
);

OAI221xp5_ASAP7_75t_L g12757 ( 
.A1(n_11075),
.A2(n_10445),
.B1(n_10791),
.B2(n_9908),
.C(n_9919),
.Y(n_12757)
);

INVx1_ASAP7_75t_L g12758 ( 
.A(n_11064),
.Y(n_12758)
);

NAND2xp5_ASAP7_75t_L g12759 ( 
.A(n_11682),
.B(n_9136),
.Y(n_12759)
);

O2A1O1Ixp33_ASAP7_75t_L g12760 ( 
.A1(n_11075),
.A2(n_10939),
.B(n_10942),
.C(n_10935),
.Y(n_12760)
);

AO21x2_ASAP7_75t_L g12761 ( 
.A1(n_11708),
.A2(n_10808),
.B(n_10159),
.Y(n_12761)
);

OAI22xp5_ASAP7_75t_L g12762 ( 
.A1(n_11439),
.A2(n_9954),
.B1(n_9970),
.B2(n_9953),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_11159),
.B(n_10086),
.Y(n_12763)
);

OAI221xp5_ASAP7_75t_SL g12764 ( 
.A1(n_11076),
.A2(n_10935),
.B1(n_10946),
.B2(n_10942),
.C(n_10939),
.Y(n_12764)
);

NAND3xp33_ASAP7_75t_L g12765 ( 
.A(n_11707),
.B(n_11749),
.C(n_11730),
.Y(n_12765)
);

AOI22xp33_ASAP7_75t_L g12766 ( 
.A1(n_12099),
.A2(n_9048),
.B1(n_8741),
.B2(n_8797),
.Y(n_12766)
);

BUFx3_ASAP7_75t_L g12767 ( 
.A(n_11103),
.Y(n_12767)
);

INVx1_ASAP7_75t_L g12768 ( 
.A(n_11065),
.Y(n_12768)
);

AOI22xp5_ASAP7_75t_L g12769 ( 
.A1(n_11706),
.A2(n_8374),
.B1(n_8493),
.B2(n_8331),
.Y(n_12769)
);

AOI22xp33_ASAP7_75t_L g12770 ( 
.A1(n_12240),
.A2(n_8741),
.B1(n_8797),
.B2(n_8659),
.Y(n_12770)
);

CKINVDCx11_ASAP7_75t_R g12771 ( 
.A(n_12186),
.Y(n_12771)
);

INVx1_ASAP7_75t_L g12772 ( 
.A(n_11067),
.Y(n_12772)
);

AOI22xp33_ASAP7_75t_L g12773 ( 
.A1(n_12245),
.A2(n_8741),
.B1(n_8797),
.B2(n_8659),
.Y(n_12773)
);

OAI22xp5_ASAP7_75t_L g12774 ( 
.A1(n_12242),
.A2(n_9999),
.B1(n_10012),
.B2(n_9970),
.Y(n_12774)
);

OAI22xp33_ASAP7_75t_L g12775 ( 
.A1(n_11076),
.A2(n_9290),
.B1(n_8134),
.B2(n_9125),
.Y(n_12775)
);

OAI22xp5_ASAP7_75t_L g12776 ( 
.A1(n_11838),
.A2(n_9999),
.B1(n_10012),
.B2(n_9970),
.Y(n_12776)
);

OR2x6_ASAP7_75t_L g12777 ( 
.A(n_11152),
.B(n_7326),
.Y(n_12777)
);

AND2x2_ASAP7_75t_L g12778 ( 
.A(n_12248),
.B(n_10395),
.Y(n_12778)
);

CKINVDCx20_ASAP7_75t_R g12779 ( 
.A(n_11817),
.Y(n_12779)
);

AOI22xp33_ASAP7_75t_L g12780 ( 
.A1(n_12104),
.A2(n_8797),
.B1(n_8823),
.B2(n_8741),
.Y(n_12780)
);

NAND2x1_ASAP7_75t_L g12781 ( 
.A(n_12170),
.B(n_9896),
.Y(n_12781)
);

AND2x2_ASAP7_75t_L g12782 ( 
.A(n_12131),
.B(n_10395),
.Y(n_12782)
);

AND2x2_ASAP7_75t_L g12783 ( 
.A(n_12147),
.B(n_10395),
.Y(n_12783)
);

NAND2xp5_ASAP7_75t_L g12784 ( 
.A(n_11707),
.B(n_9136),
.Y(n_12784)
);

INVx8_ASAP7_75t_L g12785 ( 
.A(n_11152),
.Y(n_12785)
);

BUFx12f_ASAP7_75t_L g12786 ( 
.A(n_11152),
.Y(n_12786)
);

AND2x2_ASAP7_75t_L g12787 ( 
.A(n_11815),
.B(n_10395),
.Y(n_12787)
);

AOI22xp33_ASAP7_75t_L g12788 ( 
.A1(n_12104),
.A2(n_8856),
.B1(n_8929),
.B2(n_8823),
.Y(n_12788)
);

AOI22xp33_ASAP7_75t_L g12789 ( 
.A1(n_12231),
.A2(n_8856),
.B1(n_8929),
.B2(n_8823),
.Y(n_12789)
);

NAND3xp33_ASAP7_75t_L g12790 ( 
.A(n_11730),
.B(n_10304),
.C(n_10847),
.Y(n_12790)
);

AND2x2_ASAP7_75t_L g12791 ( 
.A(n_11845),
.B(n_10395),
.Y(n_12791)
);

BUFx12f_ASAP7_75t_L g12792 ( 
.A(n_11152),
.Y(n_12792)
);

OR2x2_ASAP7_75t_L g12793 ( 
.A(n_12124),
.B(n_10783),
.Y(n_12793)
);

OR2x2_ASAP7_75t_L g12794 ( 
.A(n_12137),
.B(n_9079),
.Y(n_12794)
);

INVx2_ASAP7_75t_L g12795 ( 
.A(n_11960),
.Y(n_12795)
);

OAI22xp5_ASAP7_75t_L g12796 ( 
.A1(n_12122),
.A2(n_10012),
.B1(n_10350),
.B2(n_9999),
.Y(n_12796)
);

NAND3xp33_ASAP7_75t_L g12797 ( 
.A(n_11749),
.B(n_10847),
.C(n_9918),
.Y(n_12797)
);

AND2x2_ASAP7_75t_L g12798 ( 
.A(n_11865),
.B(n_10395),
.Y(n_12798)
);

INVx1_ASAP7_75t_L g12799 ( 
.A(n_11080),
.Y(n_12799)
);

AOI22xp33_ASAP7_75t_L g12800 ( 
.A1(n_12106),
.A2(n_8856),
.B1(n_8929),
.B2(n_8823),
.Y(n_12800)
);

AND2x2_ASAP7_75t_L g12801 ( 
.A(n_11883),
.B(n_10457),
.Y(n_12801)
);

AOI22xp33_ASAP7_75t_L g12802 ( 
.A1(n_12106),
.A2(n_12107),
.B1(n_12121),
.B2(n_12110),
.Y(n_12802)
);

OR2x2_ASAP7_75t_L g12803 ( 
.A(n_12144),
.B(n_9079),
.Y(n_12803)
);

NAND2xp5_ASAP7_75t_L g12804 ( 
.A(n_11764),
.B(n_9136),
.Y(n_12804)
);

OAI22xp33_ASAP7_75t_L g12805 ( 
.A1(n_11079),
.A2(n_9290),
.B1(n_9125),
.B2(n_8331),
.Y(n_12805)
);

NOR3xp33_ASAP7_75t_L g12806 ( 
.A(n_11902),
.B(n_10095),
.C(n_10755),
.Y(n_12806)
);

INVx1_ASAP7_75t_L g12807 ( 
.A(n_11091),
.Y(n_12807)
);

INVx3_ASAP7_75t_L g12808 ( 
.A(n_11491),
.Y(n_12808)
);

AOI21xp33_ASAP7_75t_L g12809 ( 
.A1(n_11161),
.A2(n_10918),
.B(n_10877),
.Y(n_12809)
);

AOI22xp5_ASAP7_75t_L g12810 ( 
.A1(n_11830),
.A2(n_8900),
.B1(n_8607),
.B2(n_9134),
.Y(n_12810)
);

AND2x2_ASAP7_75t_L g12811 ( 
.A(n_11885),
.B(n_10457),
.Y(n_12811)
);

OAI22xp33_ASAP7_75t_L g12812 ( 
.A1(n_11079),
.A2(n_9125),
.B1(n_8900),
.B2(n_8607),
.Y(n_12812)
);

OAI221xp5_ASAP7_75t_L g12813 ( 
.A1(n_11712),
.A2(n_9908),
.B1(n_9919),
.B2(n_9906),
.C(n_9901),
.Y(n_12813)
);

AND2x4_ASAP7_75t_L g12814 ( 
.A(n_11995),
.B(n_9833),
.Y(n_12814)
);

AOI22xp33_ASAP7_75t_L g12815 ( 
.A1(n_12240),
.A2(n_8856),
.B1(n_8929),
.B2(n_8823),
.Y(n_12815)
);

OAI211xp5_ASAP7_75t_SL g12816 ( 
.A1(n_11995),
.A2(n_10962),
.B(n_10788),
.C(n_9866),
.Y(n_12816)
);

AOI221xp5_ASAP7_75t_L g12817 ( 
.A1(n_11712),
.A2(n_11734),
.B1(n_11736),
.B2(n_11726),
.C(n_11725),
.Y(n_12817)
);

AND2x2_ASAP7_75t_L g12818 ( 
.A(n_11887),
.B(n_10457),
.Y(n_12818)
);

BUFx8_ASAP7_75t_L g12819 ( 
.A(n_11166),
.Y(n_12819)
);

AOI22xp33_ASAP7_75t_L g12820 ( 
.A1(n_12107),
.A2(n_8856),
.B1(n_8929),
.B2(n_8823),
.Y(n_12820)
);

AOI22xp33_ASAP7_75t_SL g12821 ( 
.A1(n_11151),
.A2(n_8856),
.B1(n_8984),
.B2(n_8929),
.Y(n_12821)
);

AOI22xp33_ASAP7_75t_L g12822 ( 
.A1(n_12110),
.A2(n_8984),
.B1(n_8988),
.B2(n_9183),
.Y(n_12822)
);

OAI221xp5_ASAP7_75t_L g12823 ( 
.A1(n_11725),
.A2(n_9908),
.B1(n_9919),
.B2(n_9906),
.C(n_9901),
.Y(n_12823)
);

AOI221xp5_ASAP7_75t_L g12824 ( 
.A1(n_11726),
.A2(n_9920),
.B1(n_9924),
.B2(n_9906),
.C(n_9901),
.Y(n_12824)
);

AOI22xp33_ASAP7_75t_L g12825 ( 
.A1(n_12121),
.A2(n_8984),
.B1(n_8988),
.B2(n_9183),
.Y(n_12825)
);

INVx1_ASAP7_75t_L g12826 ( 
.A(n_11092),
.Y(n_12826)
);

A2O1A1Ixp33_ASAP7_75t_L g12827 ( 
.A1(n_11391),
.A2(n_9108),
.B(n_9113),
.C(n_9105),
.Y(n_12827)
);

BUFx5_ASAP7_75t_L g12828 ( 
.A(n_11216),
.Y(n_12828)
);

AOI222xp33_ASAP7_75t_L g12829 ( 
.A1(n_11734),
.A2(n_9425),
.B1(n_9416),
.B2(n_9465),
.C1(n_9461),
.C2(n_8942),
.Y(n_12829)
);

OAI211xp5_ASAP7_75t_L g12830 ( 
.A1(n_11764),
.A2(n_10788),
.B(n_10962),
.C(n_8831),
.Y(n_12830)
);

OAI22xp5_ASAP7_75t_L g12831 ( 
.A1(n_11032),
.A2(n_10012),
.B1(n_10350),
.B2(n_9999),
.Y(n_12831)
);

OAI22xp5_ASAP7_75t_L g12832 ( 
.A1(n_11032),
.A2(n_10012),
.B1(n_10350),
.B2(n_9999),
.Y(n_12832)
);

O2A1O1Ixp33_ASAP7_75t_L g12833 ( 
.A1(n_11788),
.A2(n_10947),
.B(n_10963),
.C(n_10946),
.Y(n_12833)
);

INVx2_ASAP7_75t_L g12834 ( 
.A(n_11960),
.Y(n_12834)
);

BUFx3_ASAP7_75t_L g12835 ( 
.A(n_11150),
.Y(n_12835)
);

INVx2_ASAP7_75t_L g12836 ( 
.A(n_11960),
.Y(n_12836)
);

AOI221xp5_ASAP7_75t_L g12837 ( 
.A1(n_11736),
.A2(n_9927),
.B1(n_9933),
.B2(n_9924),
.C(n_9920),
.Y(n_12837)
);

AOI22xp33_ASAP7_75t_L g12838 ( 
.A1(n_12233),
.A2(n_8984),
.B1(n_8988),
.B2(n_9185),
.Y(n_12838)
);

AOI22xp33_ASAP7_75t_L g12839 ( 
.A1(n_12233),
.A2(n_8984),
.B1(n_8988),
.B2(n_9185),
.Y(n_12839)
);

AND2x4_ASAP7_75t_L g12840 ( 
.A(n_12002),
.B(n_9833),
.Y(n_12840)
);

NOR2xp33_ASAP7_75t_L g12841 ( 
.A(n_11150),
.B(n_9811),
.Y(n_12841)
);

OAI22xp5_ASAP7_75t_L g12842 ( 
.A1(n_11032),
.A2(n_10379),
.B1(n_10416),
.B2(n_10350),
.Y(n_12842)
);

AOI221xp5_ASAP7_75t_L g12843 ( 
.A1(n_11738),
.A2(n_9927),
.B1(n_9933),
.B2(n_9924),
.C(n_9920),
.Y(n_12843)
);

OR2x2_ASAP7_75t_L g12844 ( 
.A(n_12160),
.B(n_9079),
.Y(n_12844)
);

OAI22xp5_ASAP7_75t_L g12845 ( 
.A1(n_11201),
.A2(n_10379),
.B1(n_10416),
.B2(n_10350),
.Y(n_12845)
);

AND2x2_ASAP7_75t_L g12846 ( 
.A(n_11891),
.B(n_10457),
.Y(n_12846)
);

AOI22xp5_ASAP7_75t_L g12847 ( 
.A1(n_11219),
.A2(n_9134),
.B1(n_9179),
.B2(n_10847),
.Y(n_12847)
);

OAI22xp5_ASAP7_75t_L g12848 ( 
.A1(n_11201),
.A2(n_10416),
.B1(n_10379),
.B2(n_9184),
.Y(n_12848)
);

INVx2_ASAP7_75t_L g12849 ( 
.A(n_12084),
.Y(n_12849)
);

AO31x2_ASAP7_75t_L g12850 ( 
.A1(n_11738),
.A2(n_10947),
.A3(n_10963),
.B(n_10095),
.Y(n_12850)
);

AOI22xp5_ASAP7_75t_L g12851 ( 
.A1(n_11357),
.A2(n_9179),
.B1(n_9216),
.B2(n_9057),
.Y(n_12851)
);

BUFx10_ASAP7_75t_L g12852 ( 
.A(n_11166),
.Y(n_12852)
);

AOI22xp33_ASAP7_75t_L g12853 ( 
.A1(n_12126),
.A2(n_8984),
.B1(n_8988),
.B2(n_8847),
.Y(n_12853)
);

OAI221xp5_ASAP7_75t_L g12854 ( 
.A1(n_11742),
.A2(n_9940),
.B1(n_9946),
.B2(n_9933),
.C(n_9927),
.Y(n_12854)
);

AOI221xp5_ASAP7_75t_L g12855 ( 
.A1(n_11742),
.A2(n_9948),
.B1(n_9951),
.B2(n_9946),
.C(n_9940),
.Y(n_12855)
);

OAI211xp5_ASAP7_75t_SL g12856 ( 
.A1(n_12002),
.A2(n_9872),
.B(n_9881),
.C(n_9866),
.Y(n_12856)
);

OAI221xp5_ASAP7_75t_L g12857 ( 
.A1(n_11762),
.A2(n_9948),
.B1(n_9951),
.B2(n_9946),
.C(n_9940),
.Y(n_12857)
);

OAI21x1_ASAP7_75t_L g12858 ( 
.A1(n_12157),
.A2(n_10159),
.B(n_10317),
.Y(n_12858)
);

AOI22xp33_ASAP7_75t_L g12859 ( 
.A1(n_12126),
.A2(n_8988),
.B1(n_8847),
.B2(n_10006),
.Y(n_12859)
);

INVx4_ASAP7_75t_L g12860 ( 
.A(n_11166),
.Y(n_12860)
);

AND2x2_ASAP7_75t_L g12861 ( 
.A(n_11905),
.B(n_10457),
.Y(n_12861)
);

OAI22xp33_ASAP7_75t_L g12862 ( 
.A1(n_11837),
.A2(n_9125),
.B1(n_10918),
.B2(n_10877),
.Y(n_12862)
);

AOI22xp33_ASAP7_75t_L g12863 ( 
.A1(n_12231),
.A2(n_10016),
.B1(n_10019),
.B2(n_10006),
.Y(n_12863)
);

AOI22xp33_ASAP7_75t_L g12864 ( 
.A1(n_12127),
.A2(n_10016),
.B1(n_10019),
.B2(n_10006),
.Y(n_12864)
);

NAND2xp5_ASAP7_75t_L g12865 ( 
.A(n_11788),
.B(n_9136),
.Y(n_12865)
);

BUFx3_ASAP7_75t_L g12866 ( 
.A(n_12236),
.Y(n_12866)
);

OAI22xp5_ASAP7_75t_L g12867 ( 
.A1(n_11201),
.A2(n_10416),
.B1(n_10379),
.B2(n_9184),
.Y(n_12867)
);

AOI22xp33_ASAP7_75t_L g12868 ( 
.A1(n_12127),
.A2(n_10019),
.B1(n_10021),
.B2(n_10016),
.Y(n_12868)
);

OAI22xp5_ASAP7_75t_L g12869 ( 
.A1(n_11253),
.A2(n_10416),
.B1(n_10379),
.B2(n_9184),
.Y(n_12869)
);

NAND3xp33_ASAP7_75t_L g12870 ( 
.A(n_11977),
.B(n_12007),
.C(n_11987),
.Y(n_12870)
);

OAI21x1_ASAP7_75t_L g12871 ( 
.A1(n_12170),
.A2(n_10325),
.B(n_10317),
.Y(n_12871)
);

AOI22xp33_ASAP7_75t_L g12872 ( 
.A1(n_12136),
.A2(n_10025),
.B1(n_10035),
.B2(n_10021),
.Y(n_12872)
);

AOI22xp5_ASAP7_75t_L g12873 ( 
.A1(n_11368),
.A2(n_9216),
.B1(n_9057),
.B2(n_9267),
.Y(n_12873)
);

INVx2_ASAP7_75t_L g12874 ( 
.A(n_12084),
.Y(n_12874)
);

AOI21xp33_ASAP7_75t_L g12875 ( 
.A1(n_11243),
.A2(n_10989),
.B(n_9918),
.Y(n_12875)
);

OAI211xp5_ASAP7_75t_L g12876 ( 
.A1(n_11710),
.A2(n_8831),
.B(n_10095),
.C(n_10029),
.Y(n_12876)
);

AOI22xp33_ASAP7_75t_L g12877 ( 
.A1(n_12136),
.A2(n_10025),
.B1(n_10035),
.B2(n_10021),
.Y(n_12877)
);

NAND2x1_ASAP7_75t_L g12878 ( 
.A(n_12191),
.B(n_10325),
.Y(n_12878)
);

INVx1_ASAP7_75t_L g12879 ( 
.A(n_11096),
.Y(n_12879)
);

AND2x4_ASAP7_75t_L g12880 ( 
.A(n_12030),
.B(n_9833),
.Y(n_12880)
);

AOI22xp33_ASAP7_75t_L g12881 ( 
.A1(n_12140),
.A2(n_10035),
.B1(n_10036),
.B2(n_10025),
.Y(n_12881)
);

NAND2xp5_ASAP7_75t_L g12882 ( 
.A(n_12051),
.B(n_9136),
.Y(n_12882)
);

OAI22xp5_ASAP7_75t_L g12883 ( 
.A1(n_11253),
.A2(n_8956),
.B1(n_8817),
.B2(n_8746),
.Y(n_12883)
);

AOI22xp33_ASAP7_75t_SL g12884 ( 
.A1(n_11391),
.A2(n_9125),
.B1(n_8613),
.B2(n_10036),
.Y(n_12884)
);

INVx1_ASAP7_75t_L g12885 ( 
.A(n_11102),
.Y(n_12885)
);

INVx2_ASAP7_75t_L g12886 ( 
.A(n_12084),
.Y(n_12886)
);

AND2x2_ASAP7_75t_L g12887 ( 
.A(n_11906),
.B(n_10457),
.Y(n_12887)
);

AO221x1_ASAP7_75t_L g12888 ( 
.A1(n_11940),
.A2(n_10327),
.B1(n_10808),
.B2(n_11317),
.C(n_11298),
.Y(n_12888)
);

OR2x6_ASAP7_75t_L g12889 ( 
.A(n_11166),
.B(n_11194),
.Y(n_12889)
);

AOI222xp33_ASAP7_75t_L g12890 ( 
.A1(n_11762),
.A2(n_9425),
.B1(n_9416),
.B2(n_9465),
.C1(n_9461),
.C2(n_8942),
.Y(n_12890)
);

OAI211xp5_ASAP7_75t_SL g12891 ( 
.A1(n_12030),
.A2(n_9872),
.B(n_9881),
.C(n_9866),
.Y(n_12891)
);

AND2x2_ASAP7_75t_L g12892 ( 
.A(n_11917),
.B(n_9774),
.Y(n_12892)
);

OAI22xp33_ASAP7_75t_L g12893 ( 
.A1(n_11591),
.A2(n_10989),
.B1(n_9267),
.B2(n_8829),
.Y(n_12893)
);

INVx2_ASAP7_75t_L g12894 ( 
.A(n_11977),
.Y(n_12894)
);

NAND3xp33_ASAP7_75t_L g12895 ( 
.A(n_11977),
.B(n_9918),
.C(n_9911),
.Y(n_12895)
);

INVx1_ASAP7_75t_L g12896 ( 
.A(n_11104),
.Y(n_12896)
);

AOI22xp33_ASAP7_75t_L g12897 ( 
.A1(n_12140),
.A2(n_10045),
.B1(n_10062),
.B2(n_10036),
.Y(n_12897)
);

AOI22xp33_ASAP7_75t_SL g12898 ( 
.A1(n_11482),
.A2(n_8613),
.B1(n_10062),
.B2(n_10045),
.Y(n_12898)
);

AOI211xp5_ASAP7_75t_L g12899 ( 
.A1(n_11056),
.A2(n_10947),
.B(n_10963),
.C(n_8715),
.Y(n_12899)
);

OAI22xp33_ASAP7_75t_L g12900 ( 
.A1(n_11641),
.A2(n_8642),
.B1(n_9453),
.B2(n_8613),
.Y(n_12900)
);

OAI22xp5_ASAP7_75t_L g12901 ( 
.A1(n_11253),
.A2(n_8956),
.B1(n_8817),
.B2(n_8746),
.Y(n_12901)
);

AOI22xp33_ASAP7_75t_L g12902 ( 
.A1(n_12141),
.A2(n_10062),
.B1(n_10064),
.B2(n_10045),
.Y(n_12902)
);

INVx2_ASAP7_75t_L g12903 ( 
.A(n_11977),
.Y(n_12903)
);

A2O1A1Ixp33_ASAP7_75t_L g12904 ( 
.A1(n_11482),
.A2(n_9108),
.B(n_9113),
.C(n_9105),
.Y(n_12904)
);

AOI22xp33_ASAP7_75t_SL g12905 ( 
.A1(n_11417),
.A2(n_8613),
.B1(n_10067),
.B2(n_10064),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_11105),
.Y(n_12906)
);

AOI22xp33_ASAP7_75t_SL g12907 ( 
.A1(n_11417),
.A2(n_8613),
.B1(n_10067),
.B2(n_10064),
.Y(n_12907)
);

BUFx3_ASAP7_75t_L g12908 ( 
.A(n_11710),
.Y(n_12908)
);

INVx2_ASAP7_75t_L g12909 ( 
.A(n_11987),
.Y(n_12909)
);

AOI22xp33_ASAP7_75t_L g12910 ( 
.A1(n_12141),
.A2(n_10073),
.B1(n_10074),
.B2(n_10067),
.Y(n_12910)
);

AOI21xp33_ASAP7_75t_SL g12911 ( 
.A1(n_11654),
.A2(n_8831),
.B(n_8302),
.Y(n_12911)
);

AND2x2_ASAP7_75t_L g12912 ( 
.A(n_11961),
.B(n_9845),
.Y(n_12912)
);

A2O1A1Ixp33_ASAP7_75t_L g12913 ( 
.A1(n_11214),
.A2(n_9108),
.B(n_9113),
.C(n_9105),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_11106),
.Y(n_12914)
);

AOI21xp5_ASAP7_75t_L g12915 ( 
.A1(n_11921),
.A2(n_10611),
.B(n_10504),
.Y(n_12915)
);

OAI22xp33_ASAP7_75t_L g12916 ( 
.A1(n_11155),
.A2(n_8642),
.B1(n_9453),
.B2(n_8613),
.Y(n_12916)
);

AOI22xp33_ASAP7_75t_L g12917 ( 
.A1(n_12150),
.A2(n_10074),
.B1(n_10077),
.B2(n_10073),
.Y(n_12917)
);

INVx2_ASAP7_75t_L g12918 ( 
.A(n_11987),
.Y(n_12918)
);

INVx2_ASAP7_75t_L g12919 ( 
.A(n_11987),
.Y(n_12919)
);

OAI211xp5_ASAP7_75t_L g12920 ( 
.A1(n_11056),
.A2(n_10039),
.B(n_10072),
.C(n_9889),
.Y(n_12920)
);

AND2x4_ASAP7_75t_L g12921 ( 
.A(n_12065),
.B(n_9841),
.Y(n_12921)
);

INVx3_ASAP7_75t_L g12922 ( 
.A(n_11515),
.Y(n_12922)
);

OAI211xp5_ASAP7_75t_L g12923 ( 
.A1(n_11097),
.A2(n_10142),
.B(n_8746),
.C(n_9872),
.Y(n_12923)
);

OAI22xp33_ASAP7_75t_L g12924 ( 
.A1(n_11155),
.A2(n_10731),
.B1(n_10916),
.B2(n_9022),
.Y(n_12924)
);

AOI22xp33_ASAP7_75t_L g12925 ( 
.A1(n_12150),
.A2(n_10074),
.B1(n_10077),
.B2(n_10073),
.Y(n_12925)
);

AOI22xp33_ASAP7_75t_L g12926 ( 
.A1(n_12151),
.A2(n_10079),
.B1(n_10096),
.B2(n_10077),
.Y(n_12926)
);

OR2x6_ASAP7_75t_L g12927 ( 
.A(n_11194),
.B(n_7382),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_11107),
.Y(n_12928)
);

AOI22xp33_ASAP7_75t_L g12929 ( 
.A1(n_12151),
.A2(n_10096),
.B1(n_10099),
.B2(n_10079),
.Y(n_12929)
);

AND2x2_ASAP7_75t_L g12930 ( 
.A(n_12065),
.B(n_9934),
.Y(n_12930)
);

AOI22xp33_ASAP7_75t_L g12931 ( 
.A1(n_12156),
.A2(n_10096),
.B1(n_10099),
.B2(n_10079),
.Y(n_12931)
);

AOI222xp33_ASAP7_75t_L g12932 ( 
.A1(n_11763),
.A2(n_10122),
.B1(n_10111),
.B2(n_10124),
.C1(n_10118),
.C2(n_10099),
.Y(n_12932)
);

AOI221xp5_ASAP7_75t_L g12933 ( 
.A1(n_11763),
.A2(n_9957),
.B1(n_9961),
.B2(n_9951),
.C(n_9948),
.Y(n_12933)
);

INVx2_ASAP7_75t_L g12934 ( 
.A(n_12007),
.Y(n_12934)
);

AND2x2_ASAP7_75t_L g12935 ( 
.A(n_12094),
.B(n_9945),
.Y(n_12935)
);

OAI22xp33_ASAP7_75t_L g12936 ( 
.A1(n_11189),
.A2(n_10731),
.B1(n_10916),
.B2(n_9022),
.Y(n_12936)
);

OA21x2_ASAP7_75t_L g12937 ( 
.A1(n_11467),
.A2(n_9669),
.B(n_9668),
.Y(n_12937)
);

HB1xp67_ASAP7_75t_L g12938 ( 
.A(n_11639),
.Y(n_12938)
);

NAND2x1_ASAP7_75t_L g12939 ( 
.A(n_12191),
.B(n_10327),
.Y(n_12939)
);

NAND2xp5_ASAP7_75t_L g12940 ( 
.A(n_12051),
.B(n_9136),
.Y(n_12940)
);

AOI22xp5_ASAP7_75t_L g12941 ( 
.A1(n_11654),
.A2(n_10027),
.B1(n_9073),
.B2(n_8582),
.Y(n_12941)
);

OAI22xp33_ASAP7_75t_L g12942 ( 
.A1(n_11189),
.A2(n_10731),
.B1(n_10916),
.B2(n_9022),
.Y(n_12942)
);

AOI22xp33_ASAP7_75t_L g12943 ( 
.A1(n_12156),
.A2(n_10118),
.B1(n_10122),
.B2(n_10111),
.Y(n_12943)
);

AOI22xp5_ASAP7_75t_L g12944 ( 
.A1(n_12190),
.A2(n_10027),
.B1(n_9073),
.B2(n_8554),
.Y(n_12944)
);

AOI21xp33_ASAP7_75t_L g12945 ( 
.A1(n_12176),
.A2(n_9918),
.B(n_9911),
.Y(n_12945)
);

AOI22xp33_ASAP7_75t_SL g12946 ( 
.A1(n_11417),
.A2(n_10118),
.B1(n_10122),
.B2(n_10111),
.Y(n_12946)
);

BUFx5_ASAP7_75t_L g12947 ( 
.A(n_11216),
.Y(n_12947)
);

AOI22xp33_ASAP7_75t_L g12948 ( 
.A1(n_12158),
.A2(n_10128),
.B1(n_10132),
.B2(n_10124),
.Y(n_12948)
);

A2O1A1Ixp33_ASAP7_75t_L g12949 ( 
.A1(n_11214),
.A2(n_9120),
.B(n_9961),
.C(n_9957),
.Y(n_12949)
);

AOI22xp5_ASAP7_75t_L g12950 ( 
.A1(n_12215),
.A2(n_8554),
.B1(n_10175),
.B2(n_10151),
.Y(n_12950)
);

AO31x2_ASAP7_75t_L g12951 ( 
.A1(n_11765),
.A2(n_9961),
.A3(n_9971),
.B(n_9957),
.Y(n_12951)
);

OAI22xp33_ASAP7_75t_L g12952 ( 
.A1(n_11187),
.A2(n_10731),
.B1(n_10916),
.B2(n_9494),
.Y(n_12952)
);

CKINVDCx5p33_ASAP7_75t_R g12953 ( 
.A(n_11274),
.Y(n_12953)
);

NAND2xp5_ASAP7_75t_L g12954 ( 
.A(n_12058),
.B(n_9136),
.Y(n_12954)
);

AOI222xp33_ASAP7_75t_L g12955 ( 
.A1(n_11765),
.A2(n_10138),
.B1(n_10128),
.B2(n_10140),
.C1(n_10132),
.C2(n_10124),
.Y(n_12955)
);

INVx1_ASAP7_75t_L g12956 ( 
.A(n_11108),
.Y(n_12956)
);

OAI22xp33_ASAP7_75t_L g12957 ( 
.A1(n_11187),
.A2(n_10731),
.B1(n_10916),
.B2(n_9494),
.Y(n_12957)
);

OAI21xp5_ASAP7_75t_L g12958 ( 
.A1(n_11097),
.A2(n_11362),
.B(n_11241),
.Y(n_12958)
);

AOI22xp5_ASAP7_75t_L g12959 ( 
.A1(n_11767),
.A2(n_10191),
.B1(n_8815),
.B2(n_9976),
.Y(n_12959)
);

OAI22xp33_ASAP7_75t_L g12960 ( 
.A1(n_11298),
.A2(n_9515),
.B1(n_9255),
.B2(n_9239),
.Y(n_12960)
);

AND2x2_ASAP7_75t_L g12961 ( 
.A(n_12094),
.B(n_9945),
.Y(n_12961)
);

OR2x6_ASAP7_75t_L g12962 ( 
.A(n_11194),
.B(n_11198),
.Y(n_12962)
);

AOI221xp5_ASAP7_75t_L g12963 ( 
.A1(n_11767),
.A2(n_9976),
.B1(n_9987),
.B2(n_9980),
.C(n_9971),
.Y(n_12963)
);

OAI211xp5_ASAP7_75t_L g12964 ( 
.A1(n_12123),
.A2(n_9866),
.B(n_9881),
.C(n_9872),
.Y(n_12964)
);

OAI21x1_ASAP7_75t_L g12965 ( 
.A1(n_11241),
.A2(n_10694),
.B(n_10632),
.Y(n_12965)
);

AOI22xp33_ASAP7_75t_L g12966 ( 
.A1(n_12158),
.A2(n_10132),
.B1(n_10138),
.B2(n_10128),
.Y(n_12966)
);

INVx1_ASAP7_75t_L g12967 ( 
.A(n_11110),
.Y(n_12967)
);

INVx3_ASAP7_75t_L g12968 ( 
.A(n_11515),
.Y(n_12968)
);

INVx1_ASAP7_75t_SL g12969 ( 
.A(n_11384),
.Y(n_12969)
);

AOI22xp33_ASAP7_75t_L g12970 ( 
.A1(n_12167),
.A2(n_10140),
.B1(n_10141),
.B2(n_10138),
.Y(n_12970)
);

BUFx2_ASAP7_75t_L g12971 ( 
.A(n_12204),
.Y(n_12971)
);

NAND2xp5_ASAP7_75t_L g12972 ( 
.A(n_12058),
.B(n_12115),
.Y(n_12972)
);

AOI22xp33_ASAP7_75t_L g12973 ( 
.A1(n_12167),
.A2(n_10141),
.B1(n_10163),
.B2(n_10140),
.Y(n_12973)
);

AND2x2_ASAP7_75t_L g12974 ( 
.A(n_12123),
.B(n_10769),
.Y(n_12974)
);

AOI22xp33_ASAP7_75t_L g12975 ( 
.A1(n_12180),
.A2(n_10163),
.B1(n_10170),
.B2(n_10141),
.Y(n_12975)
);

OAI211xp5_ASAP7_75t_L g12976 ( 
.A1(n_11877),
.A2(n_9881),
.B(n_8302),
.C(n_10139),
.Y(n_12976)
);

AOI211xp5_ASAP7_75t_L g12977 ( 
.A1(n_11396),
.A2(n_8580),
.B(n_8463),
.C(n_8534),
.Y(n_12977)
);

AND2x2_ASAP7_75t_L g12978 ( 
.A(n_11137),
.B(n_10769),
.Y(n_12978)
);

HB1xp67_ASAP7_75t_L g12979 ( 
.A(n_11639),
.Y(n_12979)
);

INVx2_ASAP7_75t_L g12980 ( 
.A(n_12007),
.Y(n_12980)
);

INVx2_ASAP7_75t_L g12981 ( 
.A(n_12007),
.Y(n_12981)
);

BUFx2_ASAP7_75t_L g12982 ( 
.A(n_11306),
.Y(n_12982)
);

AOI22xp33_ASAP7_75t_L g12983 ( 
.A1(n_12180),
.A2(n_10170),
.B1(n_10182),
.B2(n_10163),
.Y(n_12983)
);

NAND2xp5_ASAP7_75t_L g12984 ( 
.A(n_12115),
.B(n_9136),
.Y(n_12984)
);

OAI22xp5_ASAP7_75t_SL g12985 ( 
.A1(n_11784),
.A2(n_7549),
.B1(n_7564),
.B2(n_7382),
.Y(n_12985)
);

OAI21x1_ASAP7_75t_L g12986 ( 
.A1(n_11889),
.A2(n_10694),
.B(n_10632),
.Y(n_12986)
);

OR2x2_ASAP7_75t_L g12987 ( 
.A(n_12202),
.B(n_9079),
.Y(n_12987)
);

INVx2_ASAP7_75t_L g12988 ( 
.A(n_12153),
.Y(n_12988)
);

OA21x2_ASAP7_75t_L g12989 ( 
.A1(n_11467),
.A2(n_9675),
.B(n_9668),
.Y(n_12989)
);

AOI221xp5_ASAP7_75t_L g12990 ( 
.A1(n_12189),
.A2(n_9976),
.B1(n_9987),
.B2(n_9980),
.C(n_9971),
.Y(n_12990)
);

BUFx3_ASAP7_75t_L g12991 ( 
.A(n_11921),
.Y(n_12991)
);

AOI22xp33_ASAP7_75t_L g12992 ( 
.A1(n_12189),
.A2(n_10182),
.B1(n_10193),
.B2(n_10170),
.Y(n_12992)
);

AO222x2_ASAP7_75t_L g12993 ( 
.A1(n_11950),
.A2(n_9757),
.B1(n_8652),
.B2(n_8419),
.C1(n_10065),
.C2(n_10017),
.Y(n_12993)
);

OAI211xp5_ASAP7_75t_L g12994 ( 
.A1(n_11877),
.A2(n_8302),
.B(n_10139),
.C(n_8833),
.Y(n_12994)
);

AO31x2_ASAP7_75t_L g12995 ( 
.A1(n_11967),
.A2(n_9987),
.A3(n_9980),
.B(n_10182),
.Y(n_12995)
);

OAI22xp5_ASAP7_75t_L g12996 ( 
.A1(n_12241),
.A2(n_8815),
.B1(n_9757),
.B2(n_10899),
.Y(n_12996)
);

OAI22xp5_ASAP7_75t_L g12997 ( 
.A1(n_11483),
.A2(n_10954),
.B1(n_8824),
.B2(n_9846),
.Y(n_12997)
);

AOI321xp33_ASAP7_75t_L g12998 ( 
.A1(n_11084),
.A2(n_10211),
.A3(n_10201),
.B1(n_10212),
.B2(n_10203),
.C(n_10193),
.Y(n_12998)
);

INVx3_ASAP7_75t_L g12999 ( 
.A(n_11515),
.Y(n_12999)
);

AND2x2_ASAP7_75t_L g13000 ( 
.A(n_11176),
.B(n_11190),
.Y(n_13000)
);

OR2x2_ASAP7_75t_L g13001 ( 
.A(n_11528),
.B(n_9079),
.Y(n_13001)
);

AOI22xp33_ASAP7_75t_L g13002 ( 
.A1(n_12192),
.A2(n_12201),
.B1(n_12205),
.B2(n_12195),
.Y(n_13002)
);

NAND2xp5_ASAP7_75t_L g13003 ( 
.A(n_12155),
.B(n_9205),
.Y(n_13003)
);

AOI22xp33_ASAP7_75t_L g13004 ( 
.A1(n_12192),
.A2(n_10201),
.B1(n_10203),
.B2(n_10193),
.Y(n_13004)
);

AOI221xp5_ASAP7_75t_L g13005 ( 
.A1(n_12195),
.A2(n_10203),
.B1(n_10212),
.B2(n_10211),
.C(n_10201),
.Y(n_13005)
);

OR2x2_ASAP7_75t_L g13006 ( 
.A(n_11893),
.B(n_9079),
.Y(n_13006)
);

OAI221xp5_ASAP7_75t_SL g13007 ( 
.A1(n_11084),
.A2(n_10212),
.B1(n_10235),
.B2(n_10228),
.C(n_10211),
.Y(n_13007)
);

AOI21xp33_ASAP7_75t_L g13008 ( 
.A1(n_12176),
.A2(n_9918),
.B(n_9911),
.Y(n_13008)
);

OAI22xp5_ASAP7_75t_L g13009 ( 
.A1(n_11950),
.A2(n_9841),
.B1(n_9886),
.B2(n_9846),
.Y(n_13009)
);

INVx3_ASAP7_75t_L g13010 ( 
.A(n_11586),
.Y(n_13010)
);

INVx2_ASAP7_75t_L g13011 ( 
.A(n_12153),
.Y(n_13011)
);

INVx1_ASAP7_75t_L g13012 ( 
.A(n_11111),
.Y(n_13012)
);

OAI22xp5_ASAP7_75t_L g13013 ( 
.A1(n_11950),
.A2(n_9841),
.B1(n_9886),
.B2(n_9846),
.Y(n_13013)
);

AOI21xp5_ASAP7_75t_L g13014 ( 
.A1(n_11182),
.A2(n_10611),
.B(n_10504),
.Y(n_13014)
);

AOI22xp33_ASAP7_75t_L g13015 ( 
.A1(n_12201),
.A2(n_10235),
.B1(n_10228),
.B2(n_9595),
.Y(n_13015)
);

INVx1_ASAP7_75t_L g13016 ( 
.A(n_11117),
.Y(n_13016)
);

OAI211xp5_ASAP7_75t_L g13017 ( 
.A1(n_11942),
.A2(n_10139),
.B(n_8833),
.C(n_9956),
.Y(n_13017)
);

NOR2xp33_ASAP7_75t_L g13018 ( 
.A(n_11683),
.B(n_9891),
.Y(n_13018)
);

AND2x2_ASAP7_75t_L g13019 ( 
.A(n_11190),
.B(n_9783),
.Y(n_13019)
);

OAI22xp5_ASAP7_75t_L g13020 ( 
.A1(n_11317),
.A2(n_9886),
.B1(n_9900),
.B2(n_9887),
.Y(n_13020)
);

INVx2_ASAP7_75t_L g13021 ( 
.A(n_12153),
.Y(n_13021)
);

OR2x6_ASAP7_75t_L g13022 ( 
.A(n_11194),
.B(n_7382),
.Y(n_13022)
);

OAI22xp33_ASAP7_75t_L g13023 ( 
.A1(n_11375),
.A2(n_9515),
.B1(n_9255),
.B2(n_9239),
.Y(n_13023)
);

INVx1_ASAP7_75t_L g13024 ( 
.A(n_11119),
.Y(n_13024)
);

AOI22xp33_ASAP7_75t_L g13025 ( 
.A1(n_12205),
.A2(n_10235),
.B1(n_10228),
.B2(n_9595),
.Y(n_13025)
);

AOI22xp33_ASAP7_75t_L g13026 ( 
.A1(n_12213),
.A2(n_9595),
.B1(n_9602),
.B2(n_9594),
.Y(n_13026)
);

OAI211xp5_ASAP7_75t_L g13027 ( 
.A1(n_11942),
.A2(n_10139),
.B(n_9916),
.C(n_9675),
.Y(n_13027)
);

INVx2_ASAP7_75t_SL g13028 ( 
.A(n_11784),
.Y(n_13028)
);

A2O1A1Ixp33_ASAP7_75t_L g13029 ( 
.A1(n_11396),
.A2(n_9120),
.B(n_8658),
.C(n_8707),
.Y(n_13029)
);

OAI222xp33_ASAP7_75t_L g13030 ( 
.A1(n_11324),
.A2(n_10530),
.B1(n_10547),
.B2(n_10406),
.C1(n_10380),
.C2(n_10310),
.Y(n_13030)
);

AOI221xp5_ASAP7_75t_L g13031 ( 
.A1(n_12213),
.A2(n_8580),
.B1(n_9602),
.B2(n_9604),
.C(n_9594),
.Y(n_13031)
);

OAI22xp33_ASAP7_75t_L g13032 ( 
.A1(n_11375),
.A2(n_9515),
.B1(n_10615),
.B2(n_10544),
.Y(n_13032)
);

NAND2xp5_ASAP7_75t_L g13033 ( 
.A(n_12155),
.B(n_9205),
.Y(n_13033)
);

AOI22xp33_ASAP7_75t_L g13034 ( 
.A1(n_12027),
.A2(n_9602),
.B1(n_9604),
.B2(n_9594),
.Y(n_13034)
);

BUFx2_ASAP7_75t_L g13035 ( 
.A(n_11306),
.Y(n_13035)
);

AOI221xp5_ASAP7_75t_L g13036 ( 
.A1(n_11589),
.A2(n_11624),
.B1(n_11651),
.B2(n_11615),
.C(n_11614),
.Y(n_13036)
);

OR2x2_ASAP7_75t_L g13037 ( 
.A(n_11122),
.B(n_9079),
.Y(n_13037)
);

INVx2_ASAP7_75t_L g13038 ( 
.A(n_12153),
.Y(n_13038)
);

OAI22xp33_ASAP7_75t_L g13039 ( 
.A1(n_11386),
.A2(n_10615),
.B1(n_10544),
.B2(n_8401),
.Y(n_13039)
);

INVx3_ASAP7_75t_L g13040 ( 
.A(n_11586),
.Y(n_13040)
);

INVx2_ASAP7_75t_L g13041 ( 
.A(n_11386),
.Y(n_13041)
);

NAND2xp5_ASAP7_75t_SL g13042 ( 
.A(n_11586),
.B(n_9911),
.Y(n_13042)
);

INVx1_ASAP7_75t_L g13043 ( 
.A(n_11126),
.Y(n_13043)
);

OAI211xp5_ASAP7_75t_L g13044 ( 
.A1(n_12032),
.A2(n_10318),
.B(n_10324),
.C(n_10269),
.Y(n_13044)
);

AND2x4_ASAP7_75t_SL g13045 ( 
.A(n_11198),
.B(n_10750),
.Y(n_13045)
);

AOI22xp33_ASAP7_75t_L g13046 ( 
.A1(n_11967),
.A2(n_9627),
.B1(n_9629),
.B2(n_9604),
.Y(n_13046)
);

AOI22xp5_ASAP7_75t_L g13047 ( 
.A1(n_11324),
.A2(n_9098),
.B1(n_9982),
.B2(n_9909),
.Y(n_13047)
);

OAI21xp33_ASAP7_75t_L g13048 ( 
.A1(n_12223),
.A2(n_9597),
.B(n_9904),
.Y(n_13048)
);

AND2x2_ASAP7_75t_L g13049 ( 
.A(n_11295),
.B(n_9783),
.Y(n_13049)
);

OR2x2_ASAP7_75t_L g13050 ( 
.A(n_11128),
.B(n_9079),
.Y(n_13050)
);

BUFx8_ASAP7_75t_SL g13051 ( 
.A(n_11052),
.Y(n_13051)
);

AOI22xp33_ASAP7_75t_L g13052 ( 
.A1(n_12027),
.A2(n_9629),
.B1(n_9635),
.B2(n_9627),
.Y(n_13052)
);

OAI22xp33_ASAP7_75t_L g13053 ( 
.A1(n_12221),
.A2(n_10615),
.B1(n_10544),
.B2(n_8401),
.Y(n_13053)
);

AOI22xp33_ASAP7_75t_L g13054 ( 
.A1(n_12076),
.A2(n_9629),
.B1(n_9635),
.B2(n_9627),
.Y(n_13054)
);

INVx2_ASAP7_75t_L g13055 ( 
.A(n_11088),
.Y(n_13055)
);

AOI21xp33_ASAP7_75t_L g13056 ( 
.A1(n_12223),
.A2(n_12253),
.B(n_11089),
.Y(n_13056)
);

AND2x4_ASAP7_75t_L g13057 ( 
.A(n_11996),
.B(n_9887),
.Y(n_13057)
);

AOI22xp33_ASAP7_75t_L g13058 ( 
.A1(n_12076),
.A2(n_9642),
.B1(n_9653),
.B2(n_9635),
.Y(n_13058)
);

AOI222xp33_ASAP7_75t_L g13059 ( 
.A1(n_11589),
.A2(n_8926),
.B1(n_8907),
.B2(n_9642),
.C1(n_9663),
.C2(n_9653),
.Y(n_13059)
);

OR2x2_ASAP7_75t_L g13060 ( 
.A(n_11134),
.B(n_9205),
.Y(n_13060)
);

INVx1_ASAP7_75t_L g13061 ( 
.A(n_11136),
.Y(n_13061)
);

INVx1_ASAP7_75t_L g13062 ( 
.A(n_11141),
.Y(n_13062)
);

AND2x2_ASAP7_75t_L g13063 ( 
.A(n_11295),
.B(n_9783),
.Y(n_13063)
);

AOI221xp5_ASAP7_75t_L g13064 ( 
.A1(n_11614),
.A2(n_9663),
.B1(n_9678),
.B2(n_9653),
.C(n_9642),
.Y(n_13064)
);

OR2x2_ASAP7_75t_L g13065 ( 
.A(n_11142),
.B(n_9205),
.Y(n_13065)
);

AOI22xp33_ASAP7_75t_L g13066 ( 
.A1(n_11993),
.A2(n_9678),
.B1(n_9679),
.B2(n_9663),
.Y(n_13066)
);

AOI22xp33_ASAP7_75t_L g13067 ( 
.A1(n_11993),
.A2(n_9679),
.B1(n_9685),
.B2(n_9678),
.Y(n_13067)
);

NAND2xp5_ASAP7_75t_SL g13068 ( 
.A(n_11324),
.B(n_9911),
.Y(n_13068)
);

NOR2x1_ASAP7_75t_SL g13069 ( 
.A(n_11249),
.B(n_10434),
.Y(n_13069)
);

OA21x2_ASAP7_75t_L g13070 ( 
.A1(n_11502),
.A2(n_9693),
.B(n_10121),
.Y(n_13070)
);

OA21x2_ASAP7_75t_L g13071 ( 
.A1(n_11502),
.A2(n_9693),
.B(n_10121),
.Y(n_13071)
);

AOI21xp5_ASAP7_75t_SL g13072 ( 
.A1(n_11249),
.A2(n_10293),
.B(n_10453),
.Y(n_13072)
);

AND2x2_ASAP7_75t_L g13073 ( 
.A(n_11363),
.B(n_9783),
.Y(n_13073)
);

INVx1_ASAP7_75t_L g13074 ( 
.A(n_11145),
.Y(n_13074)
);

AOI221xp5_ASAP7_75t_L g13075 ( 
.A1(n_11615),
.A2(n_9700),
.B1(n_9704),
.B2(n_9685),
.C(n_9679),
.Y(n_13075)
);

AOI22xp33_ASAP7_75t_L g13076 ( 
.A1(n_12050),
.A2(n_9700),
.B1(n_9704),
.B2(n_9685),
.Y(n_13076)
);

AOI21xp5_ASAP7_75t_SL g13077 ( 
.A1(n_11459),
.A2(n_10293),
.B(n_10309),
.Y(n_13077)
);

OAI21x1_ASAP7_75t_L g13078 ( 
.A1(n_11889),
.A2(n_10784),
.B(n_10761),
.Y(n_13078)
);

OAI221xp5_ASAP7_75t_L g13079 ( 
.A1(n_12253),
.A2(n_10758),
.B1(n_9712),
.B2(n_9725),
.C(n_9704),
.Y(n_13079)
);

BUFx6f_ASAP7_75t_L g13080 ( 
.A(n_11198),
.Y(n_13080)
);

AND2x4_ASAP7_75t_L g13081 ( 
.A(n_11996),
.B(n_9887),
.Y(n_13081)
);

OAI221xp5_ASAP7_75t_L g13082 ( 
.A1(n_11690),
.A2(n_9725),
.B1(n_9731),
.B2(n_9712),
.C(n_9700),
.Y(n_13082)
);

INVx1_ASAP7_75t_L g13083 ( 
.A(n_11149),
.Y(n_13083)
);

AOI222xp33_ASAP7_75t_L g13084 ( 
.A1(n_11624),
.A2(n_8926),
.B1(n_8907),
.B2(n_9712),
.C1(n_9731),
.C2(n_9725),
.Y(n_13084)
);

AOI22xp33_ASAP7_75t_L g13085 ( 
.A1(n_12077),
.A2(n_9737),
.B1(n_9751),
.B2(n_9731),
.Y(n_13085)
);

OAI22xp5_ASAP7_75t_L g13086 ( 
.A1(n_11233),
.A2(n_9900),
.B1(n_9346),
.B2(n_9283),
.Y(n_13086)
);

AND2x4_ASAP7_75t_L g13087 ( 
.A(n_11996),
.B(n_9900),
.Y(n_13087)
);

OAI22xp5_ASAP7_75t_L g13088 ( 
.A1(n_11279),
.A2(n_9346),
.B1(n_9283),
.B2(n_10476),
.Y(n_13088)
);

NAND3xp33_ASAP7_75t_L g13089 ( 
.A(n_12166),
.B(n_9918),
.C(n_9911),
.Y(n_13089)
);

AOI22xp33_ASAP7_75t_SL g13090 ( 
.A1(n_11362),
.A2(n_9751),
.B1(n_9755),
.B2(n_9737),
.Y(n_13090)
);

OAI22xp5_ASAP7_75t_L g13091 ( 
.A1(n_11335),
.A2(n_10476),
.B1(n_10551),
.B2(n_10525),
.Y(n_13091)
);

AOI22xp5_ASAP7_75t_L g13092 ( 
.A1(n_11409),
.A2(n_9098),
.B1(n_9982),
.B2(n_9909),
.Y(n_13092)
);

AOI21xp5_ASAP7_75t_L g13093 ( 
.A1(n_12161),
.A2(n_10611),
.B(n_10504),
.Y(n_13093)
);

OR2x6_ASAP7_75t_L g13094 ( 
.A(n_11198),
.B(n_7549),
.Y(n_13094)
);

INVx1_ASAP7_75t_L g13095 ( 
.A(n_11153),
.Y(n_13095)
);

INVx4_ASAP7_75t_L g13096 ( 
.A(n_11054),
.Y(n_13096)
);

OAI211xp5_ASAP7_75t_L g13097 ( 
.A1(n_11942),
.A2(n_10498),
.B(n_10500),
.C(n_10438),
.Y(n_13097)
);

OAI221xp5_ASAP7_75t_SL g13098 ( 
.A1(n_11088),
.A2(n_8865),
.B1(n_8832),
.B2(n_8687),
.C(n_9737),
.Y(n_13098)
);

NAND2xp5_ASAP7_75t_L g13099 ( 
.A(n_11639),
.B(n_9205),
.Y(n_13099)
);

AOI22xp33_ASAP7_75t_L g13100 ( 
.A1(n_12042),
.A2(n_9755),
.B1(n_9768),
.B2(n_9751),
.Y(n_13100)
);

INVx2_ASAP7_75t_L g13101 ( 
.A(n_11089),
.Y(n_13101)
);

INVx4_ASAP7_75t_L g13102 ( 
.A(n_11054),
.Y(n_13102)
);

INVx2_ASAP7_75t_L g13103 ( 
.A(n_11098),
.Y(n_13103)
);

OR2x2_ASAP7_75t_L g13104 ( 
.A(n_11157),
.B(n_9205),
.Y(n_13104)
);

AOI22xp33_ASAP7_75t_L g13105 ( 
.A1(n_12023),
.A2(n_11988),
.B1(n_11998),
.B2(n_11985),
.Y(n_13105)
);

AOI221xp5_ASAP7_75t_L g13106 ( 
.A1(n_11651),
.A2(n_9777),
.B1(n_9779),
.B2(n_9768),
.C(n_9755),
.Y(n_13106)
);

A2O1A1Ixp33_ASAP7_75t_L g13107 ( 
.A1(n_11733),
.A2(n_9120),
.B(n_8658),
.C(n_8707),
.Y(n_13107)
);

AOI22xp33_ASAP7_75t_L g13108 ( 
.A1(n_11988),
.A2(n_9777),
.B1(n_9779),
.B2(n_9768),
.Y(n_13108)
);

INVx2_ASAP7_75t_L g13109 ( 
.A(n_11098),
.Y(n_13109)
);

AOI22xp33_ASAP7_75t_SL g13110 ( 
.A1(n_11569),
.A2(n_9779),
.B1(n_9777),
.B2(n_9991),
.Y(n_13110)
);

NAND3xp33_ASAP7_75t_L g13111 ( 
.A(n_12166),
.B(n_10137),
.C(n_10061),
.Y(n_13111)
);

OAI22xp33_ASAP7_75t_L g13112 ( 
.A1(n_12221),
.A2(n_10615),
.B1(n_10544),
.B2(n_8401),
.Y(n_13112)
);

AOI22xp33_ASAP7_75t_L g13113 ( 
.A1(n_12075),
.A2(n_11998),
.B1(n_12003),
.B2(n_11985),
.Y(n_13113)
);

AO31x2_ASAP7_75t_L g13114 ( 
.A1(n_12003),
.A2(n_10083),
.A3(n_9721),
.B(n_10652),
.Y(n_13114)
);

AOI222xp33_ASAP7_75t_L g13115 ( 
.A1(n_11667),
.A2(n_8939),
.B1(n_9154),
.B2(n_9164),
.C1(n_9102),
.C2(n_9095),
.Y(n_13115)
);

INVx2_ASAP7_75t_L g13116 ( 
.A(n_11100),
.Y(n_13116)
);

AND2x2_ASAP7_75t_L g13117 ( 
.A(n_11363),
.B(n_9783),
.Y(n_13117)
);

OR2x2_ASAP7_75t_L g13118 ( 
.A(n_11169),
.B(n_9205),
.Y(n_13118)
);

AOI22xp33_ASAP7_75t_L g13119 ( 
.A1(n_12023),
.A2(n_10137),
.B1(n_10152),
.B2(n_10061),
.Y(n_13119)
);

OAI22xp5_ASAP7_75t_L g13120 ( 
.A1(n_11342),
.A2(n_10476),
.B1(n_10551),
.B2(n_10525),
.Y(n_13120)
);

INVx1_ASAP7_75t_L g13121 ( 
.A(n_11170),
.Y(n_13121)
);

CKINVDCx6p67_ASAP7_75t_R g13122 ( 
.A(n_11047),
.Y(n_13122)
);

NAND2xp5_ASAP7_75t_L g13123 ( 
.A(n_11639),
.B(n_9205),
.Y(n_13123)
);

AOI22xp33_ASAP7_75t_L g13124 ( 
.A1(n_12077),
.A2(n_10137),
.B1(n_10152),
.B2(n_10061),
.Y(n_13124)
);

AOI22xp33_ASAP7_75t_L g13125 ( 
.A1(n_12042),
.A2(n_10137),
.B1(n_10152),
.B2(n_10061),
.Y(n_13125)
);

INVx2_ASAP7_75t_L g13126 ( 
.A(n_11100),
.Y(n_13126)
);

BUFx4f_ASAP7_75t_SL g13127 ( 
.A(n_11047),
.Y(n_13127)
);

NOR2xp33_ASAP7_75t_L g13128 ( 
.A(n_11683),
.B(n_9641),
.Y(n_13128)
);

AOI22xp33_ASAP7_75t_L g13129 ( 
.A1(n_12069),
.A2(n_10137),
.B1(n_10152),
.B2(n_10061),
.Y(n_13129)
);

AND2x6_ASAP7_75t_L g13130 ( 
.A(n_11580),
.B(n_10309),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_11171),
.Y(n_13131)
);

OAI22xp33_ASAP7_75t_L g13132 ( 
.A1(n_12232),
.A2(n_10615),
.B1(n_10544),
.B2(n_8401),
.Y(n_13132)
);

NAND2xp5_ASAP7_75t_L g13133 ( 
.A(n_11744),
.B(n_9164),
.Y(n_13133)
);

A2O1A1Ixp33_ASAP7_75t_L g13134 ( 
.A1(n_11733),
.A2(n_9095),
.B(n_9102),
.C(n_8528),
.Y(n_13134)
);

AND2x2_ASAP7_75t_L g13135 ( 
.A(n_11399),
.B(n_10525),
.Y(n_13135)
);

AOI22xp5_ASAP7_75t_L g13136 ( 
.A1(n_11409),
.A2(n_10195),
.B1(n_9180),
.B2(n_10739),
.Y(n_13136)
);

AOI22xp33_ASAP7_75t_L g13137 ( 
.A1(n_12050),
.A2(n_10137),
.B1(n_10152),
.B2(n_10061),
.Y(n_13137)
);

AOI221xp5_ASAP7_75t_L g13138 ( 
.A1(n_11667),
.A2(n_10988),
.B1(n_11002),
.B2(n_10986),
.C(n_10967),
.Y(n_13138)
);

AND2x2_ASAP7_75t_L g13139 ( 
.A(n_11399),
.B(n_10551),
.Y(n_13139)
);

AOI22xp33_ASAP7_75t_SL g13140 ( 
.A1(n_11569),
.A2(n_9991),
.B1(n_9827),
.B2(n_10512),
.Y(n_13140)
);

OAI221xp5_ASAP7_75t_L g13141 ( 
.A1(n_11690),
.A2(n_9991),
.B1(n_10834),
.B2(n_10831),
.C(n_10633),
.Y(n_13141)
);

AOI22xp33_ASAP7_75t_L g13142 ( 
.A1(n_12069),
.A2(n_10216),
.B1(n_10222),
.B2(n_10152),
.Y(n_13142)
);

NAND2xp5_ASAP7_75t_L g13143 ( 
.A(n_11744),
.B(n_10195),
.Y(n_13143)
);

AOI22xp33_ASAP7_75t_SL g13144 ( 
.A1(n_11605),
.A2(n_9991),
.B1(n_9827),
.B2(n_10512),
.Y(n_13144)
);

O2A1O1Ixp5_ASAP7_75t_L g13145 ( 
.A1(n_11426),
.A2(n_11473),
.B(n_11520),
.C(n_11449),
.Y(n_13145)
);

OAI22xp5_ASAP7_75t_L g13146 ( 
.A1(n_12232),
.A2(n_10572),
.B1(n_10606),
.B2(n_10593),
.Y(n_13146)
);

OAI22xp5_ASAP7_75t_L g13147 ( 
.A1(n_11784),
.A2(n_10572),
.B1(n_10606),
.B2(n_10593),
.Y(n_13147)
);

OAI211xp5_ASAP7_75t_SL g13148 ( 
.A1(n_11604),
.A2(n_10510),
.B(n_9645),
.C(n_9694),
.Y(n_13148)
);

AOI221xp5_ASAP7_75t_L g13149 ( 
.A1(n_11109),
.A2(n_10988),
.B1(n_11002),
.B2(n_10986),
.C(n_10967),
.Y(n_13149)
);

OAI22xp5_ASAP7_75t_L g13150 ( 
.A1(n_11969),
.A2(n_10572),
.B1(n_10606),
.B2(n_10593),
.Y(n_13150)
);

NOR2x1_ASAP7_75t_L g13151 ( 
.A(n_11751),
.B(n_9641),
.Y(n_13151)
);

INVx3_ASAP7_75t_L g13152 ( 
.A(n_11409),
.Y(n_13152)
);

AND2x2_ASAP7_75t_L g13153 ( 
.A(n_11798),
.B(n_10313),
.Y(n_13153)
);

INVx1_ASAP7_75t_L g13154 ( 
.A(n_11174),
.Y(n_13154)
);

OAI22xp5_ASAP7_75t_L g13155 ( 
.A1(n_11969),
.A2(n_9180),
.B1(n_10365),
.B2(n_10313),
.Y(n_13155)
);

OAI21xp5_ASAP7_75t_L g13156 ( 
.A1(n_11699),
.A2(n_8520),
.B(n_8313),
.Y(n_13156)
);

AOI21xp5_ASAP7_75t_L g13157 ( 
.A1(n_12161),
.A2(n_10611),
.B(n_10504),
.Y(n_13157)
);

BUFx3_ASAP7_75t_L g13158 ( 
.A(n_11130),
.Y(n_13158)
);

AND2x2_ASAP7_75t_L g13159 ( 
.A(n_11798),
.B(n_10313),
.Y(n_13159)
);

INVx1_ASAP7_75t_L g13160 ( 
.A(n_11177),
.Y(n_13160)
);

INVx2_ASAP7_75t_L g13161 ( 
.A(n_11109),
.Y(n_13161)
);

AOI22xp5_ASAP7_75t_L g13162 ( 
.A1(n_11427),
.A2(n_9180),
.B1(n_10746),
.B2(n_10293),
.Y(n_13162)
);

OAI22xp5_ASAP7_75t_L g13163 ( 
.A1(n_11969),
.A2(n_9180),
.B1(n_10365),
.B2(n_10313),
.Y(n_13163)
);

INVx3_ASAP7_75t_L g13164 ( 
.A(n_11427),
.Y(n_13164)
);

INVx3_ASAP7_75t_L g13165 ( 
.A(n_11427),
.Y(n_13165)
);

AOI221xp5_ASAP7_75t_L g13166 ( 
.A1(n_11112),
.A2(n_11118),
.B1(n_11125),
.B2(n_11116),
.C(n_11114),
.Y(n_13166)
);

OAI21xp5_ASAP7_75t_SL g13167 ( 
.A1(n_11717),
.A2(n_10930),
.B(n_10909),
.Y(n_13167)
);

OAI22xp5_ASAP7_75t_L g13168 ( 
.A1(n_11860),
.A2(n_10398),
.B1(n_10465),
.B2(n_10365),
.Y(n_13168)
);

OR2x2_ASAP7_75t_L g13169 ( 
.A(n_11184),
.B(n_9265),
.Y(n_13169)
);

AND2x2_ASAP7_75t_L g13170 ( 
.A(n_11860),
.B(n_10365),
.Y(n_13170)
);

NAND3xp33_ASAP7_75t_L g13171 ( 
.A(n_12166),
.B(n_10222),
.C(n_10216),
.Y(n_13171)
);

OAI21x1_ASAP7_75t_L g13172 ( 
.A1(n_11924),
.A2(n_10784),
.B(n_10761),
.Y(n_13172)
);

OAI22xp5_ASAP7_75t_L g13173 ( 
.A1(n_11945),
.A2(n_10465),
.B1(n_10482),
.B2(n_10398),
.Y(n_13173)
);

BUFx2_ASAP7_75t_L g13174 ( 
.A(n_11127),
.Y(n_13174)
);

BUFx4f_ASAP7_75t_SL g13175 ( 
.A(n_11130),
.Y(n_13175)
);

AOI21xp5_ASAP7_75t_L g13176 ( 
.A1(n_11605),
.A2(n_9694),
.B(n_9645),
.Y(n_13176)
);

AND2x2_ASAP7_75t_L g13177 ( 
.A(n_11945),
.B(n_10398),
.Y(n_13177)
);

AOI22xp33_ASAP7_75t_L g13178 ( 
.A1(n_12075),
.A2(n_12081),
.B1(n_10222),
.B2(n_10341),
.Y(n_13178)
);

AND2x2_ASAP7_75t_L g13179 ( 
.A(n_11361),
.B(n_10398),
.Y(n_13179)
);

INVx1_ASAP7_75t_L g13180 ( 
.A(n_11185),
.Y(n_13180)
);

AND2x2_ASAP7_75t_L g13181 ( 
.A(n_11549),
.B(n_10465),
.Y(n_13181)
);

CKINVDCx20_ASAP7_75t_R g13182 ( 
.A(n_11143),
.Y(n_13182)
);

NAND2xp5_ASAP7_75t_L g13183 ( 
.A(n_11222),
.B(n_8652),
.Y(n_13183)
);

OAI211xp5_ASAP7_75t_SL g13184 ( 
.A1(n_11604),
.A2(n_9729),
.B(n_9709),
.C(n_8865),
.Y(n_13184)
);

INVx3_ASAP7_75t_L g13185 ( 
.A(n_11456),
.Y(n_13185)
);

OR2x2_ASAP7_75t_L g13186 ( 
.A(n_11188),
.B(n_9265),
.Y(n_13186)
);

AND2x2_ASAP7_75t_L g13187 ( 
.A(n_11573),
.B(n_10465),
.Y(n_13187)
);

AOI22xp33_ASAP7_75t_L g13188 ( 
.A1(n_12081),
.A2(n_10222),
.B1(n_10341),
.B2(n_10216),
.Y(n_13188)
);

AOI21xp5_ASAP7_75t_L g13189 ( 
.A1(n_11643),
.A2(n_9729),
.B(n_9709),
.Y(n_13189)
);

AOI22xp33_ASAP7_75t_L g13190 ( 
.A1(n_11374),
.A2(n_10222),
.B1(n_10341),
.B2(n_10216),
.Y(n_13190)
);

AOI21xp5_ASAP7_75t_L g13191 ( 
.A1(n_11643),
.A2(n_9003),
.B(n_9410),
.Y(n_13191)
);

OAI22xp5_ASAP7_75t_L g13192 ( 
.A1(n_11456),
.A2(n_10506),
.B1(n_10707),
.B2(n_10482),
.Y(n_13192)
);

HB1xp67_ASAP7_75t_L g13193 ( 
.A(n_11191),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_11193),
.Y(n_13194)
);

OAI22xp5_ASAP7_75t_L g13195 ( 
.A1(n_11456),
.A2(n_10506),
.B1(n_10707),
.B2(n_10482),
.Y(n_13195)
);

INVx4_ASAP7_75t_L g13196 ( 
.A(n_11683),
.Y(n_13196)
);

INVx2_ASAP7_75t_L g13197 ( 
.A(n_11112),
.Y(n_13197)
);

A2O1A1Ixp33_ASAP7_75t_L g13198 ( 
.A1(n_11699),
.A2(n_9095),
.B(n_9102),
.C(n_9121),
.Y(n_13198)
);

AO21x2_ASAP7_75t_L g13199 ( 
.A1(n_11364),
.A2(n_10865),
.B(n_10787),
.Y(n_13199)
);

BUFx4f_ASAP7_75t_SL g13200 ( 
.A(n_11143),
.Y(n_13200)
);

OAI21x1_ASAP7_75t_L g13201 ( 
.A1(n_11924),
.A2(n_10992),
.B(n_10787),
.Y(n_13201)
);

NAND2xp5_ASAP7_75t_L g13202 ( 
.A(n_11222),
.B(n_8652),
.Y(n_13202)
);

INVx2_ASAP7_75t_L g13203 ( 
.A(n_11114),
.Y(n_13203)
);

INVx1_ASAP7_75t_L g13204 ( 
.A(n_11207),
.Y(n_13204)
);

NAND2xp5_ASAP7_75t_L g13205 ( 
.A(n_11222),
.B(n_8652),
.Y(n_13205)
);

INVx2_ASAP7_75t_L g13206 ( 
.A(n_11116),
.Y(n_13206)
);

OAI21x1_ASAP7_75t_L g13207 ( 
.A1(n_11929),
.A2(n_10995),
.B(n_10992),
.Y(n_13207)
);

OAI21x1_ASAP7_75t_L g13208 ( 
.A1(n_11929),
.A2(n_10995),
.B(n_10930),
.Y(n_13208)
);

AOI22xp5_ASAP7_75t_L g13209 ( 
.A1(n_11532),
.A2(n_8862),
.B1(n_8934),
.B2(n_9501),
.Y(n_13209)
);

OAI22xp5_ASAP7_75t_SL g13210 ( 
.A1(n_11374),
.A2(n_7549),
.B1(n_7722),
.B2(n_7564),
.Y(n_13210)
);

OAI22xp5_ASAP7_75t_L g13211 ( 
.A1(n_11532),
.A2(n_10506),
.B1(n_10707),
.B2(n_10482),
.Y(n_13211)
);

NOR2xp33_ASAP7_75t_L g13212 ( 
.A(n_11683),
.B(n_10817),
.Y(n_13212)
);

AOI21x1_ASAP7_75t_L g13213 ( 
.A1(n_11597),
.A2(n_9597),
.B(n_8386),
.Y(n_13213)
);

OR2x2_ASAP7_75t_L g13214 ( 
.A(n_11209),
.B(n_9265),
.Y(n_13214)
);

AOI22xp33_ASAP7_75t_L g13215 ( 
.A1(n_11401),
.A2(n_10222),
.B1(n_10341),
.B2(n_10216),
.Y(n_13215)
);

AOI221xp5_ASAP7_75t_SL g13216 ( 
.A1(n_11970),
.A2(n_9305),
.B1(n_8832),
.B2(n_9428),
.C(n_9400),
.Y(n_13216)
);

OAI211xp5_ASAP7_75t_L g13217 ( 
.A1(n_12032),
.A2(n_10341),
.B(n_10377),
.C(n_10216),
.Y(n_13217)
);

OR2x6_ASAP7_75t_L g13218 ( 
.A(n_11401),
.B(n_7549),
.Y(n_13218)
);

INVx2_ASAP7_75t_L g13219 ( 
.A(n_11118),
.Y(n_13219)
);

AND2x2_ASAP7_75t_L g13220 ( 
.A(n_11913),
.B(n_10506),
.Y(n_13220)
);

INVx1_ASAP7_75t_L g13221 ( 
.A(n_11210),
.Y(n_13221)
);

INVx3_ASAP7_75t_L g13222 ( 
.A(n_11532),
.Y(n_13222)
);

OA21x2_ASAP7_75t_L g13223 ( 
.A1(n_11364),
.A2(n_9693),
.B(n_10121),
.Y(n_13223)
);

OAI22xp5_ASAP7_75t_L g13224 ( 
.A1(n_11593),
.A2(n_10710),
.B1(n_10714),
.B2(n_10707),
.Y(n_13224)
);

OAI22xp5_ASAP7_75t_L g13225 ( 
.A1(n_11593),
.A2(n_10714),
.B1(n_10710),
.B2(n_10861),
.Y(n_13225)
);

INVx2_ASAP7_75t_L g13226 ( 
.A(n_11125),
.Y(n_13226)
);

HB1xp67_ASAP7_75t_L g13227 ( 
.A(n_11213),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_11927),
.B(n_10710),
.Y(n_13228)
);

OAI22xp5_ASAP7_75t_SL g13229 ( 
.A1(n_11410),
.A2(n_7564),
.B1(n_7777),
.B2(n_7722),
.Y(n_13229)
);

AOI22xp33_ASAP7_75t_SL g13230 ( 
.A1(n_11504),
.A2(n_9827),
.B1(n_10559),
.B2(n_10512),
.Y(n_13230)
);

OAI22xp5_ASAP7_75t_L g13231 ( 
.A1(n_11593),
.A2(n_10714),
.B1(n_10710),
.B2(n_10312),
.Y(n_13231)
);

AOI22xp5_ASAP7_75t_L g13232 ( 
.A1(n_11609),
.A2(n_8862),
.B1(n_8934),
.B2(n_9501),
.Y(n_13232)
);

INVx2_ASAP7_75t_L g13233 ( 
.A(n_11131),
.Y(n_13233)
);

AOI22xp33_ASAP7_75t_L g13234 ( 
.A1(n_11410),
.A2(n_10377),
.B1(n_10389),
.B2(n_10341),
.Y(n_13234)
);

INVxp33_ASAP7_75t_L g13235 ( 
.A(n_11970),
.Y(n_13235)
);

AOI221xp5_ASAP7_75t_L g13236 ( 
.A1(n_11131),
.A2(n_10988),
.B1(n_11002),
.B2(n_10986),
.C(n_10967),
.Y(n_13236)
);

OAI211xp5_ASAP7_75t_SL g13237 ( 
.A1(n_11612),
.A2(n_9305),
.B(n_9671),
.C(n_9664),
.Y(n_13237)
);

BUFx2_ASAP7_75t_L g13238 ( 
.A(n_11751),
.Y(n_13238)
);

AO21x1_ASAP7_75t_L g13239 ( 
.A1(n_11133),
.A2(n_10831),
.B(n_10633),
.Y(n_13239)
);

OAI211xp5_ASAP7_75t_L g13240 ( 
.A1(n_12064),
.A2(n_10389),
.B(n_10377),
.C(n_10312),
.Y(n_13240)
);

AOI22xp33_ASAP7_75t_L g13241 ( 
.A1(n_11452),
.A2(n_10389),
.B1(n_10377),
.B2(n_8903),
.Y(n_13241)
);

AOI22xp33_ASAP7_75t_SL g13242 ( 
.A1(n_11504),
.A2(n_9827),
.B1(n_10559),
.B2(n_10512),
.Y(n_13242)
);

OAI211xp5_ASAP7_75t_SL g13243 ( 
.A1(n_11612),
.A2(n_9671),
.B(n_9713),
.C(n_9664),
.Y(n_13243)
);

AOI22xp33_ASAP7_75t_L g13244 ( 
.A1(n_11452),
.A2(n_10389),
.B1(n_10377),
.B2(n_8903),
.Y(n_13244)
);

CKINVDCx16_ASAP7_75t_R g13245 ( 
.A(n_11154),
.Y(n_13245)
);

INVx1_ASAP7_75t_L g13246 ( 
.A(n_11220),
.Y(n_13246)
);

OAI22xp5_ASAP7_75t_L g13247 ( 
.A1(n_11609),
.A2(n_10714),
.B1(n_10312),
.B2(n_10320),
.Y(n_13247)
);

AND2x2_ASAP7_75t_L g13248 ( 
.A(n_11953),
.B(n_10377),
.Y(n_13248)
);

OR2x2_ASAP7_75t_L g13249 ( 
.A(n_11223),
.B(n_10048),
.Y(n_13249)
);

AOI22xp33_ASAP7_75t_L g13250 ( 
.A1(n_11460),
.A2(n_10389),
.B1(n_11659),
.B2(n_11625),
.Y(n_13250)
);

AOI21xp33_ASAP7_75t_L g13251 ( 
.A1(n_11133),
.A2(n_10389),
.B(n_10338),
.Y(n_13251)
);

CKINVDCx5p33_ASAP7_75t_R g13252 ( 
.A(n_11154),
.Y(n_13252)
);

AOI22xp33_ASAP7_75t_SL g13253 ( 
.A1(n_11843),
.A2(n_10559),
.B1(n_8456),
.B2(n_9656),
.Y(n_13253)
);

INVx2_ASAP7_75t_L g13254 ( 
.A(n_11144),
.Y(n_13254)
);

OAI21xp5_ASAP7_75t_SL g13255 ( 
.A1(n_11717),
.A2(n_10909),
.B(n_10582),
.Y(n_13255)
);

INVx4_ASAP7_75t_L g13256 ( 
.A(n_11970),
.Y(n_13256)
);

BUFx6f_ASAP7_75t_L g13257 ( 
.A(n_11156),
.Y(n_13257)
);

AOI222xp33_ASAP7_75t_L g13258 ( 
.A1(n_11144),
.A2(n_8939),
.B1(n_9386),
.B2(n_8737),
.C1(n_8589),
.C2(n_8765),
.Y(n_13258)
);

INVx1_ASAP7_75t_L g13259 ( 
.A(n_11224),
.Y(n_13259)
);

INVx2_ASAP7_75t_L g13260 ( 
.A(n_11158),
.Y(n_13260)
);

OAI22xp33_ASAP7_75t_L g13261 ( 
.A1(n_11163),
.A2(n_8401),
.B1(n_8955),
.B2(n_8232),
.Y(n_13261)
);

OAI221xp5_ASAP7_75t_L g13262 ( 
.A1(n_11690),
.A2(n_10834),
.B1(n_10863),
.B2(n_10831),
.C(n_10633),
.Y(n_13262)
);

AOI221xp5_ASAP7_75t_L g13263 ( 
.A1(n_11158),
.A2(n_11015),
.B1(n_11009),
.B2(n_10740),
.C(n_10749),
.Y(n_13263)
);

AOI21xp5_ASAP7_75t_L g13264 ( 
.A1(n_11986),
.A2(n_8792),
.B(n_8753),
.Y(n_13264)
);

OA21x2_ASAP7_75t_L g13265 ( 
.A1(n_11514),
.A2(n_10588),
.B(n_10502),
.Y(n_13265)
);

AOI22xp33_ASAP7_75t_L g13266 ( 
.A1(n_11460),
.A2(n_11659),
.B1(n_11625),
.B2(n_11164),
.Y(n_13266)
);

OAI221xp5_ASAP7_75t_L g13267 ( 
.A1(n_11870),
.A2(n_10893),
.B1(n_10906),
.B2(n_10863),
.C(n_10834),
.Y(n_13267)
);

INVx2_ASAP7_75t_L g13268 ( 
.A(n_11162),
.Y(n_13268)
);

INVx1_ASAP7_75t_L g13269 ( 
.A(n_11228),
.Y(n_13269)
);

INVx1_ASAP7_75t_L g13270 ( 
.A(n_11229),
.Y(n_13270)
);

OAI21xp5_ASAP7_75t_SL g13271 ( 
.A1(n_11095),
.A2(n_10582),
.B(n_10578),
.Y(n_13271)
);

OAI221xp5_ASAP7_75t_L g13272 ( 
.A1(n_11870),
.A2(n_10906),
.B1(n_10893),
.B2(n_10863),
.C(n_9401),
.Y(n_13272)
);

AND2x4_ASAP7_75t_L g13273 ( 
.A(n_11814),
.B(n_11892),
.Y(n_13273)
);

AOI21xp5_ASAP7_75t_L g13274 ( 
.A1(n_11986),
.A2(n_8792),
.B(n_8753),
.Y(n_13274)
);

AOI22xp33_ASAP7_75t_SL g13275 ( 
.A1(n_11843),
.A2(n_11462),
.B1(n_11517),
.B2(n_11514),
.Y(n_13275)
);

AOI22xp33_ASAP7_75t_SL g13276 ( 
.A1(n_11462),
.A2(n_10559),
.B1(n_8456),
.B2(n_9656),
.Y(n_13276)
);

INVx4_ASAP7_75t_L g13277 ( 
.A(n_11970),
.Y(n_13277)
);

OAI22xp5_ASAP7_75t_L g13278 ( 
.A1(n_11609),
.A2(n_10320),
.B1(n_10309),
.B2(n_8232),
.Y(n_13278)
);

AO31x2_ASAP7_75t_L g13279 ( 
.A1(n_11162),
.A2(n_10655),
.A3(n_10661),
.B(n_10652),
.Y(n_13279)
);

HB1xp67_ASAP7_75t_L g13280 ( 
.A(n_11230),
.Y(n_13280)
);

AOI22xp33_ASAP7_75t_SL g13281 ( 
.A1(n_11517),
.A2(n_8456),
.B1(n_9656),
.B2(n_8449),
.Y(n_13281)
);

OAI221xp5_ASAP7_75t_L g13282 ( 
.A1(n_11870),
.A2(n_10906),
.B1(n_10893),
.B2(n_9401),
.C(n_10423),
.Y(n_13282)
);

AOI22xp33_ASAP7_75t_SL g13283 ( 
.A1(n_11629),
.A2(n_9656),
.B1(n_8449),
.B2(n_8675),
.Y(n_13283)
);

AO21x2_ASAP7_75t_L g13284 ( 
.A1(n_11163),
.A2(n_10865),
.B(n_10526),
.Y(n_13284)
);

OAI21xp33_ASAP7_75t_L g13285 ( 
.A1(n_11232),
.A2(n_9936),
.B(n_9904),
.Y(n_13285)
);

AOI22xp33_ASAP7_75t_L g13286 ( 
.A1(n_11156),
.A2(n_9509),
.B1(n_8981),
.B2(n_10320),
.Y(n_13286)
);

INVx1_ASAP7_75t_L g13287 ( 
.A(n_11234),
.Y(n_13287)
);

AOI22xp33_ASAP7_75t_L g13288 ( 
.A1(n_11164),
.A2(n_11180),
.B1(n_11195),
.B2(n_11175),
.Y(n_13288)
);

AOI22xp33_ASAP7_75t_L g13289 ( 
.A1(n_11175),
.A2(n_9509),
.B1(n_8981),
.B2(n_8936),
.Y(n_13289)
);

O2A1O1Ixp33_ASAP7_75t_SL g13290 ( 
.A1(n_11991),
.A2(n_8883),
.B(n_10155),
.C(n_9252),
.Y(n_13290)
);

INVx2_ASAP7_75t_L g13291 ( 
.A(n_11165),
.Y(n_13291)
);

BUFx6f_ASAP7_75t_L g13292 ( 
.A(n_11180),
.Y(n_13292)
);

AOI221xp5_ASAP7_75t_L g13293 ( 
.A1(n_11165),
.A2(n_11015),
.B1(n_11009),
.B2(n_10740),
.C(n_10749),
.Y(n_13293)
);

AOI221xp5_ASAP7_75t_L g13294 ( 
.A1(n_11167),
.A2(n_11015),
.B1(n_11009),
.B2(n_10740),
.C(n_10749),
.Y(n_13294)
);

NOR2xp33_ASAP7_75t_L g13295 ( 
.A(n_11195),
.B(n_11814),
.Y(n_13295)
);

CKINVDCx5p33_ASAP7_75t_R g13296 ( 
.A(n_11892),
.Y(n_13296)
);

AOI222xp33_ASAP7_75t_L g13297 ( 
.A1(n_11167),
.A2(n_9386),
.B1(n_8737),
.B2(n_8589),
.C1(n_8765),
.C2(n_8728),
.Y(n_13297)
);

AOI22xp33_ASAP7_75t_L g13298 ( 
.A1(n_11965),
.A2(n_9509),
.B1(n_8936),
.B2(n_9271),
.Y(n_13298)
);

AND2x2_ASAP7_75t_L g13299 ( 
.A(n_11964),
.B(n_9713),
.Y(n_13299)
);

AOI22xp33_ASAP7_75t_L g13300 ( 
.A1(n_11965),
.A2(n_9509),
.B1(n_9271),
.B2(n_9025),
.Y(n_13300)
);

AOI22xp33_ASAP7_75t_L g13301 ( 
.A1(n_11965),
.A2(n_9509),
.B1(n_9025),
.B2(n_8798),
.Y(n_13301)
);

OAI22xp5_ASAP7_75t_L g13302 ( 
.A1(n_11629),
.A2(n_8232),
.B1(n_8955),
.B2(n_8401),
.Y(n_13302)
);

BUFx3_ASAP7_75t_L g13303 ( 
.A(n_12033),
.Y(n_13303)
);

INVx2_ASAP7_75t_L g13304 ( 
.A(n_11172),
.Y(n_13304)
);

AOI221xp5_ASAP7_75t_L g13305 ( 
.A1(n_11172),
.A2(n_10745),
.B1(n_10771),
.B2(n_10752),
.C(n_10748),
.Y(n_13305)
);

HB1xp67_ASAP7_75t_L g13306 ( 
.A(n_11235),
.Y(n_13306)
);

INVx2_ASAP7_75t_L g13307 ( 
.A(n_11178),
.Y(n_13307)
);

BUFx2_ASAP7_75t_L g13308 ( 
.A(n_12033),
.Y(n_13308)
);

AOI22xp33_ASAP7_75t_SL g13309 ( 
.A1(n_11629),
.A2(n_8449),
.B1(n_8675),
.B2(n_8498),
.Y(n_13309)
);

AOI22xp33_ASAP7_75t_SL g13310 ( 
.A1(n_11681),
.A2(n_8498),
.B1(n_8767),
.B2(n_8675),
.Y(n_13310)
);

OAI211xp5_ASAP7_75t_L g13311 ( 
.A1(n_12032),
.A2(n_10961),
.B(n_11019),
.C(n_10999),
.Y(n_13311)
);

OAI22xp5_ASAP7_75t_SL g13312 ( 
.A1(n_11459),
.A2(n_7564),
.B1(n_7777),
.B2(n_7722),
.Y(n_13312)
);

NAND2xp5_ASAP7_75t_L g13313 ( 
.A(n_11222),
.B(n_8652),
.Y(n_13313)
);

NAND3xp33_ASAP7_75t_L g13314 ( 
.A(n_12166),
.B(n_10999),
.C(n_10961),
.Y(n_13314)
);

AND2x2_ASAP7_75t_L g13315 ( 
.A(n_11966),
.B(n_9724),
.Y(n_13315)
);

OAI22xp33_ASAP7_75t_L g13316 ( 
.A1(n_11205),
.A2(n_8401),
.B1(n_8955),
.B2(n_8232),
.Y(n_13316)
);

OR2x2_ASAP7_75t_L g13317 ( 
.A(n_12367),
.B(n_10048),
.Y(n_13317)
);

AND2x2_ASAP7_75t_L g13318 ( 
.A(n_12463),
.B(n_11580),
.Y(n_13318)
);

OR2x2_ASAP7_75t_L g13319 ( 
.A(n_12447),
.B(n_10057),
.Y(n_13319)
);

AND2x2_ASAP7_75t_L g13320 ( 
.A(n_12587),
.B(n_11997),
.Y(n_13320)
);

OR2x2_ASAP7_75t_L g13321 ( 
.A(n_12449),
.B(n_10057),
.Y(n_13321)
);

INVx2_ASAP7_75t_L g13322 ( 
.A(n_12384),
.Y(n_13322)
);

NAND2xp5_ASAP7_75t_L g13323 ( 
.A(n_12302),
.B(n_8652),
.Y(n_13323)
);

AND2x2_ASAP7_75t_L g13324 ( 
.A(n_12619),
.B(n_12022),
.Y(n_13324)
);

AND2x4_ASAP7_75t_L g13325 ( 
.A(n_12374),
.B(n_11991),
.Y(n_13325)
);

NAND2xp5_ASAP7_75t_L g13326 ( 
.A(n_12289),
.B(n_8652),
.Y(n_13326)
);

BUFx3_ASAP7_75t_L g13327 ( 
.A(n_12426),
.Y(n_13327)
);

BUFx6f_ASAP7_75t_L g13328 ( 
.A(n_12569),
.Y(n_13328)
);

AND2x2_ASAP7_75t_L g13329 ( 
.A(n_12387),
.B(n_11992),
.Y(n_13329)
);

BUFx3_ASAP7_75t_L g13330 ( 
.A(n_12549),
.Y(n_13330)
);

INVx1_ASAP7_75t_L g13331 ( 
.A(n_12466),
.Y(n_13331)
);

INVx1_ASAP7_75t_L g13332 ( 
.A(n_12550),
.Y(n_13332)
);

NAND2xp5_ASAP7_75t_L g13333 ( 
.A(n_12297),
.B(n_12751),
.Y(n_13333)
);

AOI22xp33_ASAP7_75t_L g13334 ( 
.A1(n_12448),
.A2(n_11513),
.B1(n_11425),
.B2(n_11681),
.Y(n_13334)
);

INVx2_ASAP7_75t_L g13335 ( 
.A(n_12523),
.Y(n_13335)
);

INVx1_ASAP7_75t_L g13336 ( 
.A(n_12612),
.Y(n_13336)
);

NAND2xp5_ASAP7_75t_L g13337 ( 
.A(n_12278),
.B(n_8652),
.Y(n_13337)
);

NOR2x1_ASAP7_75t_SL g13338 ( 
.A(n_12777),
.B(n_12927),
.Y(n_13338)
);

BUFx3_ASAP7_75t_L g13339 ( 
.A(n_12366),
.Y(n_13339)
);

AOI22xp33_ASAP7_75t_L g13340 ( 
.A1(n_12455),
.A2(n_11513),
.B1(n_11425),
.B2(n_11681),
.Y(n_13340)
);

INVx1_ASAP7_75t_L g13341 ( 
.A(n_12632),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_12272),
.B(n_11992),
.Y(n_13342)
);

NAND2xp5_ASAP7_75t_L g13343 ( 
.A(n_12286),
.B(n_11587),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_12272),
.B(n_12334),
.Y(n_13344)
);

INVx3_ASAP7_75t_L g13345 ( 
.A(n_12623),
.Y(n_13345)
);

BUFx2_ASAP7_75t_L g13346 ( 
.A(n_13051),
.Y(n_13346)
);

NAND2xp5_ASAP7_75t_L g13347 ( 
.A(n_12311),
.B(n_11587),
.Y(n_13347)
);

NOR2x1_ASAP7_75t_L g13348 ( 
.A(n_12304),
.B(n_11630),
.Y(n_13348)
);

INVx2_ASAP7_75t_L g13349 ( 
.A(n_12908),
.Y(n_13349)
);

INVxp67_ASAP7_75t_L g13350 ( 
.A(n_12841),
.Y(n_13350)
);

AND2x2_ASAP7_75t_L g13351 ( 
.A(n_12697),
.B(n_11630),
.Y(n_13351)
);

AOI22xp33_ASAP7_75t_L g13352 ( 
.A1(n_12320),
.A2(n_11513),
.B1(n_11425),
.B2(n_11684),
.Y(n_13352)
);

HB1xp67_ASAP7_75t_L g13353 ( 
.A(n_12282),
.Y(n_13353)
);

NAND2xp5_ASAP7_75t_L g13354 ( 
.A(n_12318),
.B(n_11587),
.Y(n_13354)
);

AND2x2_ASAP7_75t_L g13355 ( 
.A(n_12739),
.B(n_11653),
.Y(n_13355)
);

NAND2xp5_ASAP7_75t_L g13356 ( 
.A(n_12359),
.B(n_11587),
.Y(n_13356)
);

AND2x4_ASAP7_75t_SL g13357 ( 
.A(n_12686),
.B(n_12271),
.Y(n_13357)
);

HB1xp67_ASAP7_75t_L g13358 ( 
.A(n_12298),
.Y(n_13358)
);

INVx2_ASAP7_75t_L g13359 ( 
.A(n_12969),
.Y(n_13359)
);

NAND2xp5_ASAP7_75t_L g13360 ( 
.A(n_12469),
.B(n_11425),
.Y(n_13360)
);

AND2x4_ASAP7_75t_L g13361 ( 
.A(n_13151),
.B(n_11464),
.Y(n_13361)
);

NAND2xp5_ASAP7_75t_L g13362 ( 
.A(n_12322),
.B(n_11513),
.Y(n_13362)
);

BUFx6f_ASAP7_75t_L g13363 ( 
.A(n_12496),
.Y(n_13363)
);

NAND2xp5_ASAP7_75t_L g13364 ( 
.A(n_12285),
.B(n_11653),
.Y(n_13364)
);

AND2x2_ASAP7_75t_L g13365 ( 
.A(n_12262),
.B(n_11747),
.Y(n_13365)
);

AND2x4_ASAP7_75t_L g13366 ( 
.A(n_12293),
.B(n_11464),
.Y(n_13366)
);

BUFx12f_ASAP7_75t_L g13367 ( 
.A(n_12271),
.Y(n_13367)
);

AOI22xp33_ASAP7_75t_L g13368 ( 
.A1(n_12829),
.A2(n_11797),
.B1(n_11823),
.B2(n_11684),
.Y(n_13368)
);

OR2x2_ASAP7_75t_L g13369 ( 
.A(n_12490),
.B(n_10063),
.Y(n_13369)
);

AND2x2_ASAP7_75t_L g13370 ( 
.A(n_12266),
.B(n_11747),
.Y(n_13370)
);

INVx2_ASAP7_75t_L g13371 ( 
.A(n_12866),
.Y(n_13371)
);

INVx2_ASAP7_75t_L g13372 ( 
.A(n_12350),
.Y(n_13372)
);

AND2x2_ASAP7_75t_L g13373 ( 
.A(n_12729),
.B(n_11758),
.Y(n_13373)
);

INVxp67_ASAP7_75t_L g13374 ( 
.A(n_12425),
.Y(n_13374)
);

AND2x2_ASAP7_75t_L g13375 ( 
.A(n_12312),
.B(n_11758),
.Y(n_13375)
);

NAND2xp5_ASAP7_75t_L g13376 ( 
.A(n_12890),
.B(n_9058),
.Y(n_13376)
);

INVx2_ASAP7_75t_SL g13377 ( 
.A(n_12442),
.Y(n_13377)
);

INVx2_ASAP7_75t_L g13378 ( 
.A(n_13158),
.Y(n_13378)
);

HB1xp67_ASAP7_75t_L g13379 ( 
.A(n_12678),
.Y(n_13379)
);

INVx1_ASAP7_75t_L g13380 ( 
.A(n_12634),
.Y(n_13380)
);

INVx2_ASAP7_75t_SL g13381 ( 
.A(n_12292),
.Y(n_13381)
);

BUFx3_ASAP7_75t_L g13382 ( 
.A(n_12269),
.Y(n_13382)
);

NAND2xp5_ASAP7_75t_L g13383 ( 
.A(n_12287),
.B(n_9058),
.Y(n_13383)
);

INVx2_ASAP7_75t_L g13384 ( 
.A(n_12771),
.Y(n_13384)
);

INVx1_ASAP7_75t_L g13385 ( 
.A(n_12669),
.Y(n_13385)
);

HB1xp67_ASAP7_75t_L g13386 ( 
.A(n_12767),
.Y(n_13386)
);

AND2x2_ASAP7_75t_L g13387 ( 
.A(n_12315),
.B(n_11728),
.Y(n_13387)
);

INVx1_ASAP7_75t_L g13388 ( 
.A(n_12699),
.Y(n_13388)
);

INVx1_ASAP7_75t_L g13389 ( 
.A(n_12752),
.Y(n_13389)
);

AND2x2_ASAP7_75t_L g13390 ( 
.A(n_12452),
.B(n_11728),
.Y(n_13390)
);

INVx2_ASAP7_75t_L g13391 ( 
.A(n_12299),
.Y(n_13391)
);

AND2x2_ASAP7_75t_L g13392 ( 
.A(n_13045),
.B(n_11735),
.Y(n_13392)
);

NOR2xp33_ASAP7_75t_L g13393 ( 
.A(n_12433),
.B(n_11735),
.Y(n_13393)
);

BUFx2_ASAP7_75t_L g13394 ( 
.A(n_12835),
.Y(n_13394)
);

AND2x4_ASAP7_75t_L g13395 ( 
.A(n_13057),
.B(n_13081),
.Y(n_13395)
);

INVx2_ASAP7_75t_L g13396 ( 
.A(n_13257),
.Y(n_13396)
);

INVx2_ASAP7_75t_L g13397 ( 
.A(n_13257),
.Y(n_13397)
);

BUFx2_ASAP7_75t_L g13398 ( 
.A(n_12754),
.Y(n_13398)
);

INVx1_ASAP7_75t_SL g13399 ( 
.A(n_12476),
.Y(n_13399)
);

AND2x2_ASAP7_75t_L g13400 ( 
.A(n_12368),
.B(n_11490),
.Y(n_13400)
);

INVx1_ASAP7_75t_L g13401 ( 
.A(n_13193),
.Y(n_13401)
);

OR2x2_ASAP7_75t_L g13402 ( 
.A(n_12291),
.B(n_10063),
.Y(n_13402)
);

INVx2_ASAP7_75t_L g13403 ( 
.A(n_13257),
.Y(n_13403)
);

INVx2_ASAP7_75t_L g13404 ( 
.A(n_13292),
.Y(n_13404)
);

INVx1_ASAP7_75t_L g13405 ( 
.A(n_13227),
.Y(n_13405)
);

INVx1_ASAP7_75t_L g13406 ( 
.A(n_13280),
.Y(n_13406)
);

INVx1_ASAP7_75t_L g13407 ( 
.A(n_13306),
.Y(n_13407)
);

INVx2_ASAP7_75t_L g13408 ( 
.A(n_13292),
.Y(n_13408)
);

BUFx6f_ASAP7_75t_L g13409 ( 
.A(n_12382),
.Y(n_13409)
);

BUFx3_ASAP7_75t_L g13410 ( 
.A(n_12744),
.Y(n_13410)
);

BUFx2_ASAP7_75t_L g13411 ( 
.A(n_12754),
.Y(n_13411)
);

NOR2xp33_ASAP7_75t_L g13412 ( 
.A(n_12510),
.B(n_11490),
.Y(n_13412)
);

INVx2_ASAP7_75t_L g13413 ( 
.A(n_13292),
.Y(n_13413)
);

INVx1_ASAP7_75t_L g13414 ( 
.A(n_12276),
.Y(n_13414)
);

AND2x2_ASAP7_75t_L g13415 ( 
.A(n_13248),
.B(n_13273),
.Y(n_13415)
);

HB1xp67_ASAP7_75t_L g13416 ( 
.A(n_13174),
.Y(n_13416)
);

CKINVDCx5p33_ASAP7_75t_R g13417 ( 
.A(n_12450),
.Y(n_13417)
);

INVx1_ASAP7_75t_L g13418 ( 
.A(n_12279),
.Y(n_13418)
);

AND2x2_ASAP7_75t_L g13419 ( 
.A(n_13273),
.B(n_11459),
.Y(n_13419)
);

INVx3_ASAP7_75t_L g13420 ( 
.A(n_12292),
.Y(n_13420)
);

INVx2_ASAP7_75t_L g13421 ( 
.A(n_13152),
.Y(n_13421)
);

HB1xp67_ASAP7_75t_L g13422 ( 
.A(n_12339),
.Y(n_13422)
);

NAND2xp5_ASAP7_75t_L g13423 ( 
.A(n_12303),
.B(n_9058),
.Y(n_13423)
);

AOI22xp33_ASAP7_75t_SL g13424 ( 
.A1(n_12385),
.A2(n_11684),
.B1(n_11823),
.B2(n_11797),
.Y(n_13424)
);

AND2x2_ASAP7_75t_L g13425 ( 
.A(n_13179),
.B(n_11484),
.Y(n_13425)
);

INVx2_ASAP7_75t_L g13426 ( 
.A(n_13152),
.Y(n_13426)
);

INVx1_ASAP7_75t_L g13427 ( 
.A(n_12300),
.Y(n_13427)
);

AOI22xp33_ASAP7_75t_L g13428 ( 
.A1(n_12280),
.A2(n_11823),
.B1(n_11836),
.B2(n_11797),
.Y(n_13428)
);

INVx2_ASAP7_75t_L g13429 ( 
.A(n_13164),
.Y(n_13429)
);

INVx1_ASAP7_75t_L g13430 ( 
.A(n_12348),
.Y(n_13430)
);

AND2x2_ASAP7_75t_L g13431 ( 
.A(n_13181),
.B(n_11484),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_13187),
.B(n_13220),
.Y(n_13432)
);

AND2x4_ASAP7_75t_SL g13433 ( 
.A(n_12779),
.B(n_8063),
.Y(n_13433)
);

AND2x4_ASAP7_75t_L g13434 ( 
.A(n_13057),
.B(n_11484),
.Y(n_13434)
);

AO31x2_ASAP7_75t_L g13435 ( 
.A1(n_12281),
.A2(n_11192),
.A3(n_11197),
.B(n_11178),
.Y(n_13435)
);

OR2x2_ASAP7_75t_L g13436 ( 
.A(n_12352),
.B(n_10066),
.Y(n_13436)
);

INVx1_ASAP7_75t_L g13437 ( 
.A(n_12360),
.Y(n_13437)
);

BUFx2_ASAP7_75t_L g13438 ( 
.A(n_12753),
.Y(n_13438)
);

AND2x2_ASAP7_75t_L g13439 ( 
.A(n_13228),
.B(n_11619),
.Y(n_13439)
);

AND2x2_ASAP7_75t_L g13440 ( 
.A(n_12708),
.B(n_11619),
.Y(n_13440)
);

OR2x2_ASAP7_75t_L g13441 ( 
.A(n_12390),
.B(n_12419),
.Y(n_13441)
);

INVx2_ASAP7_75t_L g13442 ( 
.A(n_13164),
.Y(n_13442)
);

AND2x2_ASAP7_75t_L g13443 ( 
.A(n_12710),
.B(n_12377),
.Y(n_13443)
);

AND2x4_ASAP7_75t_L g13444 ( 
.A(n_13081),
.B(n_11619),
.Y(n_13444)
);

AOI21xp33_ASAP7_75t_L g13445 ( 
.A1(n_12370),
.A2(n_11197),
.B(n_11192),
.Y(n_13445)
);

AND2x4_ASAP7_75t_L g13446 ( 
.A(n_13087),
.B(n_11511),
.Y(n_13446)
);

AND2x2_ASAP7_75t_L g13447 ( 
.A(n_12379),
.B(n_11807),
.Y(n_13447)
);

OR2x2_ASAP7_75t_L g13448 ( 
.A(n_12342),
.B(n_10066),
.Y(n_13448)
);

INVx3_ASAP7_75t_L g13449 ( 
.A(n_12364),
.Y(n_13449)
);

INVx1_ASAP7_75t_L g13450 ( 
.A(n_12362),
.Y(n_13450)
);

INVxp67_ASAP7_75t_L g13451 ( 
.A(n_12721),
.Y(n_13451)
);

INVx2_ASAP7_75t_SL g13452 ( 
.A(n_12364),
.Y(n_13452)
);

INVx2_ASAP7_75t_L g13453 ( 
.A(n_13165),
.Y(n_13453)
);

AND2x2_ASAP7_75t_L g13454 ( 
.A(n_12400),
.B(n_11807),
.Y(n_13454)
);

BUFx2_ASAP7_75t_L g13455 ( 
.A(n_12786),
.Y(n_13455)
);

INVx2_ASAP7_75t_L g13456 ( 
.A(n_13165),
.Y(n_13456)
);

NAND2xp5_ASAP7_75t_L g13457 ( 
.A(n_12323),
.B(n_9058),
.Y(n_13457)
);

INVx2_ASAP7_75t_L g13458 ( 
.A(n_13185),
.Y(n_13458)
);

AND2x2_ASAP7_75t_L g13459 ( 
.A(n_12422),
.B(n_11807),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_12369),
.Y(n_13460)
);

OAI222xp33_ASAP7_75t_L g13461 ( 
.A1(n_12372),
.A2(n_12461),
.B1(n_12439),
.B2(n_12361),
.C1(n_12325),
.C2(n_12456),
.Y(n_13461)
);

BUFx6f_ASAP7_75t_L g13462 ( 
.A(n_12467),
.Y(n_13462)
);

INVx1_ASAP7_75t_L g13463 ( 
.A(n_12378),
.Y(n_13463)
);

BUFx2_ASAP7_75t_L g13464 ( 
.A(n_12792),
.Y(n_13464)
);

BUFx6f_ASAP7_75t_L g13465 ( 
.A(n_12531),
.Y(n_13465)
);

AND2x2_ASAP7_75t_L g13466 ( 
.A(n_12316),
.B(n_12982),
.Y(n_13466)
);

NAND2xp5_ASAP7_75t_L g13467 ( 
.A(n_12301),
.B(n_9058),
.Y(n_13467)
);

INVx2_ASAP7_75t_L g13468 ( 
.A(n_13185),
.Y(n_13468)
);

INVx2_ASAP7_75t_L g13469 ( 
.A(n_13222),
.Y(n_13469)
);

AND2x4_ASAP7_75t_L g13470 ( 
.A(n_13087),
.B(n_11511),
.Y(n_13470)
);

OR2x6_ASAP7_75t_L g13471 ( 
.A(n_12375),
.B(n_12327),
.Y(n_13471)
);

INVx2_ASAP7_75t_L g13472 ( 
.A(n_13222),
.Y(n_13472)
);

AND2x2_ASAP7_75t_L g13473 ( 
.A(n_13035),
.B(n_11899),
.Y(n_13473)
);

AND2x2_ASAP7_75t_L g13474 ( 
.A(n_13238),
.B(n_11899),
.Y(n_13474)
);

AND2x2_ASAP7_75t_L g13475 ( 
.A(n_13308),
.B(n_11899),
.Y(n_13475)
);

INVx1_ASAP7_75t_L g13476 ( 
.A(n_12381),
.Y(n_13476)
);

INVx2_ASAP7_75t_L g13477 ( 
.A(n_12561),
.Y(n_13477)
);

OR2x2_ASAP7_75t_L g13478 ( 
.A(n_12546),
.B(n_10070),
.Y(n_13478)
);

BUFx12f_ASAP7_75t_L g13479 ( 
.A(n_12629),
.Y(n_13479)
);

INVx1_ASAP7_75t_L g13480 ( 
.A(n_12412),
.Y(n_13480)
);

OR2x2_ASAP7_75t_L g13481 ( 
.A(n_12273),
.B(n_10070),
.Y(n_13481)
);

AO31x2_ASAP7_75t_L g13482 ( 
.A1(n_12346),
.A2(n_11206),
.A3(n_11208),
.B(n_11205),
.Y(n_13482)
);

INVx2_ASAP7_75t_SL g13483 ( 
.A(n_12375),
.Y(n_13483)
);

AND2x2_ASAP7_75t_L g13484 ( 
.A(n_12763),
.B(n_12154),
.Y(n_13484)
);

INVxp67_ASAP7_75t_L g13485 ( 
.A(n_12420),
.Y(n_13485)
);

INVx1_ASAP7_75t_L g13486 ( 
.A(n_12418),
.Y(n_13486)
);

INVx2_ASAP7_75t_L g13487 ( 
.A(n_13303),
.Y(n_13487)
);

OR2x6_ASAP7_75t_L g13488 ( 
.A(n_12327),
.B(n_7722),
.Y(n_13488)
);

INVx1_ASAP7_75t_L g13489 ( 
.A(n_12431),
.Y(n_13489)
);

INVx1_ASAP7_75t_L g13490 ( 
.A(n_12432),
.Y(n_13490)
);

INVx2_ASAP7_75t_L g13491 ( 
.A(n_12828),
.Y(n_13491)
);

NAND2xp5_ASAP7_75t_L g13492 ( 
.A(n_12309),
.B(n_9058),
.Y(n_13492)
);

INVx1_ASAP7_75t_L g13493 ( 
.A(n_12443),
.Y(n_13493)
);

HB1xp67_ASAP7_75t_L g13494 ( 
.A(n_12495),
.Y(n_13494)
);

OR2x2_ASAP7_75t_L g13495 ( 
.A(n_12516),
.B(n_10076),
.Y(n_13495)
);

NAND2xp5_ASAP7_75t_L g13496 ( 
.A(n_12308),
.B(n_9058),
.Y(n_13496)
);

INVx1_ASAP7_75t_L g13497 ( 
.A(n_12451),
.Y(n_13497)
);

INVx2_ASAP7_75t_L g13498 ( 
.A(n_12828),
.Y(n_13498)
);

BUFx3_ASAP7_75t_L g13499 ( 
.A(n_12643),
.Y(n_13499)
);

HB1xp67_ASAP7_75t_L g13500 ( 
.A(n_12579),
.Y(n_13500)
);

AND2x2_ASAP7_75t_L g13501 ( 
.A(n_12343),
.B(n_12154),
.Y(n_13501)
);

NAND2x1_ASAP7_75t_L g13502 ( 
.A(n_12888),
.B(n_11832),
.Y(n_13502)
);

INVx1_ASAP7_75t_L g13503 ( 
.A(n_12473),
.Y(n_13503)
);

INVx2_ASAP7_75t_L g13504 ( 
.A(n_12828),
.Y(n_13504)
);

AND2x4_ASAP7_75t_L g13505 ( 
.A(n_13028),
.B(n_11511),
.Y(n_13505)
);

AND2x2_ASAP7_75t_L g13506 ( 
.A(n_12435),
.B(n_12154),
.Y(n_13506)
);

INVx2_ASAP7_75t_SL g13507 ( 
.A(n_12652),
.Y(n_13507)
);

AND2x2_ASAP7_75t_L g13508 ( 
.A(n_12453),
.B(n_12182),
.Y(n_13508)
);

HB1xp67_ASAP7_75t_L g13509 ( 
.A(n_12606),
.Y(n_13509)
);

INVx2_ASAP7_75t_L g13510 ( 
.A(n_12828),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_12486),
.Y(n_13511)
);

NOR2xp33_ASAP7_75t_L g13512 ( 
.A(n_12647),
.B(n_10773),
.Y(n_13512)
);

AND2x2_ASAP7_75t_L g13513 ( 
.A(n_12454),
.B(n_12182),
.Y(n_13513)
);

NAND2xp5_ASAP7_75t_L g13514 ( 
.A(n_12404),
.B(n_9058),
.Y(n_13514)
);

INVx1_ASAP7_75t_L g13515 ( 
.A(n_12487),
.Y(n_13515)
);

INVx1_ASAP7_75t_L g13516 ( 
.A(n_12502),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_12508),
.Y(n_13517)
);

INVx2_ASAP7_75t_L g13518 ( 
.A(n_12828),
.Y(n_13518)
);

AND2x2_ASAP7_75t_L g13519 ( 
.A(n_12978),
.B(n_12182),
.Y(n_13519)
);

OR2x6_ASAP7_75t_SL g13520 ( 
.A(n_13296),
.B(n_10038),
.Y(n_13520)
);

INVx2_ASAP7_75t_L g13521 ( 
.A(n_12947),
.Y(n_13521)
);

INVx2_ASAP7_75t_L g13522 ( 
.A(n_12947),
.Y(n_13522)
);

AND2x2_ASAP7_75t_L g13523 ( 
.A(n_12616),
.B(n_11511),
.Y(n_13523)
);

CKINVDCx16_ASAP7_75t_R g13524 ( 
.A(n_12633),
.Y(n_13524)
);

INVx1_ASAP7_75t_L g13525 ( 
.A(n_12526),
.Y(n_13525)
);

INVx2_ASAP7_75t_L g13526 ( 
.A(n_12947),
.Y(n_13526)
);

INVx1_ASAP7_75t_L g13527 ( 
.A(n_12537),
.Y(n_13527)
);

INVx1_ASAP7_75t_L g13528 ( 
.A(n_12539),
.Y(n_13528)
);

OR2x2_ASAP7_75t_L g13529 ( 
.A(n_12704),
.B(n_10076),
.Y(n_13529)
);

NAND2xp5_ASAP7_75t_L g13530 ( 
.A(n_12264),
.B(n_9072),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_12540),
.Y(n_13531)
);

INVx2_ASAP7_75t_SL g13532 ( 
.A(n_12720),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_13135),
.B(n_10961),
.Y(n_13533)
);

AND2x2_ASAP7_75t_L g13534 ( 
.A(n_13139),
.B(n_10999),
.Y(n_13534)
);

AND2x2_ASAP7_75t_L g13535 ( 
.A(n_12480),
.B(n_11019),
.Y(n_13535)
);

INVx1_ASAP7_75t_L g13536 ( 
.A(n_12552),
.Y(n_13536)
);

AND2x4_ASAP7_75t_SL g13537 ( 
.A(n_13182),
.B(n_12417),
.Y(n_13537)
);

AND2x2_ASAP7_75t_L g13538 ( 
.A(n_12530),
.B(n_11019),
.Y(n_13538)
);

NAND2xp5_ASAP7_75t_L g13539 ( 
.A(n_12475),
.B(n_9072),
.Y(n_13539)
);

NAND2xp5_ASAP7_75t_L g13540 ( 
.A(n_12527),
.B(n_9072),
.Y(n_13540)
);

AND2x2_ASAP7_75t_L g13541 ( 
.A(n_12535),
.B(n_11426),
.Y(n_13541)
);

AND2x2_ASAP7_75t_L g13542 ( 
.A(n_12554),
.B(n_11449),
.Y(n_13542)
);

INVx2_ASAP7_75t_L g13543 ( 
.A(n_12947),
.Y(n_13543)
);

AND2x2_ASAP7_75t_L g13544 ( 
.A(n_13315),
.B(n_11473),
.Y(n_13544)
);

INVx2_ASAP7_75t_L g13545 ( 
.A(n_12947),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_12557),
.Y(n_13546)
);

INVx1_ASAP7_75t_L g13547 ( 
.A(n_12565),
.Y(n_13547)
);

INVx2_ASAP7_75t_L g13548 ( 
.A(n_12483),
.Y(n_13548)
);

AND2x4_ASAP7_75t_L g13549 ( 
.A(n_12777),
.B(n_11520),
.Y(n_13549)
);

INVx1_ASAP7_75t_L g13550 ( 
.A(n_12575),
.Y(n_13550)
);

NAND2xp5_ASAP7_75t_L g13551 ( 
.A(n_12416),
.B(n_9072),
.Y(n_13551)
);

NAND2xp5_ASAP7_75t_L g13552 ( 
.A(n_12590),
.B(n_9072),
.Y(n_13552)
);

INVx1_ASAP7_75t_L g13553 ( 
.A(n_12576),
.Y(n_13553)
);

HB1xp67_ASAP7_75t_L g13554 ( 
.A(n_12689),
.Y(n_13554)
);

AND2x2_ASAP7_75t_L g13555 ( 
.A(n_13299),
.B(n_12667),
.Y(n_13555)
);

HB1xp67_ASAP7_75t_L g13556 ( 
.A(n_12600),
.Y(n_13556)
);

AND2x4_ASAP7_75t_L g13557 ( 
.A(n_12927),
.B(n_11592),
.Y(n_13557)
);

INVx2_ASAP7_75t_L g13558 ( 
.A(n_12483),
.Y(n_13558)
);

AND2x2_ASAP7_75t_L g13559 ( 
.A(n_12892),
.B(n_11592),
.Y(n_13559)
);

AND2x4_ASAP7_75t_L g13560 ( 
.A(n_13022),
.B(n_12188),
.Y(n_13560)
);

INVxp67_ASAP7_75t_L g13561 ( 
.A(n_12662),
.Y(n_13561)
);

AND2x2_ASAP7_75t_L g13562 ( 
.A(n_12912),
.B(n_12188),
.Y(n_13562)
);

INVx3_ASAP7_75t_L g13563 ( 
.A(n_12663),
.Y(n_13563)
);

INVx2_ASAP7_75t_L g13564 ( 
.A(n_12663),
.Y(n_13564)
);

INVx1_ASAP7_75t_L g13565 ( 
.A(n_12577),
.Y(n_13565)
);

AND2x2_ASAP7_75t_SL g13566 ( 
.A(n_12597),
.B(n_9277),
.Y(n_13566)
);

INVx2_ASAP7_75t_L g13567 ( 
.A(n_12808),
.Y(n_13567)
);

INVx4_ASAP7_75t_L g13568 ( 
.A(n_12345),
.Y(n_13568)
);

INVx3_ASAP7_75t_L g13569 ( 
.A(n_12808),
.Y(n_13569)
);

INVx1_ASAP7_75t_L g13570 ( 
.A(n_12675),
.Y(n_13570)
);

BUFx3_ASAP7_75t_L g13571 ( 
.A(n_12354),
.Y(n_13571)
);

INVx1_ASAP7_75t_L g13572 ( 
.A(n_12692),
.Y(n_13572)
);

BUFx2_ASAP7_75t_SL g13573 ( 
.A(n_12397),
.Y(n_13573)
);

INVx1_ASAP7_75t_L g13574 ( 
.A(n_12702),
.Y(n_13574)
);

AND2x4_ASAP7_75t_L g13575 ( 
.A(n_13022),
.B(n_12188),
.Y(n_13575)
);

NOR2xp33_ASAP7_75t_L g13576 ( 
.A(n_12728),
.B(n_10056),
.Y(n_13576)
);

AND2x2_ASAP7_75t_L g13577 ( 
.A(n_12778),
.B(n_12188),
.Y(n_13577)
);

OR2x2_ASAP7_75t_L g13578 ( 
.A(n_12344),
.B(n_10078),
.Y(n_13578)
);

INVx3_ASAP7_75t_L g13579 ( 
.A(n_12922),
.Y(n_13579)
);

NAND2xp5_ASAP7_75t_L g13580 ( 
.A(n_12603),
.B(n_9072),
.Y(n_13580)
);

INVx2_ASAP7_75t_L g13581 ( 
.A(n_12922),
.Y(n_13581)
);

AND2x2_ASAP7_75t_L g13582 ( 
.A(n_12974),
.B(n_12199),
.Y(n_13582)
);

AND2x2_ASAP7_75t_L g13583 ( 
.A(n_12457),
.B(n_12199),
.Y(n_13583)
);

INVx1_ASAP7_75t_L g13584 ( 
.A(n_12711),
.Y(n_13584)
);

INVx1_ASAP7_75t_L g13585 ( 
.A(n_12716),
.Y(n_13585)
);

AND2x2_ASAP7_75t_L g13586 ( 
.A(n_12468),
.B(n_12199),
.Y(n_13586)
);

INVx1_ASAP7_75t_L g13587 ( 
.A(n_12740),
.Y(n_13587)
);

INVx1_ASAP7_75t_L g13588 ( 
.A(n_12750),
.Y(n_13588)
);

INVx2_ASAP7_75t_L g13589 ( 
.A(n_12968),
.Y(n_13589)
);

AND2x2_ASAP7_75t_L g13590 ( 
.A(n_12584),
.B(n_12588),
.Y(n_13590)
);

INVx5_ASAP7_75t_L g13591 ( 
.A(n_12417),
.Y(n_13591)
);

INVx5_ASAP7_75t_L g13592 ( 
.A(n_12529),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_12758),
.Y(n_13593)
);

AND2x2_ASAP7_75t_L g13594 ( 
.A(n_12782),
.B(n_12199),
.Y(n_13594)
);

AND2x2_ASAP7_75t_L g13595 ( 
.A(n_12783),
.B(n_12209),
.Y(n_13595)
);

INVx1_ASAP7_75t_L g13596 ( 
.A(n_12768),
.Y(n_13596)
);

OR2x2_ASAP7_75t_L g13597 ( 
.A(n_12793),
.B(n_10078),
.Y(n_13597)
);

NAND2xp5_ASAP7_75t_L g13598 ( 
.A(n_12631),
.B(n_9072),
.Y(n_13598)
);

AND2x2_ASAP7_75t_L g13599 ( 
.A(n_13094),
.B(n_12209),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_12772),
.Y(n_13600)
);

NAND2xp5_ASAP7_75t_L g13601 ( 
.A(n_12636),
.B(n_9072),
.Y(n_13601)
);

AOI22xp33_ASAP7_75t_L g13602 ( 
.A1(n_12410),
.A2(n_11898),
.B1(n_11836),
.B2(n_12209),
.Y(n_13602)
);

OR2x2_ASAP7_75t_L g13603 ( 
.A(n_12586),
.B(n_10084),
.Y(n_13603)
);

BUFx6f_ASAP7_75t_L g13604 ( 
.A(n_12529),
.Y(n_13604)
);

AND2x2_ASAP7_75t_L g13605 ( 
.A(n_13094),
.B(n_12209),
.Y(n_13605)
);

BUFx6f_ASAP7_75t_L g13606 ( 
.A(n_12499),
.Y(n_13606)
);

INVx2_ASAP7_75t_L g13607 ( 
.A(n_12968),
.Y(n_13607)
);

AND2x2_ASAP7_75t_L g13608 ( 
.A(n_12592),
.B(n_11972),
.Y(n_13608)
);

INVx1_ASAP7_75t_L g13609 ( 
.A(n_12799),
.Y(n_13609)
);

AND2x4_ASAP7_75t_L g13610 ( 
.A(n_12275),
.B(n_11836),
.Y(n_13610)
);

BUFx3_ASAP7_75t_L g13611 ( 
.A(n_12656),
.Y(n_13611)
);

INVx1_ASAP7_75t_L g13612 ( 
.A(n_12807),
.Y(n_13612)
);

INVx1_ASAP7_75t_L g13613 ( 
.A(n_12826),
.Y(n_13613)
);

NAND2x1_ASAP7_75t_L g13614 ( 
.A(n_12324),
.B(n_11832),
.Y(n_13614)
);

INVx2_ASAP7_75t_L g13615 ( 
.A(n_12999),
.Y(n_13615)
);

INVx2_ASAP7_75t_L g13616 ( 
.A(n_12999),
.Y(n_13616)
);

NAND2xp5_ASAP7_75t_L g13617 ( 
.A(n_12640),
.B(n_10652),
.Y(n_13617)
);

NAND2xp5_ASAP7_75t_L g13618 ( 
.A(n_12666),
.B(n_10655),
.Y(n_13618)
);

AND2x2_ASAP7_75t_L g13619 ( 
.A(n_12607),
.B(n_12001),
.Y(n_13619)
);

AND2x2_ASAP7_75t_L g13620 ( 
.A(n_12609),
.B(n_12016),
.Y(n_13620)
);

INVx1_ASAP7_75t_L g13621 ( 
.A(n_12879),
.Y(n_13621)
);

INVxp67_ASAP7_75t_SL g13622 ( 
.A(n_12321),
.Y(n_13622)
);

BUFx3_ASAP7_75t_L g13623 ( 
.A(n_12656),
.Y(n_13623)
);

OR2x2_ASAP7_75t_L g13624 ( 
.A(n_12658),
.B(n_10084),
.Y(n_13624)
);

INVx2_ASAP7_75t_L g13625 ( 
.A(n_13010),
.Y(n_13625)
);

AND2x2_ASAP7_75t_L g13626 ( 
.A(n_12626),
.B(n_12025),
.Y(n_13626)
);

NAND2xp5_ASAP7_75t_L g13627 ( 
.A(n_12670),
.B(n_10655),
.Y(n_13627)
);

INVx5_ASAP7_75t_L g13628 ( 
.A(n_12889),
.Y(n_13628)
);

INVx1_ASAP7_75t_L g13629 ( 
.A(n_12885),
.Y(n_13629)
);

NAND2xp5_ASAP7_75t_L g13630 ( 
.A(n_12326),
.B(n_10661),
.Y(n_13630)
);

AND2x4_ASAP7_75t_L g13631 ( 
.A(n_12275),
.B(n_11898),
.Y(n_13631)
);

INVx2_ASAP7_75t_L g13632 ( 
.A(n_13010),
.Y(n_13632)
);

AND2x2_ASAP7_75t_L g13633 ( 
.A(n_12641),
.B(n_12037),
.Y(n_13633)
);

AND2x2_ASAP7_75t_L g13634 ( 
.A(n_12655),
.B(n_12049),
.Y(n_13634)
);

NAND2xp5_ASAP7_75t_L g13635 ( 
.A(n_12363),
.B(n_10661),
.Y(n_13635)
);

AND2x2_ASAP7_75t_L g13636 ( 
.A(n_13000),
.B(n_12053),
.Y(n_13636)
);

BUFx2_ASAP7_75t_L g13637 ( 
.A(n_12953),
.Y(n_13637)
);

HB1xp67_ASAP7_75t_SL g13638 ( 
.A(n_12819),
.Y(n_13638)
);

INVx1_ASAP7_75t_L g13639 ( 
.A(n_12896),
.Y(n_13639)
);

INVx1_ASAP7_75t_L g13640 ( 
.A(n_12906),
.Y(n_13640)
);

INVx1_ASAP7_75t_L g13641 ( 
.A(n_12914),
.Y(n_13641)
);

AND2x2_ASAP7_75t_L g13642 ( 
.A(n_12930),
.B(n_12056),
.Y(n_13642)
);

INVx2_ASAP7_75t_L g13643 ( 
.A(n_13040),
.Y(n_13643)
);

OR2x2_ASAP7_75t_L g13644 ( 
.A(n_12694),
.B(n_10087),
.Y(n_13644)
);

AND2x2_ASAP7_75t_L g13645 ( 
.A(n_12935),
.B(n_12060),
.Y(n_13645)
);

INVx2_ASAP7_75t_L g13646 ( 
.A(n_13040),
.Y(n_13646)
);

OAI22xp5_ASAP7_75t_L g13647 ( 
.A1(n_12333),
.A2(n_8239),
.B1(n_8326),
.B2(n_8204),
.Y(n_13647)
);

BUFx6f_ASAP7_75t_L g13648 ( 
.A(n_12499),
.Y(n_13648)
);

AND2x2_ASAP7_75t_L g13649 ( 
.A(n_12961),
.B(n_12074),
.Y(n_13649)
);

HB1xp67_ASAP7_75t_L g13650 ( 
.A(n_13143),
.Y(n_13650)
);

AND2x2_ASAP7_75t_L g13651 ( 
.A(n_13153),
.B(n_12111),
.Y(n_13651)
);

INVx3_ASAP7_75t_L g13652 ( 
.A(n_13096),
.Y(n_13652)
);

INVx3_ASAP7_75t_L g13653 ( 
.A(n_13096),
.Y(n_13653)
);

INVxp67_ASAP7_75t_L g13654 ( 
.A(n_12446),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_13159),
.B(n_12125),
.Y(n_13655)
);

AND2x2_ASAP7_75t_L g13656 ( 
.A(n_13170),
.B(n_12139),
.Y(n_13656)
);

NAND2xp5_ASAP7_75t_L g13657 ( 
.A(n_12337),
.B(n_11239),
.Y(n_13657)
);

INVx1_ASAP7_75t_L g13658 ( 
.A(n_12928),
.Y(n_13658)
);

AND2x2_ASAP7_75t_L g13659 ( 
.A(n_13177),
.B(n_12668),
.Y(n_13659)
);

NAND2xp5_ASAP7_75t_L g13660 ( 
.A(n_12747),
.B(n_11240),
.Y(n_13660)
);

BUFx2_ASAP7_75t_L g13661 ( 
.A(n_12819),
.Y(n_13661)
);

HB1xp67_ASAP7_75t_L g13662 ( 
.A(n_12972),
.Y(n_13662)
);

INVx2_ASAP7_75t_L g13663 ( 
.A(n_12795),
.Y(n_13663)
);

INVx2_ASAP7_75t_L g13664 ( 
.A(n_12834),
.Y(n_13664)
);

HB1xp67_ASAP7_75t_L g13665 ( 
.A(n_12938),
.Y(n_13665)
);

AND2x2_ASAP7_75t_L g13666 ( 
.A(n_12695),
.B(n_12143),
.Y(n_13666)
);

OR2x2_ASAP7_75t_L g13667 ( 
.A(n_12265),
.B(n_10087),
.Y(n_13667)
);

INVx2_ASAP7_75t_L g13668 ( 
.A(n_12836),
.Y(n_13668)
);

OR2x2_ASAP7_75t_L g13669 ( 
.A(n_12659),
.B(n_10088),
.Y(n_13669)
);

AND2x2_ASAP7_75t_L g13670 ( 
.A(n_12701),
.B(n_12145),
.Y(n_13670)
);

HB1xp67_ASAP7_75t_L g13671 ( 
.A(n_12979),
.Y(n_13671)
);

INVx2_ASAP7_75t_L g13672 ( 
.A(n_12849),
.Y(n_13672)
);

AND2x2_ASAP7_75t_L g13673 ( 
.A(n_12814),
.B(n_12173),
.Y(n_13673)
);

INVx1_ASAP7_75t_L g13674 ( 
.A(n_12956),
.Y(n_13674)
);

AND2x4_ASAP7_75t_L g13675 ( 
.A(n_12277),
.B(n_11898),
.Y(n_13675)
);

BUFx6f_ASAP7_75t_L g13676 ( 
.A(n_12499),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_12967),
.Y(n_13677)
);

INVx1_ASAP7_75t_L g13678 ( 
.A(n_13012),
.Y(n_13678)
);

NAND2xp5_ASAP7_75t_L g13679 ( 
.A(n_12405),
.B(n_11242),
.Y(n_13679)
);

AND2x2_ASAP7_75t_L g13680 ( 
.A(n_12814),
.B(n_12840),
.Y(n_13680)
);

INVx2_ASAP7_75t_L g13681 ( 
.A(n_12874),
.Y(n_13681)
);

INVx4_ASAP7_75t_L g13682 ( 
.A(n_13127),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_13016),
.Y(n_13683)
);

AO21x2_ASAP7_75t_L g13684 ( 
.A1(n_12522),
.A2(n_11208),
.B(n_11206),
.Y(n_13684)
);

AND2x2_ASAP7_75t_L g13685 ( 
.A(n_12840),
.B(n_12880),
.Y(n_13685)
);

OR2x2_ASAP7_75t_L g13686 ( 
.A(n_12677),
.B(n_10088),
.Y(n_13686)
);

INVx2_ASAP7_75t_L g13687 ( 
.A(n_12886),
.Y(n_13687)
);

AND2x2_ASAP7_75t_L g13688 ( 
.A(n_12880),
.B(n_12210),
.Y(n_13688)
);

INVx1_ASAP7_75t_L g13689 ( 
.A(n_13024),
.Y(n_13689)
);

INVx2_ASAP7_75t_L g13690 ( 
.A(n_12894),
.Y(n_13690)
);

INVx2_ASAP7_75t_L g13691 ( 
.A(n_12903),
.Y(n_13691)
);

INVx2_ASAP7_75t_L g13692 ( 
.A(n_12909),
.Y(n_13692)
);

BUFx6f_ASAP7_75t_L g13693 ( 
.A(n_12594),
.Y(n_13693)
);

AND2x2_ASAP7_75t_L g13694 ( 
.A(n_12921),
.B(n_12224),
.Y(n_13694)
);

AND2x2_ASAP7_75t_L g13695 ( 
.A(n_12921),
.B(n_13069),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_13043),
.Y(n_13696)
);

INVx2_ASAP7_75t_L g13697 ( 
.A(n_12918),
.Y(n_13697)
);

AND2x2_ASAP7_75t_L g13698 ( 
.A(n_12274),
.B(n_9724),
.Y(n_13698)
);

NAND2xp5_ASAP7_75t_L g13699 ( 
.A(n_13059),
.B(n_11246),
.Y(n_13699)
);

INVx1_ASAP7_75t_L g13700 ( 
.A(n_13061),
.Y(n_13700)
);

AND2x4_ASAP7_75t_L g13701 ( 
.A(n_12277),
.B(n_11832),
.Y(n_13701)
);

INVx2_ASAP7_75t_L g13702 ( 
.A(n_12919),
.Y(n_13702)
);

INVx3_ASAP7_75t_L g13703 ( 
.A(n_13102),
.Y(n_13703)
);

AND2x2_ASAP7_75t_L g13704 ( 
.A(n_12274),
.B(n_9747),
.Y(n_13704)
);

BUFx6f_ASAP7_75t_L g13705 ( 
.A(n_13080),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13062),
.Y(n_13706)
);

AND2x2_ASAP7_75t_L g13707 ( 
.A(n_13128),
.B(n_13218),
.Y(n_13707)
);

INVx2_ASAP7_75t_L g13708 ( 
.A(n_12934),
.Y(n_13708)
);

AND2x2_ASAP7_75t_L g13709 ( 
.A(n_13218),
.B(n_9747),
.Y(n_13709)
);

BUFx2_ASAP7_75t_L g13710 ( 
.A(n_12661),
.Y(n_13710)
);

INVx1_ASAP7_75t_L g13711 ( 
.A(n_13074),
.Y(n_13711)
);

AND2x2_ASAP7_75t_L g13712 ( 
.A(n_12787),
.B(n_9852),
.Y(n_13712)
);

INVx2_ASAP7_75t_L g13713 ( 
.A(n_12980),
.Y(n_13713)
);

BUFx3_ASAP7_75t_L g13714 ( 
.A(n_12402),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_13083),
.Y(n_13715)
);

AND2x4_ASAP7_75t_L g13716 ( 
.A(n_12642),
.B(n_12064),
.Y(n_13716)
);

INVx1_ASAP7_75t_L g13717 ( 
.A(n_13095),
.Y(n_13717)
);

AND2x2_ASAP7_75t_L g13718 ( 
.A(n_12791),
.B(n_9852),
.Y(n_13718)
);

INVx1_ASAP7_75t_L g13719 ( 
.A(n_13121),
.Y(n_13719)
);

INVx2_ASAP7_75t_L g13720 ( 
.A(n_12981),
.Y(n_13720)
);

INVx1_ASAP7_75t_L g13721 ( 
.A(n_13131),
.Y(n_13721)
);

AND2x2_ASAP7_75t_L g13722 ( 
.A(n_12798),
.B(n_12801),
.Y(n_13722)
);

NAND2xp5_ASAP7_75t_L g13723 ( 
.A(n_13084),
.B(n_11247),
.Y(n_13723)
);

INVx2_ASAP7_75t_L g13724 ( 
.A(n_12988),
.Y(n_13724)
);

INVx1_ASAP7_75t_L g13725 ( 
.A(n_13154),
.Y(n_13725)
);

HB1xp67_ASAP7_75t_L g13726 ( 
.A(n_13011),
.Y(n_13726)
);

INVx2_ASAP7_75t_L g13727 ( 
.A(n_13021),
.Y(n_13727)
);

INVx2_ASAP7_75t_L g13728 ( 
.A(n_13038),
.Y(n_13728)
);

AND2x2_ASAP7_75t_L g13729 ( 
.A(n_12811),
.B(n_9860),
.Y(n_13729)
);

INVx1_ASAP7_75t_L g13730 ( 
.A(n_13160),
.Y(n_13730)
);

INVx2_ASAP7_75t_L g13731 ( 
.A(n_13279),
.Y(n_13731)
);

AOI21xp33_ASAP7_75t_SL g13732 ( 
.A1(n_12458),
.A2(n_11770),
.B(n_11095),
.Y(n_13732)
);

AND2x4_ASAP7_75t_L g13733 ( 
.A(n_12642),
.B(n_12596),
.Y(n_13733)
);

INVx2_ASAP7_75t_L g13734 ( 
.A(n_13279),
.Y(n_13734)
);

AOI22xp33_ASAP7_75t_L g13735 ( 
.A1(n_12492),
.A2(n_11405),
.B1(n_11350),
.B2(n_8813),
.Y(n_13735)
);

AO21x2_ASAP7_75t_L g13736 ( 
.A1(n_12371),
.A2(n_11212),
.B(n_11211),
.Y(n_13736)
);

OR2x6_ASAP7_75t_L g13737 ( 
.A(n_12477),
.B(n_7777),
.Y(n_13737)
);

INVx1_ASAP7_75t_L g13738 ( 
.A(n_13180),
.Y(n_13738)
);

AND2x2_ASAP7_75t_L g13739 ( 
.A(n_12818),
.B(n_9860),
.Y(n_13739)
);

HB1xp67_ASAP7_75t_L g13740 ( 
.A(n_12765),
.Y(n_13740)
);

INVx3_ASAP7_75t_L g13741 ( 
.A(n_13102),
.Y(n_13741)
);

INVx1_ASAP7_75t_L g13742 ( 
.A(n_13194),
.Y(n_13742)
);

HB1xp67_ASAP7_75t_L g13743 ( 
.A(n_12585),
.Y(n_13743)
);

INVx1_ASAP7_75t_L g13744 ( 
.A(n_13204),
.Y(n_13744)
);

INVx1_ASAP7_75t_L g13745 ( 
.A(n_13221),
.Y(n_13745)
);

AND2x4_ASAP7_75t_L g13746 ( 
.A(n_12596),
.B(n_12064),
.Y(n_13746)
);

INVx2_ASAP7_75t_SL g13747 ( 
.A(n_12593),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_12846),
.B(n_9926),
.Y(n_13748)
);

AND2x2_ASAP7_75t_L g13749 ( 
.A(n_12861),
.B(n_9926),
.Y(n_13749)
);

HB1xp67_ASAP7_75t_L g13750 ( 
.A(n_12687),
.Y(n_13750)
);

AND2x2_ASAP7_75t_L g13751 ( 
.A(n_12887),
.B(n_9959),
.Y(n_13751)
);

HB1xp67_ASAP7_75t_L g13752 ( 
.A(n_12690),
.Y(n_13752)
);

INVx1_ASAP7_75t_L g13753 ( 
.A(n_13246),
.Y(n_13753)
);

NOR2xp33_ASAP7_75t_L g13754 ( 
.A(n_12528),
.B(n_10230),
.Y(n_13754)
);

AND2x2_ASAP7_75t_L g13755 ( 
.A(n_13018),
.B(n_9959),
.Y(n_13755)
);

HB1xp67_ASAP7_75t_L g13756 ( 
.A(n_12703),
.Y(n_13756)
);

HB1xp67_ASAP7_75t_L g13757 ( 
.A(n_12713),
.Y(n_13757)
);

INVx2_ASAP7_75t_L g13758 ( 
.A(n_13279),
.Y(n_13758)
);

AND2x2_ASAP7_75t_L g13759 ( 
.A(n_13212),
.B(n_9963),
.Y(n_13759)
);

INVx1_ASAP7_75t_L g13760 ( 
.A(n_13259),
.Y(n_13760)
);

HB1xp67_ASAP7_75t_L g13761 ( 
.A(n_12715),
.Y(n_13761)
);

AND2x4_ASAP7_75t_SL g13762 ( 
.A(n_12570),
.B(n_8063),
.Y(n_13762)
);

AND2x2_ASAP7_75t_L g13763 ( 
.A(n_12724),
.B(n_9963),
.Y(n_13763)
);

NAND2xp5_ASAP7_75t_L g13764 ( 
.A(n_12305),
.B(n_12512),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_13269),
.Y(n_13765)
);

AND2x2_ASAP7_75t_L g13766 ( 
.A(n_12724),
.B(n_10042),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_13270),
.Y(n_13767)
);

INVx2_ASAP7_75t_L g13768 ( 
.A(n_12594),
.Y(n_13768)
);

AND2x2_ASAP7_75t_L g13769 ( 
.A(n_13245),
.B(n_10042),
.Y(n_13769)
);

NAND2xp5_ASAP7_75t_L g13770 ( 
.A(n_12595),
.B(n_11250),
.Y(n_13770)
);

OR2x2_ASAP7_75t_L g13771 ( 
.A(n_12681),
.B(n_10091),
.Y(n_13771)
);

AND2x4_ASAP7_75t_L g13772 ( 
.A(n_12635),
.B(n_9277),
.Y(n_13772)
);

AND2x2_ASAP7_75t_L g13773 ( 
.A(n_12971),
.B(n_10047),
.Y(n_13773)
);

INVx1_ASAP7_75t_L g13774 ( 
.A(n_13287),
.Y(n_13774)
);

AND2x4_ASAP7_75t_L g13775 ( 
.A(n_12635),
.B(n_9277),
.Y(n_13775)
);

INVx1_ASAP7_75t_L g13776 ( 
.A(n_13249),
.Y(n_13776)
);

AND2x2_ASAP7_75t_L g13777 ( 
.A(n_13235),
.B(n_10047),
.Y(n_13777)
);

OAI22xp5_ASAP7_75t_L g13778 ( 
.A1(n_12423),
.A2(n_8239),
.B1(n_8326),
.B2(n_8204),
.Y(n_13778)
);

INVx1_ASAP7_75t_L g13779 ( 
.A(n_13169),
.Y(n_13779)
);

INVx1_ASAP7_75t_L g13780 ( 
.A(n_13186),
.Y(n_13780)
);

INVx3_ASAP7_75t_L g13781 ( 
.A(n_13196),
.Y(n_13781)
);

INVx1_ASAP7_75t_L g13782 ( 
.A(n_13214),
.Y(n_13782)
);

INVx1_ASAP7_75t_L g13783 ( 
.A(n_13133),
.Y(n_13783)
);

INVx1_ASAP7_75t_L g13784 ( 
.A(n_12617),
.Y(n_13784)
);

OR2x2_ASAP7_75t_L g13785 ( 
.A(n_12996),
.B(n_10091),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_12310),
.Y(n_13786)
);

BUFx3_ASAP7_75t_L g13787 ( 
.A(n_12991),
.Y(n_13787)
);

HB1xp67_ASAP7_75t_L g13788 ( 
.A(n_12719),
.Y(n_13788)
);

AND2x2_ASAP7_75t_L g13789 ( 
.A(n_12314),
.B(n_10107),
.Y(n_13789)
);

INVx2_ASAP7_75t_L g13790 ( 
.A(n_12594),
.Y(n_13790)
);

INVx2_ASAP7_75t_L g13791 ( 
.A(n_12614),
.Y(n_13791)
);

AND2x2_ASAP7_75t_L g13792 ( 
.A(n_12335),
.B(n_10107),
.Y(n_13792)
);

HB1xp67_ASAP7_75t_L g13793 ( 
.A(n_12742),
.Y(n_13793)
);

AND2x2_ASAP7_75t_L g13794 ( 
.A(n_12340),
.B(n_10224),
.Y(n_13794)
);

AND2x2_ASAP7_75t_L g13795 ( 
.A(n_12353),
.B(n_10224),
.Y(n_13795)
);

INVx3_ASAP7_75t_L g13796 ( 
.A(n_13196),
.Y(n_13796)
);

INVx1_ASAP7_75t_L g13797 ( 
.A(n_12310),
.Y(n_13797)
);

INVx2_ASAP7_75t_L g13798 ( 
.A(n_12614),
.Y(n_13798)
);

INVx2_ASAP7_75t_L g13799 ( 
.A(n_12614),
.Y(n_13799)
);

AND2x2_ASAP7_75t_L g13800 ( 
.A(n_12437),
.B(n_11979),
.Y(n_13800)
);

INVx1_ASAP7_75t_L g13801 ( 
.A(n_13055),
.Y(n_13801)
);

HB1xp67_ASAP7_75t_L g13802 ( 
.A(n_12745),
.Y(n_13802)
);

AND2x2_ASAP7_75t_L g13803 ( 
.A(n_12517),
.B(n_11979),
.Y(n_13803)
);

AND2x2_ASAP7_75t_L g13804 ( 
.A(n_12560),
.B(n_11979),
.Y(n_13804)
);

INVxp67_ASAP7_75t_SL g13805 ( 
.A(n_12718),
.Y(n_13805)
);

INVx1_ASAP7_75t_L g13806 ( 
.A(n_13101),
.Y(n_13806)
);

INVx1_ASAP7_75t_SL g13807 ( 
.A(n_13175),
.Y(n_13807)
);

INVx1_ASAP7_75t_L g13808 ( 
.A(n_12503),
.Y(n_13808)
);

BUFx2_ASAP7_75t_SL g13809 ( 
.A(n_12411),
.Y(n_13809)
);

AOI22xp33_ASAP7_75t_SL g13810 ( 
.A1(n_12313),
.A2(n_12093),
.B1(n_12011),
.B2(n_11740),
.Y(n_13810)
);

OR2x2_ASAP7_75t_L g13811 ( 
.A(n_12581),
.B(n_10092),
.Y(n_13811)
);

BUFx3_ASAP7_75t_L g13812 ( 
.A(n_13200),
.Y(n_13812)
);

NAND2xp5_ASAP7_75t_L g13813 ( 
.A(n_12479),
.B(n_11257),
.Y(n_13813)
);

AND2x4_ASAP7_75t_L g13814 ( 
.A(n_12733),
.B(n_9277),
.Y(n_13814)
);

INVx2_ASAP7_75t_L g13815 ( 
.A(n_13080),
.Y(n_13815)
);

AOI22xp33_ASAP7_75t_L g13816 ( 
.A1(n_12365),
.A2(n_11405),
.B1(n_11350),
.B2(n_8813),
.Y(n_13816)
);

INVx2_ASAP7_75t_L g13817 ( 
.A(n_13080),
.Y(n_13817)
);

NAND2xp5_ASAP7_75t_L g13818 ( 
.A(n_12504),
.B(n_11259),
.Y(n_13818)
);

AOI22xp33_ASAP7_75t_L g13819 ( 
.A1(n_12338),
.A2(n_11405),
.B1(n_11350),
.B2(n_8813),
.Y(n_13819)
);

INVx1_ASAP7_75t_L g13820 ( 
.A(n_13103),
.Y(n_13820)
);

AND2x2_ASAP7_75t_L g13821 ( 
.A(n_12583),
.B(n_10247),
.Y(n_13821)
);

INVx1_ASAP7_75t_L g13822 ( 
.A(n_13109),
.Y(n_13822)
);

INVx1_ASAP7_75t_L g13823 ( 
.A(n_13116),
.Y(n_13823)
);

AND2x2_ASAP7_75t_L g13824 ( 
.A(n_12507),
.B(n_12515),
.Y(n_13824)
);

INVx1_ASAP7_75t_L g13825 ( 
.A(n_13126),
.Y(n_13825)
);

INVx2_ASAP7_75t_L g13826 ( 
.A(n_13041),
.Y(n_13826)
);

AND2x2_ASAP7_75t_L g13827 ( 
.A(n_12507),
.B(n_10247),
.Y(n_13827)
);

INVxp67_ASAP7_75t_L g13828 ( 
.A(n_13295),
.Y(n_13828)
);

NAND2xp5_ASAP7_75t_L g13829 ( 
.A(n_12329),
.B(n_11260),
.Y(n_13829)
);

INVx2_ASAP7_75t_L g13830 ( 
.A(n_13114),
.Y(n_13830)
);

INVx2_ASAP7_75t_SL g13831 ( 
.A(n_12650),
.Y(n_13831)
);

INVx3_ASAP7_75t_L g13832 ( 
.A(n_13256),
.Y(n_13832)
);

NAND2xp5_ASAP7_75t_L g13833 ( 
.A(n_12328),
.B(n_11261),
.Y(n_13833)
);

INVx1_ASAP7_75t_L g13834 ( 
.A(n_13161),
.Y(n_13834)
);

NOR2x1p5_ASAP7_75t_L g13835 ( 
.A(n_13122),
.B(n_10434),
.Y(n_13835)
);

AND2x2_ASAP7_75t_L g13836 ( 
.A(n_12515),
.B(n_10338),
.Y(n_13836)
);

INVx3_ASAP7_75t_L g13837 ( 
.A(n_13256),
.Y(n_13837)
);

BUFx2_ASAP7_75t_L g13838 ( 
.A(n_12889),
.Y(n_13838)
);

OR2x2_ASAP7_75t_L g13839 ( 
.A(n_12794),
.B(n_10092),
.Y(n_13839)
);

AND2x2_ASAP7_75t_L g13840 ( 
.A(n_12545),
.B(n_10960),
.Y(n_13840)
);

INVx2_ASAP7_75t_L g13841 ( 
.A(n_13114),
.Y(n_13841)
);

INVx1_ASAP7_75t_L g13842 ( 
.A(n_13197),
.Y(n_13842)
);

NAND2xp5_ASAP7_75t_L g13843 ( 
.A(n_12559),
.B(n_11264),
.Y(n_13843)
);

AOI22xp33_ASAP7_75t_L g13844 ( 
.A1(n_12294),
.A2(n_8813),
.B1(n_8905),
.B2(n_8799),
.Y(n_13844)
);

NAND2xp5_ASAP7_75t_L g13845 ( 
.A(n_12356),
.B(n_11267),
.Y(n_13845)
);

AND2x2_ASAP7_75t_L g13846 ( 
.A(n_12545),
.B(n_10960),
.Y(n_13846)
);

AND2x2_ASAP7_75t_L g13847 ( 
.A(n_12558),
.B(n_9936),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_13203),
.Y(n_13848)
);

AND2x2_ASAP7_75t_L g13849 ( 
.A(n_12558),
.B(n_9965),
.Y(n_13849)
);

HB1xp67_ASAP7_75t_L g13850 ( 
.A(n_12748),
.Y(n_13850)
);

OR2x2_ASAP7_75t_L g13851 ( 
.A(n_12803),
.B(n_11270),
.Y(n_13851)
);

NOR2x1_ASAP7_75t_L g13852 ( 
.A(n_13148),
.B(n_9500),
.Y(n_13852)
);

AND2x2_ASAP7_75t_L g13853 ( 
.A(n_12733),
.B(n_9965),
.Y(n_13853)
);

INVx2_ASAP7_75t_L g13854 ( 
.A(n_13114),
.Y(n_13854)
);

AND2x2_ASAP7_75t_L g13855 ( 
.A(n_12736),
.B(n_9977),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_12736),
.B(n_9977),
.Y(n_13856)
);

INVx1_ASAP7_75t_L g13857 ( 
.A(n_13206),
.Y(n_13857)
);

NAND2xp5_ASAP7_75t_L g13858 ( 
.A(n_13277),
.B(n_11272),
.Y(n_13858)
);

HB1xp67_ASAP7_75t_L g13859 ( 
.A(n_12671),
.Y(n_13859)
);

BUFx2_ASAP7_75t_L g13860 ( 
.A(n_12962),
.Y(n_13860)
);

INVx1_ASAP7_75t_L g13861 ( 
.A(n_13219),
.Y(n_13861)
);

INVx1_ASAP7_75t_L g13862 ( 
.A(n_13226),
.Y(n_13862)
);

HB1xp67_ASAP7_75t_L g13863 ( 
.A(n_12671),
.Y(n_13863)
);

INVx2_ASAP7_75t_L g13864 ( 
.A(n_12761),
.Y(n_13864)
);

AO31x2_ASAP7_75t_L g13865 ( 
.A1(n_13176),
.A2(n_13189),
.A3(n_12519),
.B(n_12394),
.Y(n_13865)
);

OR2x2_ASAP7_75t_L g13866 ( 
.A(n_12844),
.B(n_11273),
.Y(n_13866)
);

INVx1_ASAP7_75t_L g13867 ( 
.A(n_13233),
.Y(n_13867)
);

INVxp67_ASAP7_75t_SL g13868 ( 
.A(n_12336),
.Y(n_13868)
);

AND2x2_ASAP7_75t_L g13869 ( 
.A(n_13019),
.B(n_11770),
.Y(n_13869)
);

AND2x2_ASAP7_75t_L g13870 ( 
.A(n_13049),
.B(n_11818),
.Y(n_13870)
);

NAND2xp5_ASAP7_75t_L g13871 ( 
.A(n_13277),
.B(n_11275),
.Y(n_13871)
);

INVx2_ASAP7_75t_SL g13872 ( 
.A(n_12497),
.Y(n_13872)
);

INVx1_ASAP7_75t_L g13873 ( 
.A(n_13254),
.Y(n_13873)
);

INVx2_ASAP7_75t_L g13874 ( 
.A(n_12270),
.Y(n_13874)
);

OR2x2_ASAP7_75t_L g13875 ( 
.A(n_12987),
.B(n_11278),
.Y(n_13875)
);

INVx1_ASAP7_75t_L g13876 ( 
.A(n_13260),
.Y(n_13876)
);

AND2x2_ASAP7_75t_L g13877 ( 
.A(n_13063),
.B(n_11818),
.Y(n_13877)
);

HB1xp67_ASAP7_75t_L g13878 ( 
.A(n_12671),
.Y(n_13878)
);

BUFx2_ASAP7_75t_L g13879 ( 
.A(n_12962),
.Y(n_13879)
);

HB1xp67_ASAP7_75t_L g13880 ( 
.A(n_13213),
.Y(n_13880)
);

INVx2_ASAP7_75t_L g13881 ( 
.A(n_13145),
.Y(n_13881)
);

AND2x2_ASAP7_75t_L g13882 ( 
.A(n_13073),
.B(n_10554),
.Y(n_13882)
);

INVx1_ASAP7_75t_L g13883 ( 
.A(n_13268),
.Y(n_13883)
);

BUFx2_ASAP7_75t_L g13884 ( 
.A(n_12746),
.Y(n_13884)
);

INVx1_ASAP7_75t_L g13885 ( 
.A(n_13291),
.Y(n_13885)
);

INVx2_ASAP7_75t_L g13886 ( 
.A(n_13284),
.Y(n_13886)
);

NAND2xp5_ASAP7_75t_L g13887 ( 
.A(n_12950),
.B(n_11280),
.Y(n_13887)
);

AOI21xp33_ASAP7_75t_SL g13888 ( 
.A1(n_12424),
.A2(n_10568),
.B(n_7570),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13117),
.B(n_10965),
.Y(n_13889)
);

AND2x2_ASAP7_75t_L g13890 ( 
.A(n_13250),
.B(n_10965),
.Y(n_13890)
);

AND2x4_ASAP7_75t_L g13891 ( 
.A(n_12870),
.B(n_9500),
.Y(n_13891)
);

NAND2xp5_ASAP7_75t_L g13892 ( 
.A(n_13297),
.B(n_11282),
.Y(n_13892)
);

INVx2_ASAP7_75t_L g13893 ( 
.A(n_12383),
.Y(n_13893)
);

BUFx2_ASAP7_75t_L g13894 ( 
.A(n_12746),
.Y(n_13894)
);

NOR2x1_ASAP7_75t_R g13895 ( 
.A(n_12331),
.B(n_7777),
.Y(n_13895)
);

OR2x2_ASAP7_75t_L g13896 ( 
.A(n_13001),
.B(n_11285),
.Y(n_13896)
);

INVx2_ASAP7_75t_SL g13897 ( 
.A(n_12497),
.Y(n_13897)
);

INVx1_ASAP7_75t_L g13898 ( 
.A(n_13304),
.Y(n_13898)
);

INVx1_ASAP7_75t_L g13899 ( 
.A(n_13307),
.Y(n_13899)
);

BUFx3_ASAP7_75t_L g13900 ( 
.A(n_12460),
.Y(n_13900)
);

INVx1_ASAP7_75t_L g13901 ( 
.A(n_12295),
.Y(n_13901)
);

NAND2xp5_ASAP7_75t_L g13902 ( 
.A(n_13216),
.B(n_11291),
.Y(n_13902)
);

INVx2_ASAP7_75t_L g13903 ( 
.A(n_12388),
.Y(n_13903)
);

HB1xp67_ASAP7_75t_L g13904 ( 
.A(n_12997),
.Y(n_13904)
);

BUFx3_ASAP7_75t_L g13905 ( 
.A(n_12460),
.Y(n_13905)
);

BUFx3_ASAP7_75t_L g13906 ( 
.A(n_12785),
.Y(n_13906)
);

INVx2_ASAP7_75t_L g13907 ( 
.A(n_12621),
.Y(n_13907)
);

INVx2_ASAP7_75t_L g13908 ( 
.A(n_12621),
.Y(n_13908)
);

INVx1_ASAP7_75t_L g13909 ( 
.A(n_13037),
.Y(n_13909)
);

AND2x2_ASAP7_75t_L g13910 ( 
.A(n_13266),
.B(n_11013),
.Y(n_13910)
);

NAND2xp5_ASAP7_75t_L g13911 ( 
.A(n_12624),
.B(n_11292),
.Y(n_13911)
);

AND2x2_ASAP7_75t_L g13912 ( 
.A(n_13288),
.B(n_11013),
.Y(n_13912)
);

AND2x4_ASAP7_75t_L g13913 ( 
.A(n_12411),
.B(n_9500),
.Y(n_13913)
);

OR2x2_ASAP7_75t_L g13914 ( 
.A(n_13006),
.B(n_11293),
.Y(n_13914)
);

AND2x2_ASAP7_75t_L g13915 ( 
.A(n_12331),
.B(n_11017),
.Y(n_13915)
);

INVx2_ASAP7_75t_L g13916 ( 
.A(n_12688),
.Y(n_13916)
);

AND2x2_ASAP7_75t_L g13917 ( 
.A(n_12470),
.B(n_11017),
.Y(n_13917)
);

AND2x2_ASAP7_75t_L g13918 ( 
.A(n_12470),
.B(n_11796),
.Y(n_13918)
);

AND2x2_ASAP7_75t_L g13919 ( 
.A(n_13190),
.B(n_11796),
.Y(n_13919)
);

INVx1_ASAP7_75t_L g13920 ( 
.A(n_12389),
.Y(n_13920)
);

AND2x2_ASAP7_75t_L g13921 ( 
.A(n_13215),
.B(n_11796),
.Y(n_13921)
);

AND2x2_ASAP7_75t_L g13922 ( 
.A(n_13234),
.B(n_11796),
.Y(n_13922)
);

BUFx2_ASAP7_75t_L g13923 ( 
.A(n_12746),
.Y(n_13923)
);

OR2x2_ASAP7_75t_L g13924 ( 
.A(n_12706),
.B(n_11303),
.Y(n_13924)
);

AND2x2_ASAP7_75t_L g13925 ( 
.A(n_12411),
.B(n_12055),
.Y(n_13925)
);

INVx4_ASAP7_75t_L g13926 ( 
.A(n_12785),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_13099),
.Y(n_13927)
);

AND2x2_ASAP7_75t_L g13928 ( 
.A(n_12700),
.B(n_12055),
.Y(n_13928)
);

NAND2xp5_ASAP7_75t_L g13929 ( 
.A(n_12649),
.B(n_12646),
.Y(n_13929)
);

BUFx2_ASAP7_75t_L g13930 ( 
.A(n_12746),
.Y(n_13930)
);

HB1xp67_ASAP7_75t_L g13931 ( 
.A(n_13252),
.Y(n_13931)
);

NOR2xp33_ASAP7_75t_L g13932 ( 
.A(n_13044),
.B(n_10618),
.Y(n_13932)
);

INVx2_ASAP7_75t_L g13933 ( 
.A(n_12850),
.Y(n_13933)
);

NOR2x1_ASAP7_75t_L g13934 ( 
.A(n_13097),
.B(n_9500),
.Y(n_13934)
);

INVx1_ASAP7_75t_L g13935 ( 
.A(n_13123),
.Y(n_13935)
);

INVx1_ASAP7_75t_L g13936 ( 
.A(n_12568),
.Y(n_13936)
);

AND2x2_ASAP7_75t_L g13937 ( 
.A(n_12700),
.B(n_12055),
.Y(n_13937)
);

HB1xp67_ASAP7_75t_L g13938 ( 
.A(n_12848),
.Y(n_13938)
);

INVx4_ASAP7_75t_L g13939 ( 
.A(n_12860),
.Y(n_13939)
);

AND2x2_ASAP7_75t_L g13940 ( 
.A(n_12860),
.B(n_12055),
.Y(n_13940)
);

AND2x2_ASAP7_75t_L g13941 ( 
.A(n_12911),
.B(n_10725),
.Y(n_13941)
);

AND2x2_ASAP7_75t_L g13942 ( 
.A(n_12762),
.B(n_10725),
.Y(n_13942)
);

NAND2xp5_ASAP7_75t_L g13943 ( 
.A(n_12427),
.B(n_11304),
.Y(n_13943)
);

INVx2_ASAP7_75t_L g13944 ( 
.A(n_12850),
.Y(n_13944)
);

BUFx6f_ASAP7_75t_L g13945 ( 
.A(n_12852),
.Y(n_13945)
);

INVx1_ASAP7_75t_L g13946 ( 
.A(n_12471),
.Y(n_13946)
);

INVx3_ASAP7_75t_L g13947 ( 
.A(n_12852),
.Y(n_13947)
);

INVx1_ASAP7_75t_L g13948 ( 
.A(n_12471),
.Y(n_13948)
);

AND2x2_ASAP7_75t_L g13949 ( 
.A(n_12774),
.B(n_10765),
.Y(n_13949)
);

INVx1_ASAP7_75t_L g13950 ( 
.A(n_13060),
.Y(n_13950)
);

AND2x2_ASAP7_75t_L g13951 ( 
.A(n_12776),
.B(n_10765),
.Y(n_13951)
);

INVx3_ASAP7_75t_L g13952 ( 
.A(n_12781),
.Y(n_13952)
);

INVx2_ASAP7_75t_L g13953 ( 
.A(n_12850),
.Y(n_13953)
);

NAND2xp5_ASAP7_75t_L g13954 ( 
.A(n_12599),
.B(n_11309),
.Y(n_13954)
);

AND2x2_ASAP7_75t_L g13955 ( 
.A(n_12796),
.B(n_10770),
.Y(n_13955)
);

AND2x2_ASAP7_75t_L g13956 ( 
.A(n_13147),
.B(n_10770),
.Y(n_13956)
);

OR2x2_ASAP7_75t_L g13957 ( 
.A(n_12759),
.B(n_11312),
.Y(n_13957)
);

INVx2_ASAP7_75t_L g13958 ( 
.A(n_12937),
.Y(n_13958)
);

OR2x6_ASAP7_75t_L g13959 ( 
.A(n_12915),
.B(n_7788),
.Y(n_13959)
);

AND2x2_ASAP7_75t_L g13960 ( 
.A(n_13150),
.B(n_10776),
.Y(n_13960)
);

HB1xp67_ASAP7_75t_L g13961 ( 
.A(n_12867),
.Y(n_13961)
);

AND2x2_ASAP7_75t_L g13962 ( 
.A(n_12831),
.B(n_10776),
.Y(n_13962)
);

INVx2_ASAP7_75t_L g13963 ( 
.A(n_12937),
.Y(n_13963)
);

AND2x4_ASAP7_75t_SL g13964 ( 
.A(n_13047),
.B(n_7840),
.Y(n_13964)
);

BUFx2_ASAP7_75t_L g13965 ( 
.A(n_13130),
.Y(n_13965)
);

AND2x2_ASAP7_75t_L g13966 ( 
.A(n_12832),
.B(n_10796),
.Y(n_13966)
);

INVx1_ASAP7_75t_L g13967 ( 
.A(n_13065),
.Y(n_13967)
);

INVx2_ASAP7_75t_SL g13968 ( 
.A(n_13130),
.Y(n_13968)
);

AND2x2_ASAP7_75t_L g13969 ( 
.A(n_12842),
.B(n_10796),
.Y(n_13969)
);

INVx2_ASAP7_75t_SL g13970 ( 
.A(n_13130),
.Y(n_13970)
);

AND2x2_ASAP7_75t_L g13971 ( 
.A(n_12845),
.B(n_10821),
.Y(n_13971)
);

INVx1_ASAP7_75t_L g13972 ( 
.A(n_13104),
.Y(n_13972)
);

INVx2_ASAP7_75t_L g13973 ( 
.A(n_12989),
.Y(n_13973)
);

AND2x2_ASAP7_75t_L g13974 ( 
.A(n_12725),
.B(n_10821),
.Y(n_13974)
);

INVx2_ASAP7_75t_L g13975 ( 
.A(n_12989),
.Y(n_13975)
);

NAND2xp5_ASAP7_75t_L g13976 ( 
.A(n_13264),
.B(n_11313),
.Y(n_13976)
);

INVx4_ASAP7_75t_R g13977 ( 
.A(n_12985),
.Y(n_13977)
);

INVx1_ASAP7_75t_L g13978 ( 
.A(n_13118),
.Y(n_13978)
);

NAND2xp5_ASAP7_75t_L g13979 ( 
.A(n_13274),
.B(n_11319),
.Y(n_13979)
);

INVx1_ASAP7_75t_L g13980 ( 
.A(n_13050),
.Y(n_13980)
);

INVx3_ASAP7_75t_L g13981 ( 
.A(n_12878),
.Y(n_13981)
);

AND2x2_ASAP7_75t_L g13982 ( 
.A(n_12756),
.B(n_10835),
.Y(n_13982)
);

INVx1_ASAP7_75t_L g13983 ( 
.A(n_12998),
.Y(n_13983)
);

INVx1_ASAP7_75t_L g13984 ( 
.A(n_12351),
.Y(n_13984)
);

INVx2_ASAP7_75t_L g13985 ( 
.A(n_12268),
.Y(n_13985)
);

AO31x2_ASAP7_75t_L g13986 ( 
.A1(n_12414),
.A2(n_12731),
.A3(n_12712),
.B(n_12571),
.Y(n_13986)
);

AND2x2_ASAP7_75t_L g13987 ( 
.A(n_13009),
.B(n_10835),
.Y(n_13987)
);

AND2x2_ASAP7_75t_L g13988 ( 
.A(n_13013),
.B(n_10856),
.Y(n_13988)
);

INVx2_ASAP7_75t_SL g13989 ( 
.A(n_13130),
.Y(n_13989)
);

INVx1_ASAP7_75t_L g13990 ( 
.A(n_12351),
.Y(n_13990)
);

NAND2xp5_ASAP7_75t_L g13991 ( 
.A(n_12330),
.B(n_11320),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_12817),
.Y(n_13992)
);

BUFx6f_ASAP7_75t_L g13993 ( 
.A(n_12895),
.Y(n_13993)
);

INVx1_ASAP7_75t_L g13994 ( 
.A(n_12951),
.Y(n_13994)
);

INVx2_ASAP7_75t_L g13995 ( 
.A(n_12858),
.Y(n_13995)
);

INVx1_ASAP7_75t_L g13996 ( 
.A(n_12951),
.Y(n_13996)
);

AOI222xp33_ASAP7_75t_SL g13997 ( 
.A1(n_13098),
.A2(n_11565),
.B1(n_11559),
.B2(n_11566),
.C1(n_11563),
.C2(n_11558),
.Y(n_13997)
);

INVx1_ASAP7_75t_L g13998 ( 
.A(n_12951),
.Y(n_13998)
);

INVx3_ASAP7_75t_L g13999 ( 
.A(n_12939),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_12726),
.B(n_11327),
.Y(n_14000)
);

INVx3_ASAP7_75t_L g14001 ( 
.A(n_12871),
.Y(n_14001)
);

AOI22xp33_ASAP7_75t_L g14002 ( 
.A1(n_13115),
.A2(n_8813),
.B1(n_8905),
.B2(n_8799),
.Y(n_14002)
);

NAND2xp5_ASAP7_75t_L g14003 ( 
.A(n_12730),
.B(n_11330),
.Y(n_14003)
);

AND2x2_ASAP7_75t_L g14004 ( 
.A(n_13091),
.B(n_10856),
.Y(n_14004)
);

AND2x2_ASAP7_75t_L g14005 ( 
.A(n_13120),
.B(n_10873),
.Y(n_14005)
);

INVx2_ASAP7_75t_L g14006 ( 
.A(n_12538),
.Y(n_14006)
);

OR2x2_ASAP7_75t_SL g14007 ( 
.A(n_12481),
.B(n_9578),
.Y(n_14007)
);

OR2x2_ASAP7_75t_L g14008 ( 
.A(n_12784),
.B(n_12804),
.Y(n_14008)
);

AND2x2_ASAP7_75t_L g14009 ( 
.A(n_13146),
.B(n_10873),
.Y(n_14009)
);

AOI22xp33_ASAP7_75t_L g14010 ( 
.A1(n_12472),
.A2(n_8905),
.B1(n_8799),
.B2(n_11211),
.Y(n_14010)
);

HB1xp67_ASAP7_75t_L g14011 ( 
.A(n_12869),
.Y(n_14011)
);

BUFx3_ASAP7_75t_L g14012 ( 
.A(n_13210),
.Y(n_14012)
);

HB1xp67_ASAP7_75t_L g14013 ( 
.A(n_13036),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_12536),
.Y(n_14014)
);

AND2x4_ASAP7_75t_L g14015 ( 
.A(n_13314),
.B(n_10017),
.Y(n_14015)
);

OR2x2_ASAP7_75t_L g14016 ( 
.A(n_12865),
.B(n_11336),
.Y(n_14016)
);

INVx2_ASAP7_75t_L g14017 ( 
.A(n_12538),
.Y(n_14017)
);

INVx2_ASAP7_75t_L g14018 ( 
.A(n_12407),
.Y(n_14018)
);

NOR2xp33_ASAP7_75t_L g14019 ( 
.A(n_13229),
.B(n_10630),
.Y(n_14019)
);

NOR2xp67_ASAP7_75t_L g14020 ( 
.A(n_12573),
.B(n_13217),
.Y(n_14020)
);

INVx1_ASAP7_75t_L g14021 ( 
.A(n_12403),
.Y(n_14021)
);

INVx2_ASAP7_75t_L g14022 ( 
.A(n_13199),
.Y(n_14022)
);

OR2x2_ASAP7_75t_L g14023 ( 
.A(n_12882),
.B(n_11340),
.Y(n_14023)
);

NAND2xp5_ASAP7_75t_L g14024 ( 
.A(n_12732),
.B(n_11348),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_12403),
.Y(n_14025)
);

HB1xp67_ASAP7_75t_L g14026 ( 
.A(n_12940),
.Y(n_14026)
);

INVx1_ASAP7_75t_L g14027 ( 
.A(n_12403),
.Y(n_14027)
);

INVx1_ASAP7_75t_L g14028 ( 
.A(n_12995),
.Y(n_14028)
);

OR2x2_ASAP7_75t_L g14029 ( 
.A(n_12954),
.B(n_11349),
.Y(n_14029)
);

HB1xp67_ASAP7_75t_L g14030 ( 
.A(n_12984),
.Y(n_14030)
);

AND2x2_ASAP7_75t_L g14031 ( 
.A(n_13020),
.B(n_10890),
.Y(n_14031)
);

BUFx3_ASAP7_75t_L g14032 ( 
.A(n_13312),
.Y(n_14032)
);

INVx1_ASAP7_75t_L g14033 ( 
.A(n_12995),
.Y(n_14033)
);

OR2x2_ASAP7_75t_L g14034 ( 
.A(n_13003),
.B(n_11351),
.Y(n_14034)
);

AND2x2_ASAP7_75t_L g14035 ( 
.A(n_13192),
.B(n_10890),
.Y(n_14035)
);

INVx1_ASAP7_75t_L g14036 ( 
.A(n_12995),
.Y(n_14036)
);

INVx2_ASAP7_75t_L g14037 ( 
.A(n_12986),
.Y(n_14037)
);

AND2x2_ASAP7_75t_L g14038 ( 
.A(n_13195),
.B(n_10924),
.Y(n_14038)
);

INVxp67_ASAP7_75t_SL g14039 ( 
.A(n_13089),
.Y(n_14039)
);

INVx1_ASAP7_75t_L g14040 ( 
.A(n_12267),
.Y(n_14040)
);

BUFx3_ASAP7_75t_L g14041 ( 
.A(n_12797),
.Y(n_14041)
);

AND2x2_ASAP7_75t_L g14042 ( 
.A(n_13211),
.B(n_10924),
.Y(n_14042)
);

HB1xp67_ASAP7_75t_L g14043 ( 
.A(n_13033),
.Y(n_14043)
);

NOR2xp33_ASAP7_75t_L g14044 ( 
.A(n_12920),
.B(n_10638),
.Y(n_14044)
);

HB1xp67_ASAP7_75t_L g14045 ( 
.A(n_12644),
.Y(n_14045)
);

AND2x2_ASAP7_75t_L g14046 ( 
.A(n_13224),
.B(n_13231),
.Y(n_14046)
);

NAND2xp5_ASAP7_75t_L g14047 ( 
.A(n_12755),
.B(n_12766),
.Y(n_14047)
);

BUFx2_ASAP7_75t_L g14048 ( 
.A(n_13092),
.Y(n_14048)
);

INVx1_ASAP7_75t_L g14049 ( 
.A(n_12654),
.Y(n_14049)
);

OR2x2_ASAP7_75t_L g14050 ( 
.A(n_12734),
.B(n_11352),
.Y(n_14050)
);

INVx3_ASAP7_75t_L g14051 ( 
.A(n_13078),
.Y(n_14051)
);

AOI22xp33_ASAP7_75t_L g14052 ( 
.A1(n_12288),
.A2(n_8905),
.B1(n_8799),
.B2(n_11212),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13014),
.B(n_10943),
.Y(n_14053)
);

OR2x2_ASAP7_75t_L g14054 ( 
.A(n_12737),
.B(n_11356),
.Y(n_14054)
);

INVx2_ASAP7_75t_L g14055 ( 
.A(n_13070),
.Y(n_14055)
);

AND2x4_ASAP7_75t_L g14056 ( 
.A(n_13111),
.B(n_10065),
.Y(n_14056)
);

AND2x2_ASAP7_75t_L g14057 ( 
.A(n_13247),
.B(n_13168),
.Y(n_14057)
);

INVx2_ASAP7_75t_L g14058 ( 
.A(n_13070),
.Y(n_14058)
);

INVx1_ASAP7_75t_L g14059 ( 
.A(n_12660),
.Y(n_14059)
);

INVx2_ASAP7_75t_L g14060 ( 
.A(n_13071),
.Y(n_14060)
);

INVx1_ASAP7_75t_L g14061 ( 
.A(n_12727),
.Y(n_14061)
);

INVx1_ASAP7_75t_L g14062 ( 
.A(n_12413),
.Y(n_14062)
);

NAND2xp5_ASAP7_75t_L g14063 ( 
.A(n_12770),
.B(n_11358),
.Y(n_14063)
);

INVx2_ASAP7_75t_L g14064 ( 
.A(n_13071),
.Y(n_14064)
);

INVx2_ASAP7_75t_L g14065 ( 
.A(n_13172),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13173),
.B(n_10943),
.Y(n_14066)
);

INVx4_ASAP7_75t_L g14067 ( 
.A(n_13072),
.Y(n_14067)
);

INVx2_ASAP7_75t_L g14068 ( 
.A(n_13201),
.Y(n_14068)
);

OR2x2_ASAP7_75t_L g14069 ( 
.A(n_12598),
.B(n_12618),
.Y(n_14069)
);

INVx1_ASAP7_75t_L g14070 ( 
.A(n_12802),
.Y(n_14070)
);

BUFx3_ASAP7_75t_L g14071 ( 
.A(n_13225),
.Y(n_14071)
);

BUFx2_ASAP7_75t_L g14072 ( 
.A(n_12393),
.Y(n_14072)
);

AND2x4_ASAP7_75t_SL g14073 ( 
.A(n_12944),
.B(n_7840),
.Y(n_14073)
);

INVx1_ASAP7_75t_L g14074 ( 
.A(n_13002),
.Y(n_14074)
);

OR2x2_ASAP7_75t_L g14075 ( 
.A(n_12657),
.B(n_12674),
.Y(n_14075)
);

INVx2_ASAP7_75t_L g14076 ( 
.A(n_13207),
.Y(n_14076)
);

AND2x2_ASAP7_75t_L g14077 ( 
.A(n_13093),
.B(n_10469),
.Y(n_14077)
);

AND2x2_ASAP7_75t_L g14078 ( 
.A(n_13157),
.B(n_10469),
.Y(n_14078)
);

INVx2_ASAP7_75t_L g14079 ( 
.A(n_13208),
.Y(n_14079)
);

AND2x2_ASAP7_75t_L g14080 ( 
.A(n_12676),
.B(n_10492),
.Y(n_14080)
);

INVx2_ASAP7_75t_L g14081 ( 
.A(n_12965),
.Y(n_14081)
);

AO31x2_ASAP7_75t_L g14082 ( 
.A1(n_13239),
.A2(n_11215),
.A3(n_11028),
.B(n_11029),
.Y(n_14082)
);

AND2x2_ASAP7_75t_L g14083 ( 
.A(n_12941),
.B(n_10492),
.Y(n_14083)
);

BUFx2_ASAP7_75t_L g14084 ( 
.A(n_12958),
.Y(n_14084)
);

OR2x2_ASAP7_75t_L g14085 ( 
.A(n_12883),
.B(n_11359),
.Y(n_14085)
);

BUFx3_ASAP7_75t_L g14086 ( 
.A(n_13171),
.Y(n_14086)
);

BUFx2_ASAP7_75t_L g14087 ( 
.A(n_12524),
.Y(n_14087)
);

INVx2_ASAP7_75t_L g14088 ( 
.A(n_13223),
.Y(n_14088)
);

INVx3_ASAP7_75t_L g14089 ( 
.A(n_13223),
.Y(n_14089)
);

INVx2_ASAP7_75t_L g14090 ( 
.A(n_13265),
.Y(n_14090)
);

INVx3_ASAP7_75t_L g14091 ( 
.A(n_13265),
.Y(n_14091)
);

OR2x2_ASAP7_75t_L g14092 ( 
.A(n_12901),
.B(n_11360),
.Y(n_14092)
);

OR2x2_ASAP7_75t_L g14093 ( 
.A(n_12582),
.B(n_11365),
.Y(n_14093)
);

AND2x2_ASAP7_75t_L g14094 ( 
.A(n_13077),
.B(n_10507),
.Y(n_14094)
);

BUFx2_ASAP7_75t_L g14095 ( 
.A(n_12847),
.Y(n_14095)
);

AND2x2_ASAP7_75t_L g14096 ( 
.A(n_13048),
.B(n_10507),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_12319),
.Y(n_14097)
);

INVx1_ASAP7_75t_L g14098 ( 
.A(n_12833),
.Y(n_14098)
);

INVx2_ASAP7_75t_L g14099 ( 
.A(n_13068),
.Y(n_14099)
);

INVx4_ASAP7_75t_L g14100 ( 
.A(n_12735),
.Y(n_14100)
);

INVxp67_ASAP7_75t_SL g14101 ( 
.A(n_12438),
.Y(n_14101)
);

INVx1_ASAP7_75t_L g14102 ( 
.A(n_12813),
.Y(n_14102)
);

HB1xp67_ASAP7_75t_L g14103 ( 
.A(n_13183),
.Y(n_14103)
);

INVx3_ASAP7_75t_L g14104 ( 
.A(n_13202),
.Y(n_14104)
);

OR2x2_ASAP7_75t_L g14105 ( 
.A(n_12355),
.B(n_11367),
.Y(n_14105)
);

NAND2xp5_ASAP7_75t_L g14106 ( 
.A(n_12773),
.B(n_12780),
.Y(n_14106)
);

INVx2_ASAP7_75t_L g14107 ( 
.A(n_13042),
.Y(n_14107)
);

AND2x2_ASAP7_75t_L g14108 ( 
.A(n_12809),
.B(n_10511),
.Y(n_14108)
);

NAND2xp5_ASAP7_75t_L g14109 ( 
.A(n_12788),
.B(n_11372),
.Y(n_14109)
);

BUFx3_ASAP7_75t_L g14110 ( 
.A(n_12959),
.Y(n_14110)
);

NAND2x1p5_ASAP7_75t_L g14111 ( 
.A(n_13209),
.B(n_9318),
.Y(n_14111)
);

OR2x2_ASAP7_75t_L g14112 ( 
.A(n_13285),
.B(n_11373),
.Y(n_14112)
);

HB1xp67_ASAP7_75t_L g14113 ( 
.A(n_13205),
.Y(n_14113)
);

AND2x4_ASAP7_75t_L g14114 ( 
.A(n_12806),
.B(n_10075),
.Y(n_14114)
);

INVx3_ASAP7_75t_L g14115 ( 
.A(n_13313),
.Y(n_14115)
);

INVx2_ASAP7_75t_SL g14116 ( 
.A(n_13155),
.Y(n_14116)
);

INVx2_ASAP7_75t_L g14117 ( 
.A(n_13079),
.Y(n_14117)
);

INVx2_ASAP7_75t_L g14118 ( 
.A(n_13232),
.Y(n_14118)
);

AND2x4_ASAP7_75t_L g14119 ( 
.A(n_13162),
.B(n_10075),
.Y(n_14119)
);

INVxp67_ASAP7_75t_SL g14120 ( 
.A(n_12444),
.Y(n_14120)
);

INVx1_ASAP7_75t_L g14121 ( 
.A(n_12434),
.Y(n_14121)
);

INVx2_ASAP7_75t_L g14122 ( 
.A(n_12743),
.Y(n_14122)
);

INVx3_ASAP7_75t_L g14123 ( 
.A(n_12993),
.Y(n_14123)
);

INVx2_ASAP7_75t_L g14124 ( 
.A(n_12637),
.Y(n_14124)
);

AND2x2_ASAP7_75t_L g14125 ( 
.A(n_13163),
.B(n_10511),
.Y(n_14125)
);

AND2x2_ASAP7_75t_L g14126 ( 
.A(n_13119),
.B(n_10621),
.Y(n_14126)
);

AND2x4_ASAP7_75t_L g14127 ( 
.A(n_13136),
.B(n_10621),
.Y(n_14127)
);

AOI22xp5_ASAP7_75t_L g14128 ( 
.A1(n_12464),
.A2(n_8552),
.B1(n_8550),
.B2(n_12011),
.Y(n_14128)
);

OR2x2_ASAP7_75t_L g14129 ( 
.A(n_12518),
.B(n_11378),
.Y(n_14129)
);

AND2x4_ASAP7_75t_L g14130 ( 
.A(n_13124),
.B(n_10662),
.Y(n_14130)
);

INVx3_ASAP7_75t_L g14131 ( 
.A(n_12682),
.Y(n_14131)
);

INVx1_ASAP7_75t_L g14132 ( 
.A(n_12693),
.Y(n_14132)
);

AND2x2_ASAP7_75t_L g14133 ( 
.A(n_13125),
.B(n_10662),
.Y(n_14133)
);

BUFx6f_ASAP7_75t_L g14134 ( 
.A(n_12790),
.Y(n_14134)
);

INVx1_ASAP7_75t_L g14135 ( 
.A(n_12823),
.Y(n_14135)
);

HB1xp67_ASAP7_75t_L g14136 ( 
.A(n_12630),
.Y(n_14136)
);

INVx1_ASAP7_75t_L g14137 ( 
.A(n_12709),
.Y(n_14137)
);

AND2x2_ASAP7_75t_L g14138 ( 
.A(n_13129),
.B(n_10674),
.Y(n_14138)
);

HB1xp67_ASAP7_75t_L g14139 ( 
.A(n_12639),
.Y(n_14139)
);

INVx2_ASAP7_75t_L g14140 ( 
.A(n_12651),
.Y(n_14140)
);

AND2x2_ASAP7_75t_L g14141 ( 
.A(n_13137),
.B(n_10674),
.Y(n_14141)
);

AND2x2_ASAP7_75t_L g14142 ( 
.A(n_13142),
.B(n_10691),
.Y(n_14142)
);

AND2x2_ASAP7_75t_L g14143 ( 
.A(n_13188),
.B(n_12873),
.Y(n_14143)
);

AND2x2_ASAP7_75t_L g14144 ( 
.A(n_12945),
.B(n_10691),
.Y(n_14144)
);

INVx1_ASAP7_75t_L g14145 ( 
.A(n_12854),
.Y(n_14145)
);

OR2x2_ASAP7_75t_L g14146 ( 
.A(n_13056),
.B(n_11382),
.Y(n_14146)
);

HB1xp67_ASAP7_75t_L g14147 ( 
.A(n_12580),
.Y(n_14147)
);

INVx1_ASAP7_75t_L g14148 ( 
.A(n_12857),
.Y(n_14148)
);

NAND2xp5_ASAP7_75t_L g14149 ( 
.A(n_12789),
.B(n_11383),
.Y(n_14149)
);

AND2x2_ASAP7_75t_L g14150 ( 
.A(n_13008),
.B(n_9836),
.Y(n_14150)
);

AND2x2_ASAP7_75t_L g14151 ( 
.A(n_12875),
.B(n_9836),
.Y(n_14151)
);

NAND2xp5_ASAP7_75t_L g14152 ( 
.A(n_12800),
.B(n_11387),
.Y(n_14152)
);

INVx2_ASAP7_75t_L g14153 ( 
.A(n_13082),
.Y(n_14153)
);

INVx1_ASAP7_75t_L g14154 ( 
.A(n_12760),
.Y(n_14154)
);

AND2x2_ASAP7_75t_L g14155 ( 
.A(n_12684),
.B(n_9837),
.Y(n_14155)
);

OR2x2_ASAP7_75t_L g14156 ( 
.A(n_12401),
.B(n_11390),
.Y(n_14156)
);

INVx1_ASAP7_75t_L g14157 ( 
.A(n_12284),
.Y(n_14157)
);

BUFx3_ASAP7_75t_L g14158 ( 
.A(n_12698),
.Y(n_14158)
);

INVx1_ASAP7_75t_L g14159 ( 
.A(n_12296),
.Y(n_14159)
);

BUFx3_ASAP7_75t_L g14160 ( 
.A(n_12441),
.Y(n_14160)
);

AOI22xp33_ASAP7_75t_L g14161 ( 
.A1(n_12283),
.A2(n_12357),
.B1(n_12525),
.B2(n_12349),
.Y(n_14161)
);

OR2x2_ASAP7_75t_L g14162 ( 
.A(n_12482),
.B(n_11392),
.Y(n_14162)
);

NAND2xp5_ASAP7_75t_L g14163 ( 
.A(n_12815),
.B(n_11397),
.Y(n_14163)
);

INVx1_ASAP7_75t_L g14164 ( 
.A(n_12317),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_12932),
.Y(n_14165)
);

AOI22xp33_ASAP7_75t_L g14166 ( 
.A1(n_12429),
.A2(n_8905),
.B1(n_8799),
.B2(n_11215),
.Y(n_14166)
);

INVxp67_ASAP7_75t_SL g14167 ( 
.A(n_12602),
.Y(n_14167)
);

INVx2_ASAP7_75t_L g14168 ( 
.A(n_12578),
.Y(n_14168)
);

BUFx3_ASAP7_75t_L g14169 ( 
.A(n_13278),
.Y(n_14169)
);

AOI221xp5_ASAP7_75t_L g14170 ( 
.A1(n_12406),
.A2(n_11029),
.B1(n_11035),
.B2(n_11028),
.C(n_11024),
.Y(n_14170)
);

INVx2_ASAP7_75t_L g14171 ( 
.A(n_12769),
.Y(n_14171)
);

INVx1_ASAP7_75t_L g14172 ( 
.A(n_12955),
.Y(n_14172)
);

INVx3_ASAP7_75t_L g14173 ( 
.A(n_12696),
.Y(n_14173)
);

INVxp67_ASAP7_75t_L g14174 ( 
.A(n_12876),
.Y(n_14174)
);

INVx1_ASAP7_75t_L g14175 ( 
.A(n_12430),
.Y(n_14175)
);

AND2x4_ASAP7_75t_L g14176 ( 
.A(n_13029),
.B(n_10976),
.Y(n_14176)
);

AND2x2_ASAP7_75t_L g14177 ( 
.A(n_12851),
.B(n_9837),
.Y(n_14177)
);

INVx1_ASAP7_75t_L g14178 ( 
.A(n_12436),
.Y(n_14178)
);

AND2x2_ASAP7_75t_L g14179 ( 
.A(n_12358),
.B(n_9884),
.Y(n_14179)
);

BUFx12f_ASAP7_75t_L g14180 ( 
.A(n_13290),
.Y(n_14180)
);

HB1xp67_ASAP7_75t_L g14181 ( 
.A(n_13166),
.Y(n_14181)
);

INVx3_ASAP7_75t_L g14182 ( 
.A(n_12821),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_13088),
.B(n_9884),
.Y(n_14183)
);

OR2x2_ASAP7_75t_L g14184 ( 
.A(n_13007),
.B(n_11403),
.Y(n_14184)
);

NAND2xp5_ASAP7_75t_L g14185 ( 
.A(n_12820),
.B(n_11411),
.Y(n_14185)
);

INVx1_ASAP7_75t_L g14186 ( 
.A(n_13105),
.Y(n_14186)
);

CKINVDCx20_ASAP7_75t_R g14187 ( 
.A(n_13086),
.Y(n_14187)
);

INVx1_ASAP7_75t_L g14188 ( 
.A(n_13113),
.Y(n_14188)
);

OR2x2_ASAP7_75t_L g14189 ( 
.A(n_12764),
.B(n_11414),
.Y(n_14189)
);

INVx2_ASAP7_75t_L g14190 ( 
.A(n_12810),
.Y(n_14190)
);

INVxp67_ASAP7_75t_L g14191 ( 
.A(n_13311),
.Y(n_14191)
);

INVx4_ASAP7_75t_L g14192 ( 
.A(n_13240),
.Y(n_14192)
);

INVx1_ASAP7_75t_L g14193 ( 
.A(n_12638),
.Y(n_14193)
);

CKINVDCx14_ASAP7_75t_R g14194 ( 
.A(n_12445),
.Y(n_14194)
);

INVx1_ASAP7_75t_L g14195 ( 
.A(n_12307),
.Y(n_14195)
);

INVx3_ASAP7_75t_L g14196 ( 
.A(n_12520),
.Y(n_14196)
);

INVx2_ASAP7_75t_L g14197 ( 
.A(n_12620),
.Y(n_14197)
);

INVx2_ASAP7_75t_L g14198 ( 
.A(n_13141),
.Y(n_14198)
);

NAND2xp5_ASAP7_75t_L g14199 ( 
.A(n_12822),
.B(n_11418),
.Y(n_14199)
);

HB1xp67_ASAP7_75t_L g14200 ( 
.A(n_13156),
.Y(n_14200)
);

AND2x2_ASAP7_75t_L g14201 ( 
.A(n_12380),
.B(n_9651),
.Y(n_14201)
);

OR2x2_ASAP7_75t_L g14202 ( 
.A(n_12825),
.B(n_11421),
.Y(n_14202)
);

INVx2_ASAP7_75t_L g14203 ( 
.A(n_12566),
.Y(n_14203)
);

INVx2_ASAP7_75t_L g14204 ( 
.A(n_13272),
.Y(n_14204)
);

INVx1_ASAP7_75t_L g14205 ( 
.A(n_12373),
.Y(n_14205)
);

INVxp67_ASAP7_75t_L g14206 ( 
.A(n_12391),
.Y(n_14206)
);

NAND2xp5_ASAP7_75t_L g14207 ( 
.A(n_12838),
.B(n_12839),
.Y(n_14207)
);

INVx1_ASAP7_75t_L g14208 ( 
.A(n_12306),
.Y(n_14208)
);

INVx1_ASAP7_75t_L g14209 ( 
.A(n_12707),
.Y(n_14209)
);

INVx1_ASAP7_75t_L g14210 ( 
.A(n_12738),
.Y(n_14210)
);

INVx1_ASAP7_75t_L g14211 ( 
.A(n_13034),
.Y(n_14211)
);

AND2x2_ASAP7_75t_L g14212 ( 
.A(n_13251),
.B(n_9651),
.Y(n_14212)
);

AND2x2_ASAP7_75t_L g14213 ( 
.A(n_13178),
.B(n_9672),
.Y(n_14213)
);

AOI22xp33_ASAP7_75t_L g14214 ( 
.A1(n_12691),
.A2(n_11035),
.B1(n_11036),
.B2(n_11024),
.Y(n_14214)
);

HB1xp67_ASAP7_75t_L g14215 ( 
.A(n_12509),
.Y(n_14215)
);

INVx2_ASAP7_75t_L g14216 ( 
.A(n_12723),
.Y(n_14216)
);

AND2x2_ASAP7_75t_L g14217 ( 
.A(n_12494),
.B(n_9672),
.Y(n_14217)
);

AOI22xp33_ASAP7_75t_L g14218 ( 
.A1(n_12290),
.A2(n_12376),
.B1(n_12428),
.B2(n_12613),
.Y(n_14218)
);

AND2x2_ASAP7_75t_L g14219 ( 
.A(n_12534),
.B(n_10150),
.Y(n_14219)
);

NAND2xp5_ASAP7_75t_L g14220 ( 
.A(n_12440),
.B(n_12900),
.Y(n_14220)
);

INVx2_ASAP7_75t_L g14221 ( 
.A(n_13262),
.Y(n_14221)
);

AND2x2_ASAP7_75t_L g14222 ( 
.A(n_12465),
.B(n_10150),
.Y(n_14222)
);

INVx1_ASAP7_75t_L g14223 ( 
.A(n_13046),
.Y(n_14223)
);

INVx3_ASAP7_75t_L g14224 ( 
.A(n_13243),
.Y(n_14224)
);

AOI22xp33_ASAP7_75t_L g14225 ( 
.A1(n_12491),
.A2(n_11043),
.B1(n_11051),
.B2(n_11036),
.Y(n_14225)
);

NOR2xp33_ASAP7_75t_L g14226 ( 
.A(n_13184),
.B(n_10643),
.Y(n_14226)
);

OR2x2_ASAP7_75t_L g14227 ( 
.A(n_12484),
.B(n_11422),
.Y(n_14227)
);

AND2x2_ASAP7_75t_L g14228 ( 
.A(n_13241),
.B(n_10178),
.Y(n_14228)
);

INVx1_ASAP7_75t_L g14229 ( 
.A(n_13052),
.Y(n_14229)
);

INVx1_ASAP7_75t_L g14230 ( 
.A(n_13054),
.Y(n_14230)
);

BUFx3_ASAP7_75t_L g14231 ( 
.A(n_12705),
.Y(n_14231)
);

OR2x2_ASAP7_75t_L g14232 ( 
.A(n_12514),
.B(n_11429),
.Y(n_14232)
);

AND2x2_ASAP7_75t_L g14233 ( 
.A(n_13244),
.B(n_10178),
.Y(n_14233)
);

AND2x4_ASAP7_75t_SL g14234 ( 
.A(n_13286),
.B(n_7908),
.Y(n_14234)
);

OR2x2_ASAP7_75t_L g14235 ( 
.A(n_12399),
.B(n_11433),
.Y(n_14235)
);

OR2x2_ASAP7_75t_L g14236 ( 
.A(n_12511),
.B(n_11435),
.Y(n_14236)
);

INVx2_ASAP7_75t_L g14237 ( 
.A(n_13267),
.Y(n_14237)
);

INVx1_ASAP7_75t_L g14238 ( 
.A(n_13058),
.Y(n_14238)
);

AO31x2_ASAP7_75t_L g14239 ( 
.A1(n_12408),
.A2(n_11051),
.A3(n_11055),
.B(n_11043),
.Y(n_14239)
);

AND2x2_ASAP7_75t_L g14240 ( 
.A(n_12409),
.B(n_10183),
.Y(n_14240)
);

INVx3_ASAP7_75t_L g14241 ( 
.A(n_12601),
.Y(n_14241)
);

AND2x2_ASAP7_75t_L g14242 ( 
.A(n_12680),
.B(n_10183),
.Y(n_14242)
);

INVx1_ASAP7_75t_L g14243 ( 
.A(n_13066),
.Y(n_14243)
);

AND2x2_ASAP7_75t_L g14244 ( 
.A(n_12923),
.B(n_10190),
.Y(n_14244)
);

BUFx3_ASAP7_75t_L g14245 ( 
.A(n_12757),
.Y(n_14245)
);

INVx3_ASAP7_75t_L g14246 ( 
.A(n_13039),
.Y(n_14246)
);

OR2x2_ASAP7_75t_L g14247 ( 
.A(n_12853),
.B(n_11436),
.Y(n_14247)
);

INVx1_ASAP7_75t_L g14248 ( 
.A(n_13067),
.Y(n_14248)
);

AND2x4_ASAP7_75t_L g14249 ( 
.A(n_13107),
.B(n_10976),
.Y(n_14249)
);

INVx1_ASAP7_75t_L g14250 ( 
.A(n_13076),
.Y(n_14250)
);

INVx2_ASAP7_75t_SL g14251 ( 
.A(n_12474),
.Y(n_14251)
);

INVx3_ASAP7_75t_L g14252 ( 
.A(n_13053),
.Y(n_14252)
);

BUFx2_ASAP7_75t_L g14253 ( 
.A(n_12722),
.Y(n_14253)
);

INVx2_ASAP7_75t_L g14254 ( 
.A(n_12611),
.Y(n_14254)
);

INVx1_ASAP7_75t_L g14255 ( 
.A(n_13085),
.Y(n_14255)
);

OR2x2_ASAP7_75t_L g14256 ( 
.A(n_12562),
.B(n_11440),
.Y(n_14256)
);

INVx2_ASAP7_75t_L g14257 ( 
.A(n_12478),
.Y(n_14257)
);

INVx1_ASAP7_75t_L g14258 ( 
.A(n_12392),
.Y(n_14258)
);

AND2x2_ASAP7_75t_L g14259 ( 
.A(n_13289),
.B(n_10190),
.Y(n_14259)
);

INVxp67_ASAP7_75t_SL g14260 ( 
.A(n_12977),
.Y(n_14260)
);

INVx3_ASAP7_75t_L g14261 ( 
.A(n_13112),
.Y(n_14261)
);

INVx2_ASAP7_75t_L g14262 ( 
.A(n_12506),
.Y(n_14262)
);

AND2x2_ASAP7_75t_L g14263 ( 
.A(n_13310),
.B(n_10209),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_12541),
.Y(n_14264)
);

INVx1_ASAP7_75t_L g14265 ( 
.A(n_12547),
.Y(n_14265)
);

INVx1_ASAP7_75t_L g14266 ( 
.A(n_12396),
.Y(n_14266)
);

INVx1_ASAP7_75t_L g14267 ( 
.A(n_12462),
.Y(n_14267)
);

AND2x2_ASAP7_75t_L g14268 ( 
.A(n_13283),
.B(n_10209),
.Y(n_14268)
);

AND2x4_ASAP7_75t_L g14269 ( 
.A(n_13191),
.B(n_10976),
.Y(n_14269)
);

AND2x2_ASAP7_75t_L g14270 ( 
.A(n_13309),
.B(n_10213),
.Y(n_14270)
);

AND2x2_ASAP7_75t_L g14271 ( 
.A(n_13271),
.B(n_10213),
.Y(n_14271)
);

BUFx2_ASAP7_75t_L g14272 ( 
.A(n_13198),
.Y(n_14272)
);

NAND2xp5_ASAP7_75t_L g14273 ( 
.A(n_12893),
.B(n_11441),
.Y(n_14273)
);

AND2x4_ASAP7_75t_L g14274 ( 
.A(n_12904),
.B(n_10976),
.Y(n_14274)
);

INVx2_ASAP7_75t_L g14275 ( 
.A(n_12672),
.Y(n_14275)
);

AND2x2_ASAP7_75t_L g14276 ( 
.A(n_13255),
.B(n_10260),
.Y(n_14276)
);

AND2x2_ASAP7_75t_L g14277 ( 
.A(n_13167),
.B(n_10260),
.Y(n_14277)
);

INVx1_ASAP7_75t_L g14278 ( 
.A(n_12415),
.Y(n_14278)
);

OAI22xp5_ASAP7_75t_L g14279 ( 
.A1(n_12717),
.A2(n_8239),
.B1(n_8326),
.B2(n_8204),
.Y(n_14279)
);

INVx2_ASAP7_75t_L g14280 ( 
.A(n_12673),
.Y(n_14280)
);

INVx2_ASAP7_75t_L g14281 ( 
.A(n_13282),
.Y(n_14281)
);

NAND2xp5_ASAP7_75t_L g14282 ( 
.A(n_12916),
.B(n_11445),
.Y(n_14282)
);

INVx2_ASAP7_75t_L g14283 ( 
.A(n_12749),
.Y(n_14283)
);

NAND2xp5_ASAP7_75t_L g14284 ( 
.A(n_12884),
.B(n_11454),
.Y(n_14284)
);

BUFx2_ASAP7_75t_L g14285 ( 
.A(n_13134),
.Y(n_14285)
);

NAND2xp5_ASAP7_75t_L g14286 ( 
.A(n_12862),
.B(n_11463),
.Y(n_14286)
);

BUFx2_ASAP7_75t_L g14287 ( 
.A(n_12827),
.Y(n_14287)
);

BUFx3_ASAP7_75t_L g14288 ( 
.A(n_12395),
.Y(n_14288)
);

INVx2_ASAP7_75t_L g14289 ( 
.A(n_12421),
.Y(n_14289)
);

NAND2xp5_ASAP7_75t_L g14290 ( 
.A(n_12521),
.B(n_11465),
.Y(n_14290)
);

NAND2xp5_ASAP7_75t_L g14291 ( 
.A(n_13031),
.B(n_11469),
.Y(n_14291)
);

INVx1_ASAP7_75t_L g14292 ( 
.A(n_13100),
.Y(n_14292)
);

INVx2_ASAP7_75t_L g14293 ( 
.A(n_12485),
.Y(n_14293)
);

INVx2_ASAP7_75t_L g14294 ( 
.A(n_12544),
.Y(n_14294)
);

AND2x4_ASAP7_75t_L g14295 ( 
.A(n_12913),
.B(n_10011),
.Y(n_14295)
);

AOI22xp33_ASAP7_75t_L g14296 ( 
.A1(n_13258),
.A2(n_11059),
.B1(n_11061),
.B2(n_11055),
.Y(n_14296)
);

INVx2_ASAP7_75t_SL g14297 ( 
.A(n_13302),
.Y(n_14297)
);

INVx5_ASAP7_75t_L g14298 ( 
.A(n_13027),
.Y(n_14298)
);

AND2x2_ASAP7_75t_L g14299 ( 
.A(n_13275),
.B(n_10290),
.Y(n_14299)
);

INVx2_ASAP7_75t_SL g14300 ( 
.A(n_13328),
.Y(n_14300)
);

AND2x4_ASAP7_75t_L g14301 ( 
.A(n_13339),
.B(n_10675),
.Y(n_14301)
);

OAI22xp5_ASAP7_75t_L g14302 ( 
.A1(n_14123),
.A2(n_12683),
.B1(n_12714),
.B2(n_12679),
.Y(n_14302)
);

AOI22xp5_ASAP7_75t_L g14303 ( 
.A1(n_14123),
.A2(n_12501),
.B1(n_12488),
.B2(n_12653),
.Y(n_14303)
);

AND2x2_ASAP7_75t_L g14304 ( 
.A(n_13384),
.B(n_10690),
.Y(n_14304)
);

BUFx6f_ASAP7_75t_L g14305 ( 
.A(n_13328),
.Y(n_14305)
);

INVx1_ASAP7_75t_L g14306 ( 
.A(n_13665),
.Y(n_14306)
);

INVx2_ASAP7_75t_L g14307 ( 
.A(n_13327),
.Y(n_14307)
);

NOR2x1_ASAP7_75t_SL g14308 ( 
.A(n_14180),
.B(n_7788),
.Y(n_14308)
);

AOI22xp33_ASAP7_75t_L g14309 ( 
.A1(n_13983),
.A2(n_12398),
.B1(n_12332),
.B2(n_12664),
.Y(n_14309)
);

NOR2xp33_ASAP7_75t_L g14310 ( 
.A(n_13328),
.B(n_10756),
.Y(n_14310)
);

INVxp67_ASAP7_75t_SL g14311 ( 
.A(n_13374),
.Y(n_14311)
);

INVxp67_ASAP7_75t_L g14312 ( 
.A(n_13346),
.Y(n_14312)
);

INVx1_ASAP7_75t_L g14313 ( 
.A(n_13671),
.Y(n_14313)
);

INVx1_ASAP7_75t_L g14314 ( 
.A(n_13416),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_13556),
.Y(n_14315)
);

INVx2_ASAP7_75t_L g14316 ( 
.A(n_13345),
.Y(n_14316)
);

NAND2xp5_ASAP7_75t_L g14317 ( 
.A(n_13345),
.B(n_12533),
.Y(n_14317)
);

INVx1_ASAP7_75t_L g14318 ( 
.A(n_13341),
.Y(n_14318)
);

AND2x4_ASAP7_75t_L g14319 ( 
.A(n_13835),
.B(n_7747),
.Y(n_14319)
);

INVx1_ASAP7_75t_L g14320 ( 
.A(n_13341),
.Y(n_14320)
);

OAI22xp5_ASAP7_75t_L g14321 ( 
.A1(n_14298),
.A2(n_12572),
.B1(n_12574),
.B2(n_12859),
.Y(n_14321)
);

OAI22xp5_ASAP7_75t_L g14322 ( 
.A1(n_14298),
.A2(n_12625),
.B1(n_12665),
.B2(n_13140),
.Y(n_14322)
);

AND2x2_ASAP7_75t_L g14323 ( 
.A(n_13399),
.B(n_10290),
.Y(n_14323)
);

INVx2_ASAP7_75t_L g14324 ( 
.A(n_13606),
.Y(n_14324)
);

INVx1_ASAP7_75t_L g14325 ( 
.A(n_13380),
.Y(n_14325)
);

AND2x2_ASAP7_75t_L g14326 ( 
.A(n_13394),
.B(n_10331),
.Y(n_14326)
);

BUFx2_ASAP7_75t_L g14327 ( 
.A(n_14206),
.Y(n_14327)
);

INVx3_ASAP7_75t_L g14328 ( 
.A(n_13433),
.Y(n_14328)
);

BUFx2_ASAP7_75t_L g14329 ( 
.A(n_14298),
.Y(n_14329)
);

INVx2_ASAP7_75t_L g14330 ( 
.A(n_13606),
.Y(n_14330)
);

INVx2_ASAP7_75t_L g14331 ( 
.A(n_13606),
.Y(n_14331)
);

INVx1_ASAP7_75t_L g14332 ( 
.A(n_13380),
.Y(n_14332)
);

AND2x2_ASAP7_75t_L g14333 ( 
.A(n_13344),
.B(n_10331),
.Y(n_14333)
);

INVx1_ASAP7_75t_L g14334 ( 
.A(n_13385),
.Y(n_14334)
);

INVx1_ASAP7_75t_L g14335 ( 
.A(n_13385),
.Y(n_14335)
);

INVx1_ASAP7_75t_L g14336 ( 
.A(n_13388),
.Y(n_14336)
);

AOI22xp5_ASAP7_75t_L g14337 ( 
.A1(n_13983),
.A2(n_13023),
.B1(n_12960),
.B2(n_12386),
.Y(n_14337)
);

INVx2_ASAP7_75t_L g14338 ( 
.A(n_13648),
.Y(n_14338)
);

INVx1_ASAP7_75t_L g14339 ( 
.A(n_13388),
.Y(n_14339)
);

HB1xp67_ASAP7_75t_L g14340 ( 
.A(n_13379),
.Y(n_14340)
);

BUFx3_ASAP7_75t_L g14341 ( 
.A(n_13357),
.Y(n_14341)
);

NAND2x1p5_ASAP7_75t_L g14342 ( 
.A(n_13628),
.B(n_9318),
.Y(n_14342)
);

AOI22xp33_ASAP7_75t_L g14343 ( 
.A1(n_14175),
.A2(n_12263),
.B1(n_12341),
.B2(n_12347),
.Y(n_14343)
);

HB1xp67_ASAP7_75t_L g14344 ( 
.A(n_13386),
.Y(n_14344)
);

INVx2_ASAP7_75t_L g14345 ( 
.A(n_13648),
.Y(n_14345)
);

BUFx2_ASAP7_75t_SL g14346 ( 
.A(n_13330),
.Y(n_14346)
);

NAND2xp5_ASAP7_75t_L g14347 ( 
.A(n_14101),
.B(n_12513),
.Y(n_14347)
);

NAND2xp5_ASAP7_75t_L g14348 ( 
.A(n_13350),
.B(n_12543),
.Y(n_14348)
);

HB1xp67_ASAP7_75t_L g14349 ( 
.A(n_13320),
.Y(n_14349)
);

AND2x2_ASAP7_75t_L g14350 ( 
.A(n_13524),
.B(n_10391),
.Y(n_14350)
);

AND2x2_ASAP7_75t_L g14351 ( 
.A(n_13637),
.B(n_10391),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_13389),
.Y(n_14352)
);

INVx2_ASAP7_75t_L g14353 ( 
.A(n_13648),
.Y(n_14353)
);

AND2x2_ASAP7_75t_L g14354 ( 
.A(n_13318),
.B(n_10454),
.Y(n_14354)
);

NAND2xp5_ASAP7_75t_L g14355 ( 
.A(n_13451),
.B(n_12564),
.Y(n_14355)
);

INVx2_ASAP7_75t_L g14356 ( 
.A(n_13676),
.Y(n_14356)
);

AOI22xp33_ASAP7_75t_L g14357 ( 
.A1(n_14178),
.A2(n_12489),
.B1(n_12493),
.B2(n_12648),
.Y(n_14357)
);

INVx1_ASAP7_75t_L g14358 ( 
.A(n_13389),
.Y(n_14358)
);

NOR2xp33_ASAP7_75t_L g14359 ( 
.A(n_13682),
.B(n_13410),
.Y(n_14359)
);

INVx1_ASAP7_75t_L g14360 ( 
.A(n_13984),
.Y(n_14360)
);

INVx1_ASAP7_75t_L g14361 ( 
.A(n_13984),
.Y(n_14361)
);

INVx1_ASAP7_75t_L g14362 ( 
.A(n_13990),
.Y(n_14362)
);

NAND2xp5_ASAP7_75t_SL g14363 ( 
.A(n_14176),
.B(n_12775),
.Y(n_14363)
);

BUFx3_ASAP7_75t_L g14364 ( 
.A(n_13479),
.Y(n_14364)
);

INVx2_ASAP7_75t_L g14365 ( 
.A(n_13676),
.Y(n_14365)
);

INVx1_ASAP7_75t_L g14366 ( 
.A(n_13990),
.Y(n_14366)
);

INVx1_ASAP7_75t_L g14367 ( 
.A(n_13994),
.Y(n_14367)
);

AND2x2_ASAP7_75t_L g14368 ( 
.A(n_13537),
.B(n_10454),
.Y(n_14368)
);

AOI22xp33_ASAP7_75t_L g14369 ( 
.A1(n_14196),
.A2(n_12627),
.B1(n_12610),
.B2(n_12628),
.Y(n_14369)
);

OR2x2_ASAP7_75t_L g14370 ( 
.A(n_13322),
.B(n_13335),
.Y(n_14370)
);

AND2x2_ASAP7_75t_L g14371 ( 
.A(n_13762),
.B(n_7747),
.Y(n_14371)
);

INVx2_ASAP7_75t_L g14372 ( 
.A(n_13676),
.Y(n_14372)
);

AND2x2_ASAP7_75t_L g14373 ( 
.A(n_13622),
.B(n_13324),
.Y(n_14373)
);

NOR2x1_ASAP7_75t_L g14374 ( 
.A(n_14067),
.B(n_12563),
.Y(n_14374)
);

OAI22xp5_ASAP7_75t_L g14375 ( 
.A1(n_13323),
.A2(n_13144),
.B1(n_13253),
.B2(n_12567),
.Y(n_14375)
);

NAND2xp5_ASAP7_75t_L g14376 ( 
.A(n_13391),
.B(n_13015),
.Y(n_14376)
);

OR2x2_ASAP7_75t_L g14377 ( 
.A(n_13333),
.B(n_11470),
.Y(n_14377)
);

NAND2xp5_ASAP7_75t_L g14378 ( 
.A(n_14196),
.B(n_13025),
.Y(n_14378)
);

AND2x2_ASAP7_75t_L g14379 ( 
.A(n_13443),
.B(n_13329),
.Y(n_14379)
);

INVx1_ASAP7_75t_L g14380 ( 
.A(n_13996),
.Y(n_14380)
);

NOR2xp33_ASAP7_75t_L g14381 ( 
.A(n_13682),
.B(n_7788),
.Y(n_14381)
);

NAND2xp5_ASAP7_75t_L g14382 ( 
.A(n_13904),
.B(n_12863),
.Y(n_14382)
);

NAND2xp5_ASAP7_75t_L g14383 ( 
.A(n_13359),
.B(n_12864),
.Y(n_14383)
);

NAND2xp5_ASAP7_75t_L g14384 ( 
.A(n_13509),
.B(n_12868),
.Y(n_14384)
);

NAND2xp5_ASAP7_75t_L g14385 ( 
.A(n_14131),
.B(n_12872),
.Y(n_14385)
);

OR2x2_ASAP7_75t_L g14386 ( 
.A(n_14062),
.B(n_11474),
.Y(n_14386)
);

AND2x2_ASAP7_75t_L g14387 ( 
.A(n_13710),
.B(n_7826),
.Y(n_14387)
);

AND2x2_ASAP7_75t_L g14388 ( 
.A(n_13342),
.B(n_13390),
.Y(n_14388)
);

INVx4_ASAP7_75t_L g14389 ( 
.A(n_13367),
.Y(n_14389)
);

NAND2xp5_ASAP7_75t_L g14390 ( 
.A(n_14173),
.B(n_12877),
.Y(n_14390)
);

OR2x2_ASAP7_75t_L g14391 ( 
.A(n_14062),
.B(n_11475),
.Y(n_14391)
);

NOR2xp33_ASAP7_75t_L g14392 ( 
.A(n_13363),
.B(n_7788),
.Y(n_14392)
);

INVx1_ASAP7_75t_L g14393 ( 
.A(n_13998),
.Y(n_14393)
);

BUFx2_ASAP7_75t_SL g14394 ( 
.A(n_13812),
.Y(n_14394)
);

NAND2xp5_ASAP7_75t_L g14395 ( 
.A(n_14131),
.B(n_12881),
.Y(n_14395)
);

INVx1_ASAP7_75t_L g14396 ( 
.A(n_13570),
.Y(n_14396)
);

AOI22xp33_ASAP7_75t_L g14397 ( 
.A1(n_14173),
.A2(n_12591),
.B1(n_12605),
.B2(n_12604),
.Y(n_14397)
);

NAND2xp5_ASAP7_75t_L g14398 ( 
.A(n_13477),
.B(n_12897),
.Y(n_14398)
);

INVx1_ASAP7_75t_L g14399 ( 
.A(n_13570),
.Y(n_14399)
);

BUFx3_ASAP7_75t_L g14400 ( 
.A(n_13363),
.Y(n_14400)
);

NOR2xp33_ASAP7_75t_L g14401 ( 
.A(n_13363),
.B(n_7856),
.Y(n_14401)
);

OR2x2_ASAP7_75t_L g14402 ( 
.A(n_14121),
.B(n_11485),
.Y(n_14402)
);

AND2x2_ASAP7_75t_L g14403 ( 
.A(n_13573),
.B(n_7826),
.Y(n_14403)
);

NAND2xp5_ASAP7_75t_L g14404 ( 
.A(n_13353),
.B(n_12902),
.Y(n_14404)
);

INVx2_ASAP7_75t_L g14405 ( 
.A(n_13693),
.Y(n_14405)
);

BUFx2_ASAP7_75t_L g14406 ( 
.A(n_13471),
.Y(n_14406)
);

AND2x2_ASAP7_75t_L g14407 ( 
.A(n_13573),
.B(n_13466),
.Y(n_14407)
);

AND2x2_ASAP7_75t_L g14408 ( 
.A(n_13415),
.B(n_7832),
.Y(n_14408)
);

INVx1_ASAP7_75t_L g14409 ( 
.A(n_13572),
.Y(n_14409)
);

INVx1_ASAP7_75t_L g14410 ( 
.A(n_13572),
.Y(n_14410)
);

INVx1_ASAP7_75t_SL g14411 ( 
.A(n_13638),
.Y(n_14411)
);

AND2x2_ASAP7_75t_L g14412 ( 
.A(n_13824),
.B(n_7832),
.Y(n_14412)
);

AND2x2_ASAP7_75t_L g14413 ( 
.A(n_13471),
.B(n_7861),
.Y(n_14413)
);

OAI221xp5_ASAP7_75t_L g14414 ( 
.A1(n_14260),
.A2(n_12608),
.B1(n_12542),
.B2(n_12532),
.C(n_13230),
.Y(n_14414)
);

INVx2_ASAP7_75t_L g14415 ( 
.A(n_13693),
.Y(n_14415)
);

OR2x2_ASAP7_75t_L g14416 ( 
.A(n_14121),
.B(n_11487),
.Y(n_14416)
);

AND2x2_ASAP7_75t_L g14417 ( 
.A(n_13395),
.B(n_7861),
.Y(n_14417)
);

AND2x2_ASAP7_75t_L g14418 ( 
.A(n_13395),
.B(n_7903),
.Y(n_14418)
);

AND2x2_ASAP7_75t_L g14419 ( 
.A(n_13722),
.B(n_7903),
.Y(n_14419)
);

INVx2_ASAP7_75t_L g14420 ( 
.A(n_13693),
.Y(n_14420)
);

NOR2xp33_ASAP7_75t_L g14421 ( 
.A(n_13409),
.B(n_7856),
.Y(n_14421)
);

AND2x2_ASAP7_75t_L g14422 ( 
.A(n_13680),
.B(n_7907),
.Y(n_14422)
);

AND2x2_ASAP7_75t_L g14423 ( 
.A(n_13685),
.B(n_7907),
.Y(n_14423)
);

HB1xp67_ASAP7_75t_L g14424 ( 
.A(n_13931),
.Y(n_14424)
);

INVx1_ASAP7_75t_L g14425 ( 
.A(n_13574),
.Y(n_14425)
);

INVx1_ASAP7_75t_L g14426 ( 
.A(n_13574),
.Y(n_14426)
);

INVx1_ASAP7_75t_L g14427 ( 
.A(n_13658),
.Y(n_14427)
);

INVx1_ASAP7_75t_L g14428 ( 
.A(n_13658),
.Y(n_14428)
);

INVx1_ASAP7_75t_L g14429 ( 
.A(n_13674),
.Y(n_14429)
);

INVx2_ASAP7_75t_L g14430 ( 
.A(n_13705),
.Y(n_14430)
);

INVx2_ASAP7_75t_L g14431 ( 
.A(n_13705),
.Y(n_14431)
);

INVx1_ASAP7_75t_L g14432 ( 
.A(n_13674),
.Y(n_14432)
);

INVx2_ASAP7_75t_L g14433 ( 
.A(n_13705),
.Y(n_14433)
);

INVxp67_ASAP7_75t_SL g14434 ( 
.A(n_13409),
.Y(n_14434)
);

NAND2xp5_ASAP7_75t_L g14435 ( 
.A(n_13358),
.B(n_12910),
.Y(n_14435)
);

INVx5_ASAP7_75t_L g14436 ( 
.A(n_13604),
.Y(n_14436)
);

AND2x4_ASAP7_75t_L g14437 ( 
.A(n_13733),
.B(n_7956),
.Y(n_14437)
);

INVx1_ASAP7_75t_L g14438 ( 
.A(n_13677),
.Y(n_14438)
);

HB1xp67_ASAP7_75t_L g14439 ( 
.A(n_13349),
.Y(n_14439)
);

INVx1_ASAP7_75t_L g14440 ( 
.A(n_13677),
.Y(n_14440)
);

OR2x2_ASAP7_75t_L g14441 ( 
.A(n_13578),
.B(n_11488),
.Y(n_14441)
);

AND2x2_ASAP7_75t_L g14442 ( 
.A(n_13432),
.B(n_7956),
.Y(n_14442)
);

OR2x2_ASAP7_75t_L g14443 ( 
.A(n_13740),
.B(n_11492),
.Y(n_14443)
);

OR2x2_ASAP7_75t_L g14444 ( 
.A(n_14013),
.B(n_11505),
.Y(n_14444)
);

INVx1_ASAP7_75t_L g14445 ( 
.A(n_13678),
.Y(n_14445)
);

INVx1_ASAP7_75t_L g14446 ( 
.A(n_13678),
.Y(n_14446)
);

BUFx3_ASAP7_75t_L g14447 ( 
.A(n_13409),
.Y(n_14447)
);

OR2x2_ASAP7_75t_L g14448 ( 
.A(n_14258),
.B(n_11506),
.Y(n_14448)
);

INVx2_ASAP7_75t_L g14449 ( 
.A(n_13714),
.Y(n_14449)
);

OR2x2_ASAP7_75t_L g14450 ( 
.A(n_14258),
.B(n_11509),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_13683),
.Y(n_14451)
);

NAND4xp25_ASAP7_75t_L g14452 ( 
.A(n_13348),
.B(n_12830),
.C(n_13237),
.D(n_12645),
.Y(n_14452)
);

AND2x2_ASAP7_75t_L g14453 ( 
.A(n_13420),
.B(n_8053),
.Y(n_14453)
);

OR2x2_ASAP7_75t_L g14454 ( 
.A(n_13699),
.B(n_13723),
.Y(n_14454)
);

INVx1_ASAP7_75t_L g14455 ( 
.A(n_13683),
.Y(n_14455)
);

AND2x4_ASAP7_75t_L g14456 ( 
.A(n_13733),
.B(n_8053),
.Y(n_14456)
);

INVx1_ASAP7_75t_L g14457 ( 
.A(n_13765),
.Y(n_14457)
);

INVx2_ASAP7_75t_L g14458 ( 
.A(n_13563),
.Y(n_14458)
);

INVx1_ASAP7_75t_L g14459 ( 
.A(n_13765),
.Y(n_14459)
);

OAI22xp5_ASAP7_75t_L g14460 ( 
.A1(n_13326),
.A2(n_13276),
.B1(n_13281),
.B2(n_12615),
.Y(n_14460)
);

AND2x2_ASAP7_75t_L g14461 ( 
.A(n_13420),
.B(n_8058),
.Y(n_14461)
);

INVx2_ASAP7_75t_L g14462 ( 
.A(n_13563),
.Y(n_14462)
);

AND2x2_ASAP7_75t_L g14463 ( 
.A(n_13449),
.B(n_8058),
.Y(n_14463)
);

AND2x4_ASAP7_75t_L g14464 ( 
.A(n_13449),
.B(n_10011),
.Y(n_14464)
);

HB1xp67_ASAP7_75t_L g14465 ( 
.A(n_13372),
.Y(n_14465)
);

INVx1_ASAP7_75t_L g14466 ( 
.A(n_13767),
.Y(n_14466)
);

INVx2_ASAP7_75t_L g14467 ( 
.A(n_13569),
.Y(n_14467)
);

INVx2_ASAP7_75t_L g14468 ( 
.A(n_13569),
.Y(n_14468)
);

INVx1_ASAP7_75t_L g14469 ( 
.A(n_13767),
.Y(n_14469)
);

NAND2xp5_ASAP7_75t_L g14470 ( 
.A(n_14048),
.B(n_12917),
.Y(n_14470)
);

OAI22xp5_ASAP7_75t_L g14471 ( 
.A1(n_14182),
.A2(n_12622),
.B1(n_13242),
.B2(n_12805),
.Y(n_14471)
);

OR2x6_ASAP7_75t_L g14472 ( 
.A(n_13398),
.B(n_7856),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_13481),
.Y(n_14473)
);

INVx2_ASAP7_75t_R g14474 ( 
.A(n_14264),
.Y(n_14474)
);

HB1xp67_ASAP7_75t_L g14475 ( 
.A(n_13726),
.Y(n_14475)
);

NAND2xp5_ASAP7_75t_L g14476 ( 
.A(n_14147),
.B(n_12925),
.Y(n_14476)
);

BUFx2_ASAP7_75t_L g14477 ( 
.A(n_13520),
.Y(n_14477)
);

INVx1_ASAP7_75t_L g14478 ( 
.A(n_13786),
.Y(n_14478)
);

AND2x2_ASAP7_75t_L g14479 ( 
.A(n_13532),
.B(n_9746),
.Y(n_14479)
);

INVx1_ASAP7_75t_L g14480 ( 
.A(n_13797),
.Y(n_14480)
);

INVx1_ASAP7_75t_L g14481 ( 
.A(n_13331),
.Y(n_14481)
);

AND2x2_ASAP7_75t_L g14482 ( 
.A(n_13523),
.B(n_9746),
.Y(n_14482)
);

INVx1_ASAP7_75t_L g14483 ( 
.A(n_13332),
.Y(n_14483)
);

NAND2xp5_ASAP7_75t_L g14484 ( 
.A(n_13662),
.B(n_12926),
.Y(n_14484)
);

BUFx6f_ASAP7_75t_L g14485 ( 
.A(n_13462),
.Y(n_14485)
);

AND2x2_ASAP7_75t_SL g14486 ( 
.A(n_14272),
.B(n_10015),
.Y(n_14486)
);

NAND2xp5_ASAP7_75t_L g14487 ( 
.A(n_14182),
.B(n_12929),
.Y(n_14487)
);

HB1xp67_ASAP7_75t_L g14488 ( 
.A(n_13938),
.Y(n_14488)
);

BUFx2_ASAP7_75t_L g14489 ( 
.A(n_13787),
.Y(n_14489)
);

INVx1_ASAP7_75t_L g14490 ( 
.A(n_13336),
.Y(n_14490)
);

AND2x2_ASAP7_75t_L g14491 ( 
.A(n_13447),
.B(n_9785),
.Y(n_14491)
);

INVx1_ASAP7_75t_L g14492 ( 
.A(n_13936),
.Y(n_14492)
);

INVx2_ASAP7_75t_L g14493 ( 
.A(n_13579),
.Y(n_14493)
);

AND2x4_ASAP7_75t_L g14494 ( 
.A(n_13361),
.B(n_10015),
.Y(n_14494)
);

BUFx2_ASAP7_75t_L g14495 ( 
.A(n_13325),
.Y(n_14495)
);

INVx2_ASAP7_75t_L g14496 ( 
.A(n_13579),
.Y(n_14496)
);

AND2x2_ASAP7_75t_L g14497 ( 
.A(n_13454),
.B(n_9785),
.Y(n_14497)
);

INVx1_ASAP7_75t_L g14498 ( 
.A(n_13936),
.Y(n_14498)
);

AND2x2_ASAP7_75t_L g14499 ( 
.A(n_13459),
.B(n_9786),
.Y(n_14499)
);

OR2x2_ASAP7_75t_L g14500 ( 
.A(n_13784),
.B(n_11516),
.Y(n_14500)
);

AOI22xp33_ASAP7_75t_L g14501 ( 
.A1(n_13816),
.A2(n_12498),
.B1(n_13026),
.B2(n_13108),
.Y(n_14501)
);

INVx4_ASAP7_75t_SL g14502 ( 
.A(n_13604),
.Y(n_14502)
);

AOI22xp33_ASAP7_75t_L g14503 ( 
.A1(n_14254),
.A2(n_12459),
.B1(n_12907),
.B2(n_12905),
.Y(n_14503)
);

INVx2_ASAP7_75t_L g14504 ( 
.A(n_13628),
.Y(n_14504)
);

INVx1_ASAP7_75t_L g14505 ( 
.A(n_13946),
.Y(n_14505)
);

AO22x1_ASAP7_75t_L g14506 ( 
.A1(n_13805),
.A2(n_7570),
.B1(n_7536),
.B2(n_10015),
.Y(n_14506)
);

AND2x2_ASAP7_75t_L g14507 ( 
.A(n_13392),
.B(n_9786),
.Y(n_14507)
);

OR2x2_ASAP7_75t_L g14508 ( 
.A(n_13448),
.B(n_11518),
.Y(n_14508)
);

NOR2xp33_ASAP7_75t_L g14509 ( 
.A(n_13462),
.B(n_7856),
.Y(n_14509)
);

INVx3_ASAP7_75t_L g14510 ( 
.A(n_13462),
.Y(n_14510)
);

INVx1_ASAP7_75t_L g14511 ( 
.A(n_13946),
.Y(n_14511)
);

BUFx3_ASAP7_75t_L g14512 ( 
.A(n_13465),
.Y(n_14512)
);

NAND2xp5_ASAP7_75t_L g14513 ( 
.A(n_13650),
.B(n_12931),
.Y(n_14513)
);

INVx1_ASAP7_75t_L g14514 ( 
.A(n_13948),
.Y(n_14514)
);

AOI22xp33_ASAP7_75t_L g14515 ( 
.A1(n_14132),
.A2(n_12589),
.B1(n_13298),
.B2(n_13300),
.Y(n_14515)
);

NAND2xp5_ASAP7_75t_L g14516 ( 
.A(n_13422),
.B(n_12943),
.Y(n_14516)
);

INVx1_ASAP7_75t_L g14517 ( 
.A(n_13948),
.Y(n_14517)
);

AND2x2_ASAP7_75t_L g14518 ( 
.A(n_13577),
.B(n_13654),
.Y(n_14518)
);

INVx2_ASAP7_75t_L g14519 ( 
.A(n_13628),
.Y(n_14519)
);

NAND2xp5_ASAP7_75t_L g14520 ( 
.A(n_13494),
.B(n_12948),
.Y(n_14520)
);

AND2x2_ASAP7_75t_L g14521 ( 
.A(n_13438),
.B(n_9832),
.Y(n_14521)
);

OR2x2_ASAP7_75t_L g14522 ( 
.A(n_14236),
.B(n_13317),
.Y(n_14522)
);

AND2x2_ASAP7_75t_L g14523 ( 
.A(n_13455),
.B(n_9832),
.Y(n_14523)
);

NAND2xp5_ASAP7_75t_L g14524 ( 
.A(n_13500),
.B(n_12966),
.Y(n_14524)
);

INVx2_ASAP7_75t_L g14525 ( 
.A(n_13993),
.Y(n_14525)
);

NAND2xp5_ASAP7_75t_L g14526 ( 
.A(n_14181),
.B(n_12970),
.Y(n_14526)
);

INVx1_ASAP7_75t_L g14527 ( 
.A(n_13565),
.Y(n_14527)
);

INVx1_ASAP7_75t_L g14528 ( 
.A(n_13565),
.Y(n_14528)
);

NAND2xp5_ASAP7_75t_L g14529 ( 
.A(n_13554),
.B(n_12973),
.Y(n_14529)
);

HB1xp67_ASAP7_75t_L g14530 ( 
.A(n_13961),
.Y(n_14530)
);

INVx2_ASAP7_75t_L g14531 ( 
.A(n_13993),
.Y(n_14531)
);

AND2x4_ASAP7_75t_L g14532 ( 
.A(n_13361),
.B(n_10015),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_13779),
.Y(n_14533)
);

INVx2_ASAP7_75t_L g14534 ( 
.A(n_13993),
.Y(n_14534)
);

INVx2_ASAP7_75t_L g14535 ( 
.A(n_13838),
.Y(n_14535)
);

BUFx3_ASAP7_75t_L g14536 ( 
.A(n_13465),
.Y(n_14536)
);

INVx1_ASAP7_75t_L g14537 ( 
.A(n_13780),
.Y(n_14537)
);

OR2x2_ASAP7_75t_L g14538 ( 
.A(n_13679),
.B(n_14050),
.Y(n_14538)
);

NAND2xp5_ASAP7_75t_L g14539 ( 
.A(n_14264),
.B(n_12975),
.Y(n_14539)
);

NAND2xp5_ASAP7_75t_L g14540 ( 
.A(n_14265),
.B(n_12983),
.Y(n_14540)
);

NAND2xp5_ASAP7_75t_L g14541 ( 
.A(n_14265),
.B(n_12992),
.Y(n_14541)
);

NAND2xp5_ASAP7_75t_L g14542 ( 
.A(n_13347),
.B(n_13004),
.Y(n_14542)
);

OR2x2_ASAP7_75t_L g14543 ( 
.A(n_14054),
.B(n_11526),
.Y(n_14543)
);

OR2x6_ASAP7_75t_L g14544 ( 
.A(n_13411),
.B(n_7999),
.Y(n_14544)
);

INVx1_ASAP7_75t_L g14545 ( 
.A(n_13782),
.Y(n_14545)
);

INVx1_ASAP7_75t_L g14546 ( 
.A(n_13776),
.Y(n_14546)
);

OR2x2_ASAP7_75t_L g14547 ( 
.A(n_13892),
.B(n_11529),
.Y(n_14547)
);

INVx1_ASAP7_75t_L g14548 ( 
.A(n_13401),
.Y(n_14548)
);

HB1xp67_ASAP7_75t_L g14549 ( 
.A(n_14011),
.Y(n_14549)
);

OR2x2_ASAP7_75t_L g14550 ( 
.A(n_13764),
.B(n_11530),
.Y(n_14550)
);

NAND2xp5_ASAP7_75t_L g14551 ( 
.A(n_13354),
.B(n_8419),
.Y(n_14551)
);

BUFx3_ASAP7_75t_L g14552 ( 
.A(n_13465),
.Y(n_14552)
);

NAND2xp5_ASAP7_75t_L g14553 ( 
.A(n_13690),
.B(n_8419),
.Y(n_14553)
);

AND2x2_ASAP7_75t_L g14554 ( 
.A(n_13464),
.B(n_7536),
.Y(n_14554)
);

BUFx2_ASAP7_75t_L g14555 ( 
.A(n_13325),
.Y(n_14555)
);

AND2x2_ASAP7_75t_L g14556 ( 
.A(n_13555),
.B(n_8883),
.Y(n_14556)
);

NOR2xp33_ASAP7_75t_L g14557 ( 
.A(n_13807),
.B(n_7999),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_13401),
.Y(n_14558)
);

AND2x2_ASAP7_75t_L g14559 ( 
.A(n_13373),
.B(n_8345),
.Y(n_14559)
);

NAND2xp5_ASAP7_75t_L g14560 ( 
.A(n_13691),
.B(n_8419),
.Y(n_14560)
);

HB1xp67_ASAP7_75t_L g14561 ( 
.A(n_13487),
.Y(n_14561)
);

AND2x2_ASAP7_75t_L g14562 ( 
.A(n_13365),
.B(n_8345),
.Y(n_14562)
);

NAND4xp25_ASAP7_75t_L g14563 ( 
.A(n_14020),
.B(n_12500),
.C(n_12976),
.D(n_12856),
.Y(n_14563)
);

AND2x2_ASAP7_75t_L g14564 ( 
.A(n_13370),
.B(n_8345),
.Y(n_14564)
);

AND2x4_ASAP7_75t_L g14565 ( 
.A(n_13381),
.B(n_10023),
.Y(n_14565)
);

NAND2xp5_ASAP7_75t_L g14566 ( 
.A(n_13692),
.B(n_8419),
.Y(n_14566)
);

INVx1_ASAP7_75t_L g14567 ( 
.A(n_13405),
.Y(n_14567)
);

NAND2xp5_ASAP7_75t_L g14568 ( 
.A(n_13697),
.B(n_8419),
.Y(n_14568)
);

INVx2_ASAP7_75t_L g14569 ( 
.A(n_13860),
.Y(n_14569)
);

INVx1_ASAP7_75t_L g14570 ( 
.A(n_13405),
.Y(n_14570)
);

HB1xp67_ASAP7_75t_L g14571 ( 
.A(n_13482),
.Y(n_14571)
);

OR2x2_ASAP7_75t_L g14572 ( 
.A(n_13833),
.B(n_11533),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_13406),
.Y(n_14573)
);

AND2x2_ASAP7_75t_L g14574 ( 
.A(n_13484),
.B(n_8382),
.Y(n_14574)
);

NOR2x1_ASAP7_75t_L g14575 ( 
.A(n_14067),
.B(n_12741),
.Y(n_14575)
);

INVx2_ASAP7_75t_L g14576 ( 
.A(n_13879),
.Y(n_14576)
);

INVx2_ASAP7_75t_L g14577 ( 
.A(n_13378),
.Y(n_14577)
);

AND2x2_ASAP7_75t_L g14578 ( 
.A(n_13519),
.B(n_8382),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_13406),
.Y(n_14579)
);

INVx2_ASAP7_75t_L g14580 ( 
.A(n_13371),
.Y(n_14580)
);

AND2x4_ASAP7_75t_L g14581 ( 
.A(n_13452),
.B(n_13483),
.Y(n_14581)
);

NAND2xp5_ASAP7_75t_L g14582 ( 
.A(n_13702),
.B(n_8419),
.Y(n_14582)
);

AND2x2_ASAP7_75t_L g14583 ( 
.A(n_13661),
.B(n_8382),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_13594),
.B(n_8427),
.Y(n_14584)
);

HB1xp67_ASAP7_75t_L g14585 ( 
.A(n_13482),
.Y(n_14585)
);

OR2x2_ASAP7_75t_L g14586 ( 
.A(n_14045),
.B(n_11536),
.Y(n_14586)
);

INVx3_ASAP7_75t_L g14587 ( 
.A(n_13382),
.Y(n_14587)
);

AND2x2_ASAP7_75t_L g14588 ( 
.A(n_13595),
.B(n_8427),
.Y(n_14588)
);

NOR2x1_ASAP7_75t_L g14589 ( 
.A(n_13809),
.B(n_13017),
.Y(n_14589)
);

OR2x2_ASAP7_75t_L g14590 ( 
.A(n_13954),
.B(n_11537),
.Y(n_14590)
);

INVxp67_ASAP7_75t_SL g14591 ( 
.A(n_13512),
.Y(n_14591)
);

AOI21xp33_ASAP7_75t_L g14592 ( 
.A1(n_13920),
.A2(n_13032),
.B(n_12899),
.Y(n_14592)
);

INVx2_ASAP7_75t_L g14593 ( 
.A(n_13473),
.Y(n_14593)
);

AND2x2_ASAP7_75t_L g14594 ( 
.A(n_13562),
.B(n_8427),
.Y(n_14594)
);

AND2x2_ASAP7_75t_L g14595 ( 
.A(n_13400),
.B(n_8317),
.Y(n_14595)
);

AND2x2_ASAP7_75t_L g14596 ( 
.A(n_13582),
.B(n_8317),
.Y(n_14596)
);

OR2x2_ASAP7_75t_L g14597 ( 
.A(n_13667),
.B(n_11538),
.Y(n_14597)
);

AOI22xp33_ASAP7_75t_L g14598 ( 
.A1(n_14132),
.A2(n_12898),
.B1(n_13110),
.B2(n_12548),
.Y(n_14598)
);

INVxp67_ASAP7_75t_SL g14599 ( 
.A(n_13499),
.Y(n_14599)
);

AND2x2_ASAP7_75t_L g14600 ( 
.A(n_13610),
.B(n_8317),
.Y(n_14600)
);

BUFx2_ASAP7_75t_L g14601 ( 
.A(n_13701),
.Y(n_14601)
);

AND2x2_ASAP7_75t_L g14602 ( 
.A(n_13610),
.B(n_8317),
.Y(n_14602)
);

AND2x2_ASAP7_75t_L g14603 ( 
.A(n_13631),
.B(n_8317),
.Y(n_14603)
);

INVx2_ASAP7_75t_L g14604 ( 
.A(n_13474),
.Y(n_14604)
);

AND2x2_ASAP7_75t_L g14605 ( 
.A(n_13631),
.B(n_8381),
.Y(n_14605)
);

AND2x4_ASAP7_75t_L g14606 ( 
.A(n_13366),
.B(n_10023),
.Y(n_14606)
);

AND2x2_ASAP7_75t_L g14607 ( 
.A(n_13675),
.B(n_13338),
.Y(n_14607)
);

OAI21xp5_ASAP7_75t_L g14608 ( 
.A1(n_13461),
.A2(n_12994),
.B(n_11741),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_13407),
.Y(n_14609)
);

INVx3_ASAP7_75t_L g14610 ( 
.A(n_13611),
.Y(n_14610)
);

INVx1_ASAP7_75t_L g14611 ( 
.A(n_13407),
.Y(n_14611)
);

AOI22xp33_ASAP7_75t_L g14612 ( 
.A1(n_14137),
.A2(n_12551),
.B1(n_12553),
.B2(n_13301),
.Y(n_14612)
);

NOR2x1p5_ASAP7_75t_L g14613 ( 
.A(n_13623),
.B(n_10434),
.Y(n_14613)
);

INVx1_ASAP7_75t_L g14614 ( 
.A(n_13436),
.Y(n_14614)
);

BUFx2_ASAP7_75t_L g14615 ( 
.A(n_13701),
.Y(n_14615)
);

NOR2xp33_ASAP7_75t_L g14616 ( 
.A(n_13568),
.B(n_7999),
.Y(n_14616)
);

NAND2xp5_ASAP7_75t_L g14617 ( 
.A(n_13708),
.B(n_8419),
.Y(n_14617)
);

INVx2_ASAP7_75t_L g14618 ( 
.A(n_13475),
.Y(n_14618)
);

HB1xp67_ASAP7_75t_L g14619 ( 
.A(n_13482),
.Y(n_14619)
);

NAND2xp5_ASAP7_75t_L g14620 ( 
.A(n_13713),
.B(n_11540),
.Y(n_14620)
);

AND2x4_ASAP7_75t_L g14621 ( 
.A(n_13366),
.B(n_10023),
.Y(n_14621)
);

AND2x2_ASAP7_75t_L g14622 ( 
.A(n_13675),
.B(n_8381),
.Y(n_14622)
);

AOI22xp33_ASAP7_75t_L g14623 ( 
.A1(n_14137),
.A2(n_13090),
.B1(n_12685),
.B2(n_12946),
.Y(n_14623)
);

INVx2_ASAP7_75t_L g14624 ( 
.A(n_13781),
.Y(n_14624)
);

AND2x2_ASAP7_75t_L g14625 ( 
.A(n_13338),
.B(n_13868),
.Y(n_14625)
);

BUFx2_ASAP7_75t_L g14626 ( 
.A(n_13446),
.Y(n_14626)
);

INVx2_ASAP7_75t_L g14627 ( 
.A(n_13781),
.Y(n_14627)
);

NOR2xp33_ASAP7_75t_L g14628 ( 
.A(n_13568),
.B(n_7999),
.Y(n_14628)
);

HB1xp67_ASAP7_75t_L g14629 ( 
.A(n_13485),
.Y(n_14629)
);

AND2x2_ASAP7_75t_L g14630 ( 
.A(n_13882),
.B(n_8381),
.Y(n_14630)
);

INVx1_ASAP7_75t_L g14631 ( 
.A(n_13495),
.Y(n_14631)
);

OAI21xp5_ASAP7_75t_SL g14632 ( 
.A1(n_13424),
.A2(n_12891),
.B(n_12816),
.Y(n_14632)
);

INVx1_ASAP7_75t_L g14633 ( 
.A(n_14006),
.Y(n_14633)
);

OR2x2_ASAP7_75t_L g14634 ( 
.A(n_13770),
.B(n_11547),
.Y(n_14634)
);

BUFx2_ASAP7_75t_SL g14635 ( 
.A(n_13591),
.Y(n_14635)
);

INVx1_ASAP7_75t_L g14636 ( 
.A(n_14017),
.Y(n_14636)
);

INVx1_ASAP7_75t_L g14637 ( 
.A(n_14028),
.Y(n_14637)
);

INVx1_ASAP7_75t_L g14638 ( 
.A(n_14033),
.Y(n_14638)
);

INVxp67_ASAP7_75t_SL g14639 ( 
.A(n_13571),
.Y(n_14639)
);

AOI22xp33_ASAP7_75t_L g14640 ( 
.A1(n_14294),
.A2(n_12990),
.B1(n_13005),
.B2(n_12936),
.Y(n_14640)
);

HB1xp67_ASAP7_75t_L g14641 ( 
.A(n_13743),
.Y(n_14641)
);

INVx2_ASAP7_75t_L g14642 ( 
.A(n_13796),
.Y(n_14642)
);

AND2x2_ASAP7_75t_L g14643 ( 
.A(n_13561),
.B(n_8381),
.Y(n_14643)
);

AOI22xp33_ASAP7_75t_L g14644 ( 
.A1(n_14293),
.A2(n_12942),
.B1(n_12924),
.B2(n_13064),
.Y(n_14644)
);

NAND3xp33_ASAP7_75t_L g14645 ( 
.A(n_13997),
.B(n_13920),
.C(n_14267),
.Y(n_14645)
);

BUFx2_ASAP7_75t_L g14646 ( 
.A(n_13446),
.Y(n_14646)
);

INVx2_ASAP7_75t_L g14647 ( 
.A(n_13796),
.Y(n_14647)
);

AND2x2_ASAP7_75t_L g14648 ( 
.A(n_13583),
.B(n_8381),
.Y(n_14648)
);

HB1xp67_ASAP7_75t_L g14649 ( 
.A(n_13750),
.Y(n_14649)
);

INVx1_ASAP7_75t_L g14650 ( 
.A(n_14036),
.Y(n_14650)
);

INVx1_ASAP7_75t_L g14651 ( 
.A(n_13584),
.Y(n_14651)
);

OR2x2_ASAP7_75t_L g14652 ( 
.A(n_14093),
.B(n_11552),
.Y(n_14652)
);

AND2x2_ASAP7_75t_L g14653 ( 
.A(n_13586),
.B(n_8381),
.Y(n_14653)
);

OAI22xp5_ASAP7_75t_L g14654 ( 
.A1(n_14194),
.A2(n_12556),
.B1(n_12505),
.B2(n_12949),
.Y(n_14654)
);

AND2x4_ASAP7_75t_SL g14655 ( 
.A(n_13576),
.B(n_7908),
.Y(n_14655)
);

INVx2_ASAP7_75t_L g14656 ( 
.A(n_13832),
.Y(n_14656)
);

OR2x2_ASAP7_75t_L g14657 ( 
.A(n_13660),
.B(n_11553),
.Y(n_14657)
);

INVx1_ASAP7_75t_L g14658 ( 
.A(n_13585),
.Y(n_14658)
);

INVx2_ASAP7_75t_L g14659 ( 
.A(n_13832),
.Y(n_14659)
);

INVx1_ASAP7_75t_L g14660 ( 
.A(n_13587),
.Y(n_14660)
);

AND2x4_ASAP7_75t_L g14661 ( 
.A(n_13434),
.B(n_10023),
.Y(n_14661)
);

INVx1_ASAP7_75t_L g14662 ( 
.A(n_13588),
.Y(n_14662)
);

AOI22xp33_ASAP7_75t_L g14663 ( 
.A1(n_14165),
.A2(n_13106),
.B1(n_13075),
.B2(n_12824),
.Y(n_14663)
);

AND2x2_ASAP7_75t_L g14664 ( 
.A(n_13673),
.B(n_8385),
.Y(n_14664)
);

NAND2xp5_ASAP7_75t_L g14665 ( 
.A(n_13720),
.B(n_13724),
.Y(n_14665)
);

AND2x2_ASAP7_75t_L g14666 ( 
.A(n_13688),
.B(n_8385),
.Y(n_14666)
);

INVx2_ASAP7_75t_L g14667 ( 
.A(n_13837),
.Y(n_14667)
);

NAND2xp5_ASAP7_75t_L g14668 ( 
.A(n_13727),
.B(n_11557),
.Y(n_14668)
);

INVx1_ASAP7_75t_L g14669 ( 
.A(n_13593),
.Y(n_14669)
);

AND2x4_ASAP7_75t_SL g14670 ( 
.A(n_13604),
.B(n_13387),
.Y(n_14670)
);

INVx1_ASAP7_75t_L g14671 ( 
.A(n_13596),
.Y(n_14671)
);

INVx3_ASAP7_75t_L g14672 ( 
.A(n_13470),
.Y(n_14672)
);

INVx2_ASAP7_75t_L g14673 ( 
.A(n_13837),
.Y(n_14673)
);

INVx4_ASAP7_75t_L g14674 ( 
.A(n_13591),
.Y(n_14674)
);

NAND2xp5_ASAP7_75t_L g14675 ( 
.A(n_13728),
.B(n_11560),
.Y(n_14675)
);

INVx1_ASAP7_75t_L g14676 ( 
.A(n_13600),
.Y(n_14676)
);

INVx1_ASAP7_75t_L g14677 ( 
.A(n_13609),
.Y(n_14677)
);

AND2x2_ASAP7_75t_L g14678 ( 
.A(n_13694),
.B(n_8385),
.Y(n_14678)
);

NAND2xp5_ASAP7_75t_L g14679 ( 
.A(n_13356),
.B(n_11564),
.Y(n_14679)
);

INVx1_ASAP7_75t_L g14680 ( 
.A(n_13612),
.Y(n_14680)
);

AND2x2_ASAP7_75t_L g14681 ( 
.A(n_13769),
.B(n_8385),
.Y(n_14681)
);

AND2x2_ASAP7_75t_L g14682 ( 
.A(n_13659),
.B(n_8385),
.Y(n_14682)
);

INVx1_ASAP7_75t_L g14683 ( 
.A(n_13613),
.Y(n_14683)
);

HB1xp67_ASAP7_75t_L g14684 ( 
.A(n_13752),
.Y(n_14684)
);

BUFx2_ASAP7_75t_L g14685 ( 
.A(n_14267),
.Y(n_14685)
);

INVx1_ASAP7_75t_L g14686 ( 
.A(n_13621),
.Y(n_14686)
);

AND2x2_ASAP7_75t_L g14687 ( 
.A(n_13506),
.B(n_8385),
.Y(n_14687)
);

INVx1_ASAP7_75t_L g14688 ( 
.A(n_13629),
.Y(n_14688)
);

INVx1_ASAP7_75t_L g14689 ( 
.A(n_13639),
.Y(n_14689)
);

AND2x2_ASAP7_75t_L g14690 ( 
.A(n_13508),
.B(n_8394),
.Y(n_14690)
);

INVxp67_ASAP7_75t_SL g14691 ( 
.A(n_13360),
.Y(n_14691)
);

INVx1_ASAP7_75t_L g14692 ( 
.A(n_13640),
.Y(n_14692)
);

INVxp67_ASAP7_75t_L g14693 ( 
.A(n_13393),
.Y(n_14693)
);

OR2x2_ASAP7_75t_L g14694 ( 
.A(n_13635),
.B(n_11567),
.Y(n_14694)
);

NAND2x1p5_ASAP7_75t_SL g14695 ( 
.A(n_13872),
.B(n_7859),
.Y(n_14695)
);

INVxp67_ASAP7_75t_L g14696 ( 
.A(n_13412),
.Y(n_14696)
);

INVx1_ASAP7_75t_L g14697 ( 
.A(n_13641),
.Y(n_14697)
);

INVx2_ASAP7_75t_L g14698 ( 
.A(n_14086),
.Y(n_14698)
);

HB1xp67_ASAP7_75t_L g14699 ( 
.A(n_13756),
.Y(n_14699)
);

NAND2xp5_ASAP7_75t_L g14700 ( 
.A(n_13757),
.B(n_11568),
.Y(n_14700)
);

NAND2xp5_ASAP7_75t_SL g14701 ( 
.A(n_14176),
.B(n_12952),
.Y(n_14701)
);

AND2x4_ASAP7_75t_L g14702 ( 
.A(n_13434),
.B(n_10054),
.Y(n_14702)
);

NAND2xp5_ASAP7_75t_L g14703 ( 
.A(n_13761),
.B(n_11572),
.Y(n_14703)
);

AND2x4_ASAP7_75t_L g14704 ( 
.A(n_13444),
.B(n_10054),
.Y(n_14704)
);

NAND2xp5_ASAP7_75t_L g14705 ( 
.A(n_13788),
.B(n_11576),
.Y(n_14705)
);

INVx2_ASAP7_75t_L g14706 ( 
.A(n_13396),
.Y(n_14706)
);

AOI22xp33_ASAP7_75t_SL g14707 ( 
.A1(n_14287),
.A2(n_12964),
.B1(n_12011),
.B2(n_12093),
.Y(n_14707)
);

AND2x2_ASAP7_75t_L g14708 ( 
.A(n_13513),
.B(n_8394),
.Y(n_14708)
);

OR2x2_ASAP7_75t_L g14709 ( 
.A(n_13402),
.B(n_11581),
.Y(n_14709)
);

AND2x4_ASAP7_75t_L g14710 ( 
.A(n_13444),
.B(n_10054),
.Y(n_14710)
);

INVx1_ASAP7_75t_L g14711 ( 
.A(n_13689),
.Y(n_14711)
);

INVx1_ASAP7_75t_L g14712 ( 
.A(n_13696),
.Y(n_14712)
);

AND2x2_ASAP7_75t_L g14713 ( 
.A(n_13636),
.B(n_8394),
.Y(n_14713)
);

INVx1_ASAP7_75t_L g14714 ( 
.A(n_13700),
.Y(n_14714)
);

INVx1_ASAP7_75t_L g14715 ( 
.A(n_13706),
.Y(n_14715)
);

INVx1_ASAP7_75t_L g14716 ( 
.A(n_13711),
.Y(n_14716)
);

INVxp67_ASAP7_75t_L g14717 ( 
.A(n_13754),
.Y(n_14717)
);

AND2x4_ASAP7_75t_L g14718 ( 
.A(n_13900),
.B(n_10054),
.Y(n_14718)
);

INVx1_ASAP7_75t_L g14719 ( 
.A(n_13715),
.Y(n_14719)
);

AND2x2_ASAP7_75t_L g14720 ( 
.A(n_13590),
.B(n_8394),
.Y(n_14720)
);

NAND2xp5_ASAP7_75t_L g14721 ( 
.A(n_13793),
.B(n_13802),
.Y(n_14721)
);

OR2x2_ASAP7_75t_L g14722 ( 
.A(n_13319),
.B(n_11584),
.Y(n_14722)
);

INVx1_ASAP7_75t_L g14723 ( 
.A(n_13717),
.Y(n_14723)
);

AOI22xp33_ASAP7_75t_SL g14724 ( 
.A1(n_14285),
.A2(n_12093),
.B1(n_11521),
.B2(n_11450),
.Y(n_14724)
);

NAND2xp5_ASAP7_75t_L g14725 ( 
.A(n_13850),
.B(n_11585),
.Y(n_14725)
);

NAND2xp5_ASAP7_75t_L g14726 ( 
.A(n_14209),
.B(n_11588),
.Y(n_14726)
);

AND2x4_ASAP7_75t_L g14727 ( 
.A(n_13905),
.B(n_13906),
.Y(n_14727)
);

INVx1_ASAP7_75t_L g14728 ( 
.A(n_13719),
.Y(n_14728)
);

AND2x2_ASAP7_75t_L g14729 ( 
.A(n_13544),
.B(n_8394),
.Y(n_14729)
);

INVx1_ASAP7_75t_L g14730 ( 
.A(n_13721),
.Y(n_14730)
);

INVx1_ASAP7_75t_L g14731 ( 
.A(n_13725),
.Y(n_14731)
);

NAND2xp5_ASAP7_75t_L g14732 ( 
.A(n_14210),
.B(n_11595),
.Y(n_14732)
);

AND2x4_ASAP7_75t_L g14733 ( 
.A(n_13897),
.B(n_8394),
.Y(n_14733)
);

INVx2_ASAP7_75t_SL g14734 ( 
.A(n_13591),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_13730),
.Y(n_14735)
);

INVx2_ASAP7_75t_L g14736 ( 
.A(n_13397),
.Y(n_14736)
);

INVx2_ASAP7_75t_L g14737 ( 
.A(n_13403),
.Y(n_14737)
);

INVxp67_ASAP7_75t_SL g14738 ( 
.A(n_13362),
.Y(n_14738)
);

INVx2_ASAP7_75t_L g14739 ( 
.A(n_13404),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_13738),
.Y(n_14740)
);

AND2x2_ASAP7_75t_L g14741 ( 
.A(n_13847),
.B(n_13849),
.Y(n_14741)
);

AND2x2_ASAP7_75t_L g14742 ( 
.A(n_13375),
.B(n_8403),
.Y(n_14742)
);

AND2x2_ASAP7_75t_L g14743 ( 
.A(n_13541),
.B(n_8403),
.Y(n_14743)
);

AND2x2_ASAP7_75t_L g14744 ( 
.A(n_13542),
.B(n_8403),
.Y(n_14744)
);

OAI222xp33_ASAP7_75t_L g14745 ( 
.A1(n_13376),
.A2(n_12812),
.B1(n_12957),
.B2(n_13030),
.C1(n_11074),
.C2(n_11061),
.Y(n_14745)
);

HB1xp67_ASAP7_75t_L g14746 ( 
.A(n_13408),
.Y(n_14746)
);

INVx1_ASAP7_75t_L g14747 ( 
.A(n_13742),
.Y(n_14747)
);

OR2x2_ASAP7_75t_L g14748 ( 
.A(n_13321),
.B(n_13369),
.Y(n_14748)
);

AOI22xp5_ASAP7_75t_L g14749 ( 
.A1(n_14167),
.A2(n_12555),
.B1(n_12843),
.B2(n_12837),
.Y(n_14749)
);

OR2x2_ASAP7_75t_L g14750 ( 
.A(n_13603),
.B(n_11596),
.Y(n_14750)
);

INVx2_ASAP7_75t_L g14751 ( 
.A(n_13413),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_13744),
.Y(n_14752)
);

INVx1_ASAP7_75t_L g14753 ( 
.A(n_13745),
.Y(n_14753)
);

INVx2_ASAP7_75t_L g14754 ( 
.A(n_13768),
.Y(n_14754)
);

INVx1_ASAP7_75t_L g14755 ( 
.A(n_13753),
.Y(n_14755)
);

INVx1_ASAP7_75t_L g14756 ( 
.A(n_13760),
.Y(n_14756)
);

AND2x2_ASAP7_75t_SL g14757 ( 
.A(n_13918),
.B(n_9578),
.Y(n_14757)
);

INVx1_ASAP7_75t_L g14758 ( 
.A(n_13774),
.Y(n_14758)
);

INVx2_ASAP7_75t_SL g14759 ( 
.A(n_13592),
.Y(n_14759)
);

AND2x2_ASAP7_75t_L g14760 ( 
.A(n_13419),
.B(n_8403),
.Y(n_14760)
);

INVx1_ASAP7_75t_L g14761 ( 
.A(n_13414),
.Y(n_14761)
);

NAND2xp5_ASAP7_75t_L g14762 ( 
.A(n_14193),
.B(n_11600),
.Y(n_14762)
);

INVx2_ASAP7_75t_L g14763 ( 
.A(n_13790),
.Y(n_14763)
);

INVx2_ASAP7_75t_L g14764 ( 
.A(n_13791),
.Y(n_14764)
);

OR2x2_ASAP7_75t_L g14765 ( 
.A(n_14105),
.B(n_11601),
.Y(n_14765)
);

BUFx3_ASAP7_75t_L g14766 ( 
.A(n_13417),
.Y(n_14766)
);

INVx3_ASAP7_75t_L g14767 ( 
.A(n_13470),
.Y(n_14767)
);

AND2x2_ASAP7_75t_L g14768 ( 
.A(n_13773),
.B(n_8403),
.Y(n_14768)
);

NAND2xp5_ASAP7_75t_L g14769 ( 
.A(n_13826),
.B(n_11602),
.Y(n_14769)
);

NAND2xp5_ASAP7_75t_L g14770 ( 
.A(n_13976),
.B(n_11603),
.Y(n_14770)
);

AND2x4_ASAP7_75t_L g14771 ( 
.A(n_13747),
.B(n_8403),
.Y(n_14771)
);

OR2x2_ASAP7_75t_L g14772 ( 
.A(n_13478),
.B(n_11607),
.Y(n_14772)
);

INVxp67_ASAP7_75t_SL g14773 ( 
.A(n_13377),
.Y(n_14773)
);

INVx1_ASAP7_75t_SL g14774 ( 
.A(n_13884),
.Y(n_14774)
);

NOR2xp33_ASAP7_75t_L g14775 ( 
.A(n_13592),
.B(n_8004),
.Y(n_14775)
);

INVx6_ASAP7_75t_L g14776 ( 
.A(n_13592),
.Y(n_14776)
);

INVxp67_ASAP7_75t_L g14777 ( 
.A(n_13809),
.Y(n_14777)
);

INVx1_ASAP7_75t_L g14778 ( 
.A(n_13418),
.Y(n_14778)
);

INVxp67_ASAP7_75t_L g14779 ( 
.A(n_14226),
.Y(n_14779)
);

AND2x2_ASAP7_75t_L g14780 ( 
.A(n_13853),
.B(n_8435),
.Y(n_14780)
);

INVxp67_ASAP7_75t_SL g14781 ( 
.A(n_14018),
.Y(n_14781)
);

INVx1_ASAP7_75t_L g14782 ( 
.A(n_13427),
.Y(n_14782)
);

AOI22xp33_ASAP7_75t_L g14783 ( 
.A1(n_14172),
.A2(n_14207),
.B1(n_14278),
.B2(n_14164),
.Y(n_14783)
);

INVx2_ASAP7_75t_L g14784 ( 
.A(n_13798),
.Y(n_14784)
);

INVxp67_ASAP7_75t_SL g14785 ( 
.A(n_13343),
.Y(n_14785)
);

INVx1_ASAP7_75t_L g14786 ( 
.A(n_13430),
.Y(n_14786)
);

AND2x2_ASAP7_75t_L g14787 ( 
.A(n_13855),
.B(n_8435),
.Y(n_14787)
);

INVx1_ASAP7_75t_L g14788 ( 
.A(n_13437),
.Y(n_14788)
);

INVx2_ASAP7_75t_L g14789 ( 
.A(n_13799),
.Y(n_14789)
);

NAND2xp5_ASAP7_75t_L g14790 ( 
.A(n_13979),
.B(n_11611),
.Y(n_14790)
);

AND2x2_ASAP7_75t_L g14791 ( 
.A(n_13856),
.B(n_8435),
.Y(n_14791)
);

HB1xp67_ASAP7_75t_L g14792 ( 
.A(n_13351),
.Y(n_14792)
);

INVx1_ASAP7_75t_L g14793 ( 
.A(n_13450),
.Y(n_14793)
);

INVx1_ASAP7_75t_L g14794 ( 
.A(n_13460),
.Y(n_14794)
);

NAND2xp5_ASAP7_75t_L g14795 ( 
.A(n_14154),
.B(n_11618),
.Y(n_14795)
);

OR2x2_ASAP7_75t_L g14796 ( 
.A(n_13529),
.B(n_11620),
.Y(n_14796)
);

INVx1_ASAP7_75t_L g14797 ( 
.A(n_13463),
.Y(n_14797)
);

AND2x2_ASAP7_75t_L g14798 ( 
.A(n_13533),
.B(n_8435),
.Y(n_14798)
);

AND2x2_ASAP7_75t_L g14799 ( 
.A(n_13534),
.B(n_13666),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_13476),
.Y(n_14800)
);

AND2x2_ASAP7_75t_L g14801 ( 
.A(n_13670),
.B(n_8435),
.Y(n_14801)
);

BUFx2_ASAP7_75t_L g14802 ( 
.A(n_13737),
.Y(n_14802)
);

AND2x4_ASAP7_75t_L g14803 ( 
.A(n_13831),
.B(n_8435),
.Y(n_14803)
);

AND2x2_ASAP7_75t_L g14804 ( 
.A(n_13501),
.B(n_8450),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_13480),
.Y(n_14805)
);

AND2x2_ASAP7_75t_L g14806 ( 
.A(n_13608),
.B(n_13619),
.Y(n_14806)
);

AND2x2_ASAP7_75t_L g14807 ( 
.A(n_13620),
.B(n_8450),
.Y(n_14807)
);

INVx1_ASAP7_75t_L g14808 ( 
.A(n_13486),
.Y(n_14808)
);

AND2x2_ASAP7_75t_L g14809 ( 
.A(n_13626),
.B(n_8450),
.Y(n_14809)
);

INVx2_ASAP7_75t_L g14810 ( 
.A(n_13815),
.Y(n_14810)
);

NAND2xp5_ASAP7_75t_L g14811 ( 
.A(n_13663),
.B(n_11621),
.Y(n_14811)
);

AND2x2_ASAP7_75t_L g14812 ( 
.A(n_13633),
.B(n_8450),
.Y(n_14812)
);

INVx1_ASAP7_75t_L g14813 ( 
.A(n_13489),
.Y(n_14813)
);

INVx2_ASAP7_75t_L g14814 ( 
.A(n_13817),
.Y(n_14814)
);

INVx2_ASAP7_75t_L g14815 ( 
.A(n_14056),
.Y(n_14815)
);

AND2x2_ASAP7_75t_L g14816 ( 
.A(n_13634),
.B(n_8450),
.Y(n_14816)
);

AND2x2_ASAP7_75t_L g14817 ( 
.A(n_13695),
.B(n_8450),
.Y(n_14817)
);

NAND2xp5_ASAP7_75t_L g14818 ( 
.A(n_13664),
.B(n_11622),
.Y(n_14818)
);

INVx1_ASAP7_75t_SL g14819 ( 
.A(n_13894),
.Y(n_14819)
);

INVx1_ASAP7_75t_L g14820 ( 
.A(n_13490),
.Y(n_14820)
);

INVx1_ASAP7_75t_L g14821 ( 
.A(n_13493),
.Y(n_14821)
);

INVx1_ASAP7_75t_SL g14822 ( 
.A(n_13923),
.Y(n_14822)
);

AOI22xp33_ASAP7_75t_L g14823 ( 
.A1(n_14278),
.A2(n_12933),
.B1(n_12963),
.B2(n_12855),
.Y(n_14823)
);

INVx1_ASAP7_75t_L g14824 ( 
.A(n_13497),
.Y(n_14824)
);

AOI22xp5_ASAP7_75t_L g14825 ( 
.A1(n_14266),
.A2(n_13149),
.B1(n_13236),
.B2(n_13138),
.Y(n_14825)
);

NOR2xp33_ASAP7_75t_SL g14826 ( 
.A(n_14100),
.B(n_10486),
.Y(n_14826)
);

BUFx2_ASAP7_75t_L g14827 ( 
.A(n_13737),
.Y(n_14827)
);

HB1xp67_ASAP7_75t_L g14828 ( 
.A(n_13355),
.Y(n_14828)
);

INVx2_ASAP7_75t_L g14829 ( 
.A(n_14056),
.Y(n_14829)
);

NAND2xp5_ASAP7_75t_L g14830 ( 
.A(n_13668),
.B(n_11626),
.Y(n_14830)
);

OR2x2_ASAP7_75t_L g14831 ( 
.A(n_14136),
.B(n_11628),
.Y(n_14831)
);

AOI22xp33_ASAP7_75t_L g14832 ( 
.A1(n_14266),
.A2(n_13293),
.B1(n_13294),
.B2(n_13263),
.Y(n_14832)
);

INVx1_ASAP7_75t_L g14833 ( 
.A(n_13503),
.Y(n_14833)
);

INVx2_ASAP7_75t_L g14834 ( 
.A(n_13548),
.Y(n_14834)
);

OR2x2_ASAP7_75t_L g14835 ( 
.A(n_14139),
.B(n_11631),
.Y(n_14835)
);

BUFx2_ASAP7_75t_L g14836 ( 
.A(n_13488),
.Y(n_14836)
);

AND2x2_ASAP7_75t_L g14837 ( 
.A(n_13440),
.B(n_8004),
.Y(n_14837)
);

AND2x2_ASAP7_75t_L g14838 ( 
.A(n_13917),
.B(n_8004),
.Y(n_14838)
);

AND2x2_ASAP7_75t_L g14839 ( 
.A(n_13827),
.B(n_8004),
.Y(n_14839)
);

INVxp67_ASAP7_75t_SL g14840 ( 
.A(n_13507),
.Y(n_14840)
);

INVx1_ASAP7_75t_SL g14841 ( 
.A(n_13930),
.Y(n_14841)
);

AND2x2_ASAP7_75t_L g14842 ( 
.A(n_13836),
.B(n_8014),
.Y(n_14842)
);

INVx2_ASAP7_75t_L g14843 ( 
.A(n_13558),
.Y(n_14843)
);

INVx1_ASAP7_75t_L g14844 ( 
.A(n_13511),
.Y(n_14844)
);

NAND2x1p5_ASAP7_75t_SL g14845 ( 
.A(n_13968),
.B(n_7859),
.Y(n_14845)
);

AND2x2_ASAP7_75t_L g14846 ( 
.A(n_13535),
.B(n_8014),
.Y(n_14846)
);

OR2x2_ASAP7_75t_L g14847 ( 
.A(n_13441),
.B(n_11633),
.Y(n_14847)
);

AND2x4_ASAP7_75t_L g14848 ( 
.A(n_13652),
.B(n_10303),
.Y(n_14848)
);

BUFx2_ASAP7_75t_L g14849 ( 
.A(n_13488),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_13515),
.Y(n_14850)
);

AND2x2_ASAP7_75t_L g14851 ( 
.A(n_13538),
.B(n_8014),
.Y(n_14851)
);

INVx2_ASAP7_75t_L g14852 ( 
.A(n_13564),
.Y(n_14852)
);

INVxp67_ASAP7_75t_L g14853 ( 
.A(n_13965),
.Y(n_14853)
);

INVx2_ASAP7_75t_L g14854 ( 
.A(n_13567),
.Y(n_14854)
);

INVx2_ASAP7_75t_L g14855 ( 
.A(n_13581),
.Y(n_14855)
);

AND2x2_ASAP7_75t_L g14856 ( 
.A(n_13651),
.B(n_8014),
.Y(n_14856)
);

AND2x2_ASAP7_75t_L g14857 ( 
.A(n_13655),
.B(n_8067),
.Y(n_14857)
);

AND2x2_ASAP7_75t_L g14858 ( 
.A(n_13656),
.B(n_8067),
.Y(n_14858)
);

AND2x2_ASAP7_75t_L g14859 ( 
.A(n_13425),
.B(n_8067),
.Y(n_14859)
);

HB1xp67_ASAP7_75t_L g14860 ( 
.A(n_13828),
.Y(n_14860)
);

INVx2_ASAP7_75t_L g14861 ( 
.A(n_13589),
.Y(n_14861)
);

INVx2_ASAP7_75t_L g14862 ( 
.A(n_13607),
.Y(n_14862)
);

INVx1_ASAP7_75t_L g14863 ( 
.A(n_13516),
.Y(n_14863)
);

AND2x2_ASAP7_75t_L g14864 ( 
.A(n_13431),
.B(n_8067),
.Y(n_14864)
);

INVx1_ASAP7_75t_L g14865 ( 
.A(n_13517),
.Y(n_14865)
);

NAND2xp5_ASAP7_75t_L g14866 ( 
.A(n_13672),
.B(n_11646),
.Y(n_14866)
);

AND2x4_ASAP7_75t_L g14867 ( 
.A(n_13652),
.B(n_10303),
.Y(n_14867)
);

AND2x2_ASAP7_75t_L g14868 ( 
.A(n_13439),
.B(n_8071),
.Y(n_14868)
);

INVx2_ASAP7_75t_L g14869 ( 
.A(n_13615),
.Y(n_14869)
);

AOI22xp33_ASAP7_75t_L g14870 ( 
.A1(n_13808),
.A2(n_11068),
.B1(n_11074),
.B2(n_11059),
.Y(n_14870)
);

INVxp67_ASAP7_75t_SL g14871 ( 
.A(n_13880),
.Y(n_14871)
);

INVx3_ASAP7_75t_L g14872 ( 
.A(n_13505),
.Y(n_14872)
);

AND2x2_ASAP7_75t_L g14873 ( 
.A(n_13642),
.B(n_8071),
.Y(n_14873)
);

AND2x2_ASAP7_75t_L g14874 ( 
.A(n_13645),
.B(n_8071),
.Y(n_14874)
);

OR2x2_ASAP7_75t_L g14875 ( 
.A(n_13681),
.B(n_11647),
.Y(n_14875)
);

INVx2_ASAP7_75t_L g14876 ( 
.A(n_13616),
.Y(n_14876)
);

INVx2_ASAP7_75t_SL g14877 ( 
.A(n_13505),
.Y(n_14877)
);

INVx2_ASAP7_75t_L g14878 ( 
.A(n_13625),
.Y(n_14878)
);

AND2x2_ASAP7_75t_L g14879 ( 
.A(n_13649),
.B(n_8071),
.Y(n_14879)
);

NAND2xp5_ASAP7_75t_L g14880 ( 
.A(n_13687),
.B(n_11657),
.Y(n_14880)
);

INVx2_ASAP7_75t_L g14881 ( 
.A(n_13632),
.Y(n_14881)
);

INVx2_ASAP7_75t_L g14882 ( 
.A(n_13643),
.Y(n_14882)
);

OR2x2_ASAP7_75t_L g14883 ( 
.A(n_13597),
.B(n_11658),
.Y(n_14883)
);

CKINVDCx20_ASAP7_75t_R g14884 ( 
.A(n_14187),
.Y(n_14884)
);

INVx3_ASAP7_75t_L g14885 ( 
.A(n_13926),
.Y(n_14885)
);

AND2x2_ASAP7_75t_L g14886 ( 
.A(n_13559),
.B(n_11662),
.Y(n_14886)
);

NOR2xp33_ASAP7_75t_L g14887 ( 
.A(n_13926),
.B(n_6742),
.Y(n_14887)
);

AND2x2_ASAP7_75t_L g14888 ( 
.A(n_13869),
.B(n_11668),
.Y(n_14888)
);

OR2x2_ASAP7_75t_L g14889 ( 
.A(n_13624),
.B(n_11673),
.Y(n_14889)
);

AND2x2_ASAP7_75t_L g14890 ( 
.A(n_13870),
.B(n_11674),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_13525),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_13527),
.Y(n_14892)
);

INVx1_ASAP7_75t_L g14893 ( 
.A(n_13528),
.Y(n_14893)
);

BUFx3_ASAP7_75t_L g14894 ( 
.A(n_13707),
.Y(n_14894)
);

BUFx2_ASAP7_75t_L g14895 ( 
.A(n_13852),
.Y(n_14895)
);

AND2x2_ASAP7_75t_L g14896 ( 
.A(n_13877),
.B(n_11676),
.Y(n_14896)
);

NAND2xp5_ASAP7_75t_L g14897 ( 
.A(n_14098),
.B(n_11680),
.Y(n_14897)
);

NAND2xp5_ASAP7_75t_L g14898 ( 
.A(n_13902),
.B(n_11685),
.Y(n_14898)
);

AND2x4_ASAP7_75t_SL g14899 ( 
.A(n_13959),
.B(n_7908),
.Y(n_14899)
);

BUFx3_ASAP7_75t_L g14900 ( 
.A(n_14012),
.Y(n_14900)
);

AND2x2_ASAP7_75t_L g14901 ( 
.A(n_13755),
.B(n_11687),
.Y(n_14901)
);

INVx1_ASAP7_75t_L g14902 ( 
.A(n_13531),
.Y(n_14902)
);

INVx2_ASAP7_75t_L g14903 ( 
.A(n_13646),
.Y(n_14903)
);

HB1xp67_ASAP7_75t_L g14904 ( 
.A(n_13421),
.Y(n_14904)
);

INVx2_ASAP7_75t_L g14905 ( 
.A(n_14015),
.Y(n_14905)
);

OAI22xp5_ASAP7_75t_L g14906 ( 
.A1(n_13530),
.A2(n_8376),
.B1(n_10582),
.B2(n_10578),
.Y(n_14906)
);

AND2x2_ASAP7_75t_L g14907 ( 
.A(n_13599),
.B(n_11691),
.Y(n_14907)
);

INVx1_ASAP7_75t_L g14908 ( 
.A(n_13536),
.Y(n_14908)
);

BUFx2_ASAP7_75t_L g14909 ( 
.A(n_13653),
.Y(n_14909)
);

NAND2xp5_ASAP7_75t_SL g14910 ( 
.A(n_14249),
.B(n_13732),
.Y(n_14910)
);

AND2x2_ASAP7_75t_L g14911 ( 
.A(n_13605),
.B(n_11695),
.Y(n_14911)
);

AOI22xp33_ASAP7_75t_L g14912 ( 
.A1(n_13808),
.A2(n_11068),
.B1(n_13305),
.B2(n_11531),
.Y(n_14912)
);

AND2x4_ASAP7_75t_L g14913 ( 
.A(n_13653),
.B(n_10303),
.Y(n_14913)
);

AND2x2_ASAP7_75t_L g14914 ( 
.A(n_13915),
.B(n_11696),
.Y(n_14914)
);

AND2x2_ASAP7_75t_L g14915 ( 
.A(n_13840),
.B(n_11697),
.Y(n_14915)
);

AND2x2_ASAP7_75t_L g14916 ( 
.A(n_13846),
.B(n_11698),
.Y(n_14916)
);

AND2x2_ASAP7_75t_L g14917 ( 
.A(n_13759),
.B(n_11700),
.Y(n_14917)
);

AND2x2_ASAP7_75t_L g14918 ( 
.A(n_13777),
.B(n_11701),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_13546),
.Y(n_14919)
);

AND2x2_ASAP7_75t_L g14920 ( 
.A(n_13712),
.B(n_11702),
.Y(n_14920)
);

INVx1_ASAP7_75t_L g14921 ( 
.A(n_13547),
.Y(n_14921)
);

OAI22xp5_ASAP7_75t_L g14922 ( 
.A1(n_13368),
.A2(n_8376),
.B1(n_10622),
.B2(n_10578),
.Y(n_14922)
);

HB1xp67_ASAP7_75t_L g14923 ( 
.A(n_13426),
.Y(n_14923)
);

INVx2_ASAP7_75t_L g14924 ( 
.A(n_14015),
.Y(n_14924)
);

INVx1_ASAP7_75t_L g14925 ( 
.A(n_13550),
.Y(n_14925)
);

INVx1_ASAP7_75t_L g14926 ( 
.A(n_13553),
.Y(n_14926)
);

HB1xp67_ASAP7_75t_L g14927 ( 
.A(n_13429),
.Y(n_14927)
);

NAND2xp5_ASAP7_75t_L g14928 ( 
.A(n_13783),
.B(n_11709),
.Y(n_14928)
);

OR2x2_ASAP7_75t_L g14929 ( 
.A(n_13644),
.B(n_11716),
.Y(n_14929)
);

AND2x2_ASAP7_75t_L g14930 ( 
.A(n_13718),
.B(n_8296),
.Y(n_14930)
);

INVx1_ASAP7_75t_L g14931 ( 
.A(n_14021),
.Y(n_14931)
);

HB1xp67_ASAP7_75t_L g14932 ( 
.A(n_13442),
.Y(n_14932)
);

INVx1_ASAP7_75t_L g14933 ( 
.A(n_14025),
.Y(n_14933)
);

INVx1_ASAP7_75t_L g14934 ( 
.A(n_14027),
.Y(n_14934)
);

AND2x2_ASAP7_75t_L g14935 ( 
.A(n_13729),
.B(n_8296),
.Y(n_14935)
);

AND2x2_ASAP7_75t_L g14936 ( 
.A(n_13739),
.B(n_8296),
.Y(n_14936)
);

INVx2_ASAP7_75t_L g14937 ( 
.A(n_13453),
.Y(n_14937)
);

HB1xp67_ASAP7_75t_L g14938 ( 
.A(n_13456),
.Y(n_14938)
);

AND2x2_ASAP7_75t_L g14939 ( 
.A(n_13748),
.B(n_8296),
.Y(n_14939)
);

INVx2_ASAP7_75t_L g14940 ( 
.A(n_13458),
.Y(n_14940)
);

INVx1_ASAP7_75t_L g14941 ( 
.A(n_13801),
.Y(n_14941)
);

INVx1_ASAP7_75t_L g14942 ( 
.A(n_13806),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_13820),
.Y(n_14943)
);

BUFx2_ASAP7_75t_L g14944 ( 
.A(n_13703),
.Y(n_14944)
);

NAND2xp5_ASAP7_75t_L g14945 ( 
.A(n_14275),
.B(n_8933),
.Y(n_14945)
);

AND2x4_ASAP7_75t_L g14946 ( 
.A(n_13703),
.B(n_10303),
.Y(n_14946)
);

AND2x2_ASAP7_75t_L g14947 ( 
.A(n_13749),
.B(n_8296),
.Y(n_14947)
);

AOI22xp5_ASAP7_75t_L g14948 ( 
.A1(n_13496),
.A2(n_8552),
.B1(n_8550),
.B2(n_11419),
.Y(n_14948)
);

OR2x2_ASAP7_75t_L g14949 ( 
.A(n_13669),
.B(n_11721),
.Y(n_14949)
);

NAND2xp5_ASAP7_75t_L g14950 ( 
.A(n_14280),
.B(n_8933),
.Y(n_14950)
);

AND2x2_ASAP7_75t_L g14951 ( 
.A(n_13751),
.B(n_8306),
.Y(n_14951)
);

OR2x2_ASAP7_75t_L g14952 ( 
.A(n_13686),
.B(n_11724),
.Y(n_14952)
);

AND2x4_ASAP7_75t_L g14953 ( 
.A(n_13741),
.B(n_10323),
.Y(n_14953)
);

HB1xp67_ASAP7_75t_L g14954 ( 
.A(n_13468),
.Y(n_14954)
);

INVx2_ASAP7_75t_SL g14955 ( 
.A(n_13614),
.Y(n_14955)
);

NAND2xp5_ASAP7_75t_L g14956 ( 
.A(n_13845),
.B(n_8933),
.Y(n_14956)
);

AND2x2_ASAP7_75t_L g14957 ( 
.A(n_13910),
.B(n_8306),
.Y(n_14957)
);

AND2x2_ASAP7_75t_L g14958 ( 
.A(n_13912),
.B(n_8306),
.Y(n_14958)
);

INVx2_ASAP7_75t_L g14959 ( 
.A(n_13469),
.Y(n_14959)
);

HB1xp67_ASAP7_75t_L g14960 ( 
.A(n_13472),
.Y(n_14960)
);

AND2x2_ASAP7_75t_L g14961 ( 
.A(n_13709),
.B(n_8306),
.Y(n_14961)
);

INVx1_ASAP7_75t_L g14962 ( 
.A(n_13822),
.Y(n_14962)
);

AOI22xp33_ASAP7_75t_L g14963 ( 
.A1(n_14211),
.A2(n_11531),
.B1(n_11496),
.B2(n_11419),
.Y(n_14963)
);

AND2x2_ASAP7_75t_L g14964 ( 
.A(n_13964),
.B(n_8306),
.Y(n_14964)
);

INVx1_ASAP7_75t_L g14965 ( 
.A(n_13823),
.Y(n_14965)
);

AND2x4_ASAP7_75t_L g14966 ( 
.A(n_13741),
.B(n_10323),
.Y(n_14966)
);

AND2x4_ASAP7_75t_L g14967 ( 
.A(n_13939),
.B(n_10323),
.Y(n_14967)
);

NAND2xp5_ASAP7_75t_L g14968 ( 
.A(n_14283),
.B(n_8933),
.Y(n_14968)
);

INVx2_ASAP7_75t_L g14969 ( 
.A(n_13925),
.Y(n_14969)
);

INVx1_ASAP7_75t_L g14970 ( 
.A(n_13825),
.Y(n_14970)
);

AND2x2_ASAP7_75t_L g14971 ( 
.A(n_13698),
.B(n_8377),
.Y(n_14971)
);

INVx1_ASAP7_75t_L g14972 ( 
.A(n_13834),
.Y(n_14972)
);

AND2x2_ASAP7_75t_L g14973 ( 
.A(n_13704),
.B(n_8377),
.Y(n_14973)
);

OR2x2_ASAP7_75t_L g14974 ( 
.A(n_13771),
.B(n_11727),
.Y(n_14974)
);

INVx1_ASAP7_75t_L g14975 ( 
.A(n_13842),
.Y(n_14975)
);

INVx1_ASAP7_75t_L g14976 ( 
.A(n_13848),
.Y(n_14976)
);

INVx2_ASAP7_75t_L g14977 ( 
.A(n_13889),
.Y(n_14977)
);

CKINVDCx5p33_ASAP7_75t_R g14978 ( 
.A(n_13959),
.Y(n_14978)
);

NAND2xp5_ASAP7_75t_L g14979 ( 
.A(n_14014),
.B(n_8933),
.Y(n_14979)
);

NOR2xp33_ASAP7_75t_L g14980 ( 
.A(n_13939),
.B(n_6805),
.Y(n_14980)
);

BUFx3_ASAP7_75t_L g14981 ( 
.A(n_14032),
.Y(n_14981)
);

INVx1_ASAP7_75t_L g14982 ( 
.A(n_13857),
.Y(n_14982)
);

OR2x2_ASAP7_75t_L g14983 ( 
.A(n_14184),
.B(n_11729),
.Y(n_14983)
);

NAND2xp5_ASAP7_75t_L g14984 ( 
.A(n_13943),
.B(n_8933),
.Y(n_14984)
);

OR2x2_ASAP7_75t_L g14985 ( 
.A(n_14085),
.B(n_11731),
.Y(n_14985)
);

INVx1_ASAP7_75t_L g14986 ( 
.A(n_13861),
.Y(n_14986)
);

BUFx2_ASAP7_75t_L g14987 ( 
.A(n_13865),
.Y(n_14987)
);

INVx2_ASAP7_75t_L g14988 ( 
.A(n_13928),
.Y(n_14988)
);

AND2x2_ASAP7_75t_L g14989 ( 
.A(n_13772),
.B(n_8377),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_13862),
.Y(n_14990)
);

INVx1_ASAP7_75t_L g14991 ( 
.A(n_13867),
.Y(n_14991)
);

HB1xp67_ASAP7_75t_L g14992 ( 
.A(n_13435),
.Y(n_14992)
);

AND2x2_ASAP7_75t_L g14993 ( 
.A(n_13772),
.B(n_8377),
.Y(n_14993)
);

INVx1_ASAP7_75t_L g14994 ( 
.A(n_13873),
.Y(n_14994)
);

AND2x2_ASAP7_75t_L g14995 ( 
.A(n_13775),
.B(n_8377),
.Y(n_14995)
);

NOR2xp33_ASAP7_75t_L g14996 ( 
.A(n_13945),
.B(n_6883),
.Y(n_14996)
);

INVx2_ASAP7_75t_L g14997 ( 
.A(n_13937),
.Y(n_14997)
);

AND2x4_ASAP7_75t_L g14998 ( 
.A(n_13970),
.B(n_10323),
.Y(n_14998)
);

INVx1_ASAP7_75t_L g14999 ( 
.A(n_13876),
.Y(n_14999)
);

INVx1_ASAP7_75t_L g15000 ( 
.A(n_13883),
.Y(n_15000)
);

INVx3_ASAP7_75t_L g15001 ( 
.A(n_13716),
.Y(n_15001)
);

INVxp67_ASAP7_75t_SL g15002 ( 
.A(n_13916),
.Y(n_15002)
);

OR2x2_ASAP7_75t_L g15003 ( 
.A(n_14092),
.B(n_13657),
.Y(n_15003)
);

AND2x4_ASAP7_75t_L g15004 ( 
.A(n_13989),
.B(n_10387),
.Y(n_15004)
);

INVx1_ASAP7_75t_SL g15005 ( 
.A(n_13560),
.Y(n_15005)
);

INVx2_ASAP7_75t_L g15006 ( 
.A(n_13940),
.Y(n_15006)
);

INVx1_ASAP7_75t_L g15007 ( 
.A(n_13885),
.Y(n_15007)
);

AND2x4_ASAP7_75t_L g15008 ( 
.A(n_13746),
.B(n_10387),
.Y(n_15008)
);

AND2x4_ASAP7_75t_L g15009 ( 
.A(n_13746),
.B(n_10387),
.Y(n_15009)
);

OAI22xp5_ASAP7_75t_L g15010 ( 
.A1(n_14007),
.A2(n_8376),
.B1(n_10622),
.B2(n_8401),
.Y(n_15010)
);

HB1xp67_ASAP7_75t_L g15011 ( 
.A(n_13435),
.Y(n_15011)
);

INVx2_ASAP7_75t_L g15012 ( 
.A(n_13731),
.Y(n_15012)
);

AND2x2_ASAP7_75t_L g15013 ( 
.A(n_13775),
.B(n_11894),
.Y(n_15013)
);

AOI22xp33_ASAP7_75t_SL g15014 ( 
.A1(n_14245),
.A2(n_14084),
.B1(n_14215),
.B2(n_14220),
.Y(n_15014)
);

INVxp67_ASAP7_75t_SL g15015 ( 
.A(n_14174),
.Y(n_15015)
);

OR2x2_ASAP7_75t_SL g15016 ( 
.A(n_14069),
.B(n_10538),
.Y(n_15016)
);

NOR2xp33_ASAP7_75t_L g15017 ( 
.A(n_13945),
.B(n_10486),
.Y(n_15017)
);

AND2x4_ASAP7_75t_L g15018 ( 
.A(n_13716),
.B(n_10387),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_13898),
.Y(n_15019)
);

INVx2_ASAP7_75t_L g15020 ( 
.A(n_13734),
.Y(n_15020)
);

INVx4_ASAP7_75t_R g15021 ( 
.A(n_14041),
.Y(n_15021)
);

INVx1_ASAP7_75t_L g15022 ( 
.A(n_13899),
.Y(n_15022)
);

AND2x2_ASAP7_75t_L g15023 ( 
.A(n_13814),
.B(n_11894),
.Y(n_15023)
);

AND2x2_ASAP7_75t_L g15024 ( 
.A(n_13814),
.B(n_11908),
.Y(n_15024)
);

INVx1_ASAP7_75t_L g15025 ( 
.A(n_13617),
.Y(n_15025)
);

AOI22xp33_ASAP7_75t_SL g15026 ( 
.A1(n_14200),
.A2(n_11521),
.B1(n_11450),
.B2(n_11447),
.Y(n_15026)
);

INVx1_ASAP7_75t_L g15027 ( 
.A(n_13618),
.Y(n_15027)
);

INVx1_ASAP7_75t_L g15028 ( 
.A(n_13627),
.Y(n_15028)
);

INVx2_ASAP7_75t_L g15029 ( 
.A(n_13758),
.Y(n_15029)
);

NAND2xp5_ASAP7_75t_L g15030 ( 
.A(n_14118),
.B(n_8933),
.Y(n_15030)
);

OR2x2_ASAP7_75t_L g15031 ( 
.A(n_13887),
.B(n_11732),
.Y(n_15031)
);

AND2x4_ASAP7_75t_L g15032 ( 
.A(n_13560),
.B(n_10396),
.Y(n_15032)
);

INVx1_ASAP7_75t_L g15033 ( 
.A(n_13859),
.Y(n_15033)
);

HB1xp67_ASAP7_75t_L g15034 ( 
.A(n_13435),
.Y(n_15034)
);

HB1xp67_ASAP7_75t_L g15035 ( 
.A(n_13985),
.Y(n_15035)
);

INVx2_ASAP7_75t_L g15036 ( 
.A(n_13830),
.Y(n_15036)
);

HB1xp67_ASAP7_75t_L g15037 ( 
.A(n_13881),
.Y(n_15037)
);

INVx2_ASAP7_75t_SL g15038 ( 
.A(n_13614),
.Y(n_15038)
);

INVx1_ASAP7_75t_L g15039 ( 
.A(n_13863),
.Y(n_15039)
);

INVx1_ASAP7_75t_L g15040 ( 
.A(n_13878),
.Y(n_15040)
);

AND2x2_ASAP7_75t_L g15041 ( 
.A(n_13763),
.B(n_11908),
.Y(n_15041)
);

OR2x2_ASAP7_75t_L g15042 ( 
.A(n_13785),
.B(n_11737),
.Y(n_15042)
);

AND2x4_ASAP7_75t_L g15043 ( 
.A(n_13575),
.B(n_10396),
.Y(n_15043)
);

AOI22xp33_ASAP7_75t_L g15044 ( 
.A1(n_14223),
.A2(n_11531),
.B1(n_11496),
.B2(n_11419),
.Y(n_15044)
);

OR2x2_ASAP7_75t_L g15045 ( 
.A(n_13811),
.B(n_11739),
.Y(n_15045)
);

NAND2xp5_ASAP7_75t_L g15046 ( 
.A(n_14120),
.B(n_8933),
.Y(n_15046)
);

OR2x2_ASAP7_75t_L g15047 ( 
.A(n_14189),
.B(n_11748),
.Y(n_15047)
);

AND2x2_ASAP7_75t_L g15048 ( 
.A(n_13766),
.B(n_9538),
.Y(n_15048)
);

INVx1_ASAP7_75t_L g15049 ( 
.A(n_13841),
.Y(n_15049)
);

INVx3_ASAP7_75t_L g15050 ( 
.A(n_13575),
.Y(n_15050)
);

INVx2_ASAP7_75t_L g15051 ( 
.A(n_13854),
.Y(n_15051)
);

BUFx3_ASAP7_75t_L g15052 ( 
.A(n_14072),
.Y(n_15052)
);

INVx1_ASAP7_75t_L g15053 ( 
.A(n_13933),
.Y(n_15053)
);

INVx1_ASAP7_75t_L g15054 ( 
.A(n_13944),
.Y(n_15054)
);

INVx2_ASAP7_75t_L g15055 ( 
.A(n_14001),
.Y(n_15055)
);

OR2x2_ASAP7_75t_L g15056 ( 
.A(n_14291),
.B(n_11752),
.Y(n_15056)
);

AND2x2_ASAP7_75t_L g15057 ( 
.A(n_13789),
.B(n_9538),
.Y(n_15057)
);

INVx1_ASAP7_75t_L g15058 ( 
.A(n_13953),
.Y(n_15058)
);

INVx1_ASAP7_75t_L g15059 ( 
.A(n_14146),
.Y(n_15059)
);

INVx1_ASAP7_75t_L g15060 ( 
.A(n_13950),
.Y(n_15060)
);

OR2x2_ASAP7_75t_L g15061 ( 
.A(n_14235),
.B(n_11759),
.Y(n_15061)
);

INVx2_ASAP7_75t_L g15062 ( 
.A(n_14001),
.Y(n_15062)
);

INVx1_ASAP7_75t_L g15063 ( 
.A(n_13950),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_13967),
.Y(n_15064)
);

AND2x2_ASAP7_75t_L g15065 ( 
.A(n_13792),
.B(n_9538),
.Y(n_15065)
);

NAND2xp5_ASAP7_75t_L g15066 ( 
.A(n_14273),
.B(n_8966),
.Y(n_15066)
);

INVx2_ASAP7_75t_SL g15067 ( 
.A(n_13945),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_13967),
.Y(n_15068)
);

INVx1_ASAP7_75t_L g15069 ( 
.A(n_13972),
.Y(n_15069)
);

INVx1_ASAP7_75t_L g15070 ( 
.A(n_13972),
.Y(n_15070)
);

AND2x2_ASAP7_75t_L g15071 ( 
.A(n_13794),
.B(n_13795),
.Y(n_15071)
);

INVx2_ASAP7_75t_L g15072 ( 
.A(n_13947),
.Y(n_15072)
);

NAND2xp5_ASAP7_75t_L g15073 ( 
.A(n_13337),
.B(n_8966),
.Y(n_15073)
);

INVx1_ASAP7_75t_L g15074 ( 
.A(n_13978),
.Y(n_15074)
);

AND2x4_ASAP7_75t_L g15075 ( 
.A(n_13913),
.B(n_13947),
.Y(n_15075)
);

INVx2_ASAP7_75t_L g15076 ( 
.A(n_13491),
.Y(n_15076)
);

BUFx2_ASAP7_75t_L g15077 ( 
.A(n_13934),
.Y(n_15077)
);

OR2x2_ASAP7_75t_L g15078 ( 
.A(n_13818),
.B(n_11766),
.Y(n_15078)
);

INVx2_ASAP7_75t_L g15079 ( 
.A(n_13498),
.Y(n_15079)
);

INVx1_ASAP7_75t_L g15080 ( 
.A(n_13978),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_13980),
.Y(n_15081)
);

AND2x2_ASAP7_75t_L g15082 ( 
.A(n_13800),
.B(n_9539),
.Y(n_15082)
);

INVx1_ASAP7_75t_L g15083 ( 
.A(n_13980),
.Y(n_15083)
);

OR2x2_ASAP7_75t_L g15084 ( 
.A(n_13829),
.B(n_11769),
.Y(n_15084)
);

AND2x2_ASAP7_75t_L g15085 ( 
.A(n_13803),
.B(n_9539),
.Y(n_15085)
);

INVx1_ASAP7_75t_SL g15086 ( 
.A(n_13913),
.Y(n_15086)
);

INVx1_ASAP7_75t_L g15087 ( 
.A(n_13909),
.Y(n_15087)
);

AND2x2_ASAP7_75t_L g15088 ( 
.A(n_13804),
.B(n_9539),
.Y(n_15088)
);

INVx2_ASAP7_75t_SL g15089 ( 
.A(n_13549),
.Y(n_15089)
);

AND2x2_ASAP7_75t_L g15090 ( 
.A(n_13942),
.B(n_9569),
.Y(n_15090)
);

INVx2_ASAP7_75t_L g15091 ( 
.A(n_13504),
.Y(n_15091)
);

INVx3_ASAP7_75t_L g15092 ( 
.A(n_13549),
.Y(n_15092)
);

INVx1_ASAP7_75t_L g15093 ( 
.A(n_13858),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_13871),
.Y(n_15094)
);

NAND2xp5_ASAP7_75t_L g15095 ( 
.A(n_14289),
.B(n_8966),
.Y(n_15095)
);

INVx2_ASAP7_75t_L g15096 ( 
.A(n_13510),
.Y(n_15096)
);

AOI22xp33_ASAP7_75t_L g15097 ( 
.A1(n_14229),
.A2(n_11496),
.B1(n_11451),
.B2(n_11455),
.Y(n_15097)
);

INVx1_ASAP7_75t_L g15098 ( 
.A(n_13907),
.Y(n_15098)
);

INVx1_ASAP7_75t_L g15099 ( 
.A(n_13908),
.Y(n_15099)
);

INVx1_ASAP7_75t_L g15100 ( 
.A(n_14230),
.Y(n_15100)
);

INVx1_ASAP7_75t_L g15101 ( 
.A(n_14238),
.Y(n_15101)
);

INVxp33_ASAP7_75t_SL g15102 ( 
.A(n_13895),
.Y(n_15102)
);

AND2x2_ASAP7_75t_L g15103 ( 
.A(n_13949),
.B(n_13951),
.Y(n_15103)
);

AND2x2_ASAP7_75t_L g15104 ( 
.A(n_13955),
.B(n_9569),
.Y(n_15104)
);

BUFx2_ASAP7_75t_L g15105 ( 
.A(n_13865),
.Y(n_15105)
);

INVx1_ASAP7_75t_L g15106 ( 
.A(n_14243),
.Y(n_15106)
);

NAND2xp5_ASAP7_75t_L g15107 ( 
.A(n_14162),
.B(n_8966),
.Y(n_15107)
);

INVx1_ASAP7_75t_L g15108 ( 
.A(n_14248),
.Y(n_15108)
);

BUFx2_ASAP7_75t_L g15109 ( 
.A(n_14071),
.Y(n_15109)
);

INVx1_ASAP7_75t_L g15110 ( 
.A(n_14250),
.Y(n_15110)
);

BUFx3_ASAP7_75t_L g15111 ( 
.A(n_13932),
.Y(n_15111)
);

AND2x2_ASAP7_75t_L g15112 ( 
.A(n_13821),
.B(n_9569),
.Y(n_15112)
);

INVx2_ASAP7_75t_SL g15113 ( 
.A(n_13557),
.Y(n_15113)
);

CKINVDCx6p67_ASAP7_75t_R g15114 ( 
.A(n_14100),
.Y(n_15114)
);

INVx1_ASAP7_75t_L g15115 ( 
.A(n_14255),
.Y(n_15115)
);

INVx2_ASAP7_75t_L g15116 ( 
.A(n_13518),
.Y(n_15116)
);

NOR2x1_ASAP7_75t_L g15117 ( 
.A(n_14192),
.B(n_13132),
.Y(n_15117)
);

AND2x4_ASAP7_75t_SL g15118 ( 
.A(n_14019),
.B(n_7908),
.Y(n_15118)
);

BUFx2_ASAP7_75t_L g15119 ( 
.A(n_14158),
.Y(n_15119)
);

INVx2_ASAP7_75t_L g15120 ( 
.A(n_13521),
.Y(n_15120)
);

INVx1_ASAP7_75t_L g15121 ( 
.A(n_14292),
.Y(n_15121)
);

AND2x2_ASAP7_75t_L g15122 ( 
.A(n_13956),
.B(n_9580),
.Y(n_15122)
);

NAND2xp5_ASAP7_75t_L g15123 ( 
.A(n_14231),
.B(n_8966),
.Y(n_15123)
);

INVx1_ASAP7_75t_L g15124 ( 
.A(n_14112),
.Y(n_15124)
);

AND2x2_ASAP7_75t_L g15125 ( 
.A(n_13960),
.B(n_9580),
.Y(n_15125)
);

OR2x2_ASAP7_75t_L g15126 ( 
.A(n_14256),
.B(n_11772),
.Y(n_15126)
);

INVx2_ASAP7_75t_SL g15127 ( 
.A(n_13557),
.Y(n_15127)
);

INVx1_ASAP7_75t_L g15128 ( 
.A(n_13927),
.Y(n_15128)
);

AND2x2_ASAP7_75t_L g15129 ( 
.A(n_14057),
.B(n_9580),
.Y(n_15129)
);

AND2x2_ASAP7_75t_L g15130 ( 
.A(n_14073),
.B(n_14046),
.Y(n_15130)
);

OR2x2_ASAP7_75t_L g15131 ( 
.A(n_14199),
.B(n_11773),
.Y(n_15131)
);

AND2x2_ASAP7_75t_L g15132 ( 
.A(n_14044),
.B(n_9165),
.Y(n_15132)
);

BUFx6f_ASAP7_75t_L g15133 ( 
.A(n_13891),
.Y(n_15133)
);

NAND2xp5_ASAP7_75t_L g15134 ( 
.A(n_14227),
.B(n_8966),
.Y(n_15134)
);

INVx2_ASAP7_75t_L g15135 ( 
.A(n_13522),
.Y(n_15135)
);

INVx1_ASAP7_75t_L g15136 ( 
.A(n_13927),
.Y(n_15136)
);

AND2x2_ASAP7_75t_L g15137 ( 
.A(n_14094),
.B(n_9165),
.Y(n_15137)
);

AND2x2_ASAP7_75t_L g15138 ( 
.A(n_14179),
.B(n_9165),
.Y(n_15138)
);

BUFx2_ASAP7_75t_SL g15139 ( 
.A(n_14341),
.Y(n_15139)
);

AND2x4_ASAP7_75t_SL g15140 ( 
.A(n_14305),
.B(n_13891),
.Y(n_15140)
);

INVx2_ASAP7_75t_L g15141 ( 
.A(n_14884),
.Y(n_15141)
);

AND2x2_ASAP7_75t_L g15142 ( 
.A(n_14394),
.B(n_14224),
.Y(n_15142)
);

HB1xp67_ASAP7_75t_L g15143 ( 
.A(n_15109),
.Y(n_15143)
);

INVx2_ASAP7_75t_L g15144 ( 
.A(n_14485),
.Y(n_15144)
);

AND2x2_ASAP7_75t_L g15145 ( 
.A(n_14346),
.B(n_14224),
.Y(n_15145)
);

INVx2_ASAP7_75t_L g15146 ( 
.A(n_14485),
.Y(n_15146)
);

INVxp67_ASAP7_75t_L g15147 ( 
.A(n_14305),
.Y(n_15147)
);

AND2x2_ASAP7_75t_L g15148 ( 
.A(n_14350),
.B(n_14116),
.Y(n_15148)
);

NAND2xp5_ASAP7_75t_L g15149 ( 
.A(n_14373),
.B(n_14216),
.Y(n_15149)
);

INVx2_ASAP7_75t_L g15150 ( 
.A(n_14489),
.Y(n_15150)
);

AND2x2_ASAP7_75t_L g15151 ( 
.A(n_14407),
.B(n_14191),
.Y(n_15151)
);

INVxp67_ASAP7_75t_L g15152 ( 
.A(n_15119),
.Y(n_15152)
);

NOR2xp33_ASAP7_75t_L g15153 ( 
.A(n_14411),
.B(n_14192),
.Y(n_15153)
);

OR2x2_ASAP7_75t_L g15154 ( 
.A(n_14488),
.B(n_14202),
.Y(n_15154)
);

INVx1_ASAP7_75t_L g15155 ( 
.A(n_14475),
.Y(n_15155)
);

BUFx2_ASAP7_75t_SL g15156 ( 
.A(n_14300),
.Y(n_15156)
);

AND2x4_ASAP7_75t_L g15157 ( 
.A(n_14301),
.B(n_14107),
.Y(n_15157)
);

HB1xp67_ASAP7_75t_L g15158 ( 
.A(n_14987),
.Y(n_15158)
);

AND2x2_ASAP7_75t_L g15159 ( 
.A(n_14301),
.B(n_14134),
.Y(n_15159)
);

INVx2_ASAP7_75t_SL g15160 ( 
.A(n_14670),
.Y(n_15160)
);

BUFx2_ASAP7_75t_L g15161 ( 
.A(n_14987),
.Y(n_15161)
);

INVx1_ASAP7_75t_L g15162 ( 
.A(n_14641),
.Y(n_15162)
);

INVx1_ASAP7_75t_L g15163 ( 
.A(n_14649),
.Y(n_15163)
);

INVx2_ASAP7_75t_L g15164 ( 
.A(n_14495),
.Y(n_15164)
);

INVx2_ASAP7_75t_L g15165 ( 
.A(n_14555),
.Y(n_15165)
);

INVx2_ASAP7_75t_L g15166 ( 
.A(n_14601),
.Y(n_15166)
);

AND2x2_ASAP7_75t_L g15167 ( 
.A(n_14379),
.B(n_14134),
.Y(n_15167)
);

AND2x2_ASAP7_75t_L g15168 ( 
.A(n_14625),
.B(n_14134),
.Y(n_15168)
);

INVx1_ASAP7_75t_L g15169 ( 
.A(n_14684),
.Y(n_15169)
);

INVx1_ASAP7_75t_L g15170 ( 
.A(n_14699),
.Y(n_15170)
);

NAND2xp5_ASAP7_75t_L g15171 ( 
.A(n_14311),
.B(n_14117),
.Y(n_15171)
);

INVx1_ASAP7_75t_L g15172 ( 
.A(n_14340),
.Y(n_15172)
);

INVx5_ASAP7_75t_L g15173 ( 
.A(n_14389),
.Y(n_15173)
);

INVx1_ASAP7_75t_L g15174 ( 
.A(n_14344),
.Y(n_15174)
);

BUFx3_ASAP7_75t_L g15175 ( 
.A(n_14406),
.Y(n_15175)
);

INVx1_ASAP7_75t_L g15176 ( 
.A(n_14571),
.Y(n_15176)
);

AND2x2_ASAP7_75t_L g15177 ( 
.A(n_14328),
.B(n_14083),
.Y(n_15177)
);

INVx5_ASAP7_75t_L g15178 ( 
.A(n_14776),
.Y(n_15178)
);

INVx2_ASAP7_75t_L g15179 ( 
.A(n_14615),
.Y(n_15179)
);

NAND2xp5_ASAP7_75t_L g15180 ( 
.A(n_14349),
.B(n_14095),
.Y(n_15180)
);

INVx1_ASAP7_75t_L g15181 ( 
.A(n_14585),
.Y(n_15181)
);

INVx5_ASAP7_75t_L g15182 ( 
.A(n_14776),
.Y(n_15182)
);

INVx2_ASAP7_75t_L g15183 ( 
.A(n_14447),
.Y(n_15183)
);

AND2x2_ASAP7_75t_L g15184 ( 
.A(n_14806),
.B(n_13987),
.Y(n_15184)
);

HB1xp67_ASAP7_75t_L g15185 ( 
.A(n_15105),
.Y(n_15185)
);

OR2x2_ASAP7_75t_L g15186 ( 
.A(n_14530),
.B(n_14129),
.Y(n_15186)
);

INVx1_ASAP7_75t_L g15187 ( 
.A(n_14619),
.Y(n_15187)
);

OAI21xp33_ASAP7_75t_L g15188 ( 
.A1(n_14563),
.A2(n_14106),
.B(n_14047),
.Y(n_15188)
);

INVx4_ASAP7_75t_L g15189 ( 
.A(n_14436),
.Y(n_15189)
);

AND2x2_ASAP7_75t_L g15190 ( 
.A(n_14607),
.B(n_13988),
.Y(n_15190)
);

INVx3_ASAP7_75t_L g15191 ( 
.A(n_14400),
.Y(n_15191)
);

OR2x6_ASAP7_75t_L g15192 ( 
.A(n_14307),
.B(n_13364),
.Y(n_15192)
);

INVx2_ASAP7_75t_L g15193 ( 
.A(n_14512),
.Y(n_15193)
);

AND2x2_ASAP7_75t_L g15194 ( 
.A(n_14388),
.B(n_13890),
.Y(n_15194)
);

HB1xp67_ASAP7_75t_L g15195 ( 
.A(n_15105),
.Y(n_15195)
);

INVx1_ASAP7_75t_L g15196 ( 
.A(n_14992),
.Y(n_15196)
);

INVx2_ASAP7_75t_L g15197 ( 
.A(n_14536),
.Y(n_15197)
);

AOI22xp5_ASAP7_75t_L g15198 ( 
.A1(n_14378),
.A2(n_14161),
.B1(n_14153),
.B2(n_13514),
.Y(n_15198)
);

INVx5_ASAP7_75t_SL g15199 ( 
.A(n_15114),
.Y(n_15199)
);

INVxp67_ASAP7_75t_SL g15200 ( 
.A(n_14549),
.Y(n_15200)
);

INVx2_ASAP7_75t_L g15201 ( 
.A(n_14552),
.Y(n_15201)
);

OR2x6_ASAP7_75t_L g15202 ( 
.A(n_14472),
.B(n_13526),
.Y(n_15202)
);

BUFx6f_ASAP7_75t_L g15203 ( 
.A(n_14364),
.Y(n_15203)
);

INVx3_ASAP7_75t_L g15204 ( 
.A(n_14581),
.Y(n_15204)
);

AND2x2_ASAP7_75t_L g15205 ( 
.A(n_14387),
.B(n_13974),
.Y(n_15205)
);

AND2x2_ASAP7_75t_L g15206 ( 
.A(n_14304),
.B(n_13982),
.Y(n_15206)
);

INVx1_ASAP7_75t_L g15207 ( 
.A(n_15011),
.Y(n_15207)
);

INVx2_ASAP7_75t_L g15208 ( 
.A(n_14342),
.Y(n_15208)
);

INVx1_ASAP7_75t_L g15209 ( 
.A(n_15034),
.Y(n_15209)
);

BUFx3_ASAP7_75t_L g15210 ( 
.A(n_14894),
.Y(n_15210)
);

INVx1_ASAP7_75t_L g15211 ( 
.A(n_14629),
.Y(n_15211)
);

AND2x2_ASAP7_75t_L g15212 ( 
.A(n_14799),
.B(n_14111),
.Y(n_15212)
);

INVx2_ASAP7_75t_L g15213 ( 
.A(n_14610),
.Y(n_15213)
);

INVx1_ASAP7_75t_L g15214 ( 
.A(n_14424),
.Y(n_15214)
);

AND2x2_ASAP7_75t_L g15215 ( 
.A(n_14403),
.B(n_14004),
.Y(n_15215)
);

INVx1_ASAP7_75t_L g15216 ( 
.A(n_14860),
.Y(n_15216)
);

INVx3_ASAP7_75t_L g15217 ( 
.A(n_14581),
.Y(n_15217)
);

BUFx3_ASAP7_75t_L g15218 ( 
.A(n_14766),
.Y(n_15218)
);

BUFx2_ASAP7_75t_L g15219 ( 
.A(n_14329),
.Y(n_15219)
);

INVx2_ASAP7_75t_L g15220 ( 
.A(n_14510),
.Y(n_15220)
);

AOI22xp33_ASAP7_75t_L g15221 ( 
.A1(n_14454),
.A2(n_13901),
.B1(n_14197),
.B2(n_14198),
.Y(n_15221)
);

INVx2_ASAP7_75t_L g15222 ( 
.A(n_14587),
.Y(n_15222)
);

AND2x2_ASAP7_75t_L g15223 ( 
.A(n_14434),
.B(n_14005),
.Y(n_15223)
);

INVx1_ASAP7_75t_L g15224 ( 
.A(n_14748),
.Y(n_15224)
);

AND2x2_ASAP7_75t_L g15225 ( 
.A(n_14981),
.B(n_14099),
.Y(n_15225)
);

HB1xp67_ASAP7_75t_L g15226 ( 
.A(n_14312),
.Y(n_15226)
);

INVxp67_ASAP7_75t_SL g15227 ( 
.A(n_14329),
.Y(n_15227)
);

INVx1_ASAP7_75t_L g15228 ( 
.A(n_15033),
.Y(n_15228)
);

AND2x2_ASAP7_75t_L g15229 ( 
.A(n_14773),
.B(n_14177),
.Y(n_15229)
);

AND2x2_ASAP7_75t_L g15230 ( 
.A(n_14518),
.B(n_13962),
.Y(n_15230)
);

AND2x2_ASAP7_75t_L g15231 ( 
.A(n_14900),
.B(n_13966),
.Y(n_15231)
);

INVxp67_ASAP7_75t_L g15232 ( 
.A(n_14359),
.Y(n_15232)
);

OR2x2_ASAP7_75t_L g15233 ( 
.A(n_14327),
.B(n_13924),
.Y(n_15233)
);

BUFx2_ASAP7_75t_L g15234 ( 
.A(n_14374),
.Y(n_15234)
);

INVx2_ASAP7_75t_L g15235 ( 
.A(n_14626),
.Y(n_15235)
);

AOI22xp33_ASAP7_75t_L g15236 ( 
.A1(n_14385),
.A2(n_14221),
.B1(n_14237),
.B2(n_13819),
.Y(n_15236)
);

INVx1_ASAP7_75t_L g15237 ( 
.A(n_15039),
.Y(n_15237)
);

AND2x2_ASAP7_75t_L g15238 ( 
.A(n_14310),
.B(n_13969),
.Y(n_15238)
);

AND2x2_ASAP7_75t_L g15239 ( 
.A(n_14368),
.B(n_13971),
.Y(n_15239)
);

NAND2xp5_ASAP7_75t_L g15240 ( 
.A(n_14327),
.B(n_14160),
.Y(n_15240)
);

BUFx3_ASAP7_75t_L g15241 ( 
.A(n_14646),
.Y(n_15241)
);

BUFx6f_ASAP7_75t_L g15242 ( 
.A(n_14436),
.Y(n_15242)
);

INVx2_ASAP7_75t_L g15243 ( 
.A(n_14436),
.Y(n_15243)
);

INVx1_ASAP7_75t_L g15244 ( 
.A(n_15040),
.Y(n_15244)
);

INVxp67_ASAP7_75t_SL g15245 ( 
.A(n_14575),
.Y(n_15245)
);

INVx2_ASAP7_75t_L g15246 ( 
.A(n_14872),
.Y(n_15246)
);

INVx1_ASAP7_75t_L g15247 ( 
.A(n_14360),
.Y(n_15247)
);

INVx2_ASAP7_75t_L g15248 ( 
.A(n_14502),
.Y(n_15248)
);

INVx1_ASAP7_75t_L g15249 ( 
.A(n_14361),
.Y(n_15249)
);

INVx1_ASAP7_75t_L g15250 ( 
.A(n_14362),
.Y(n_15250)
);

INVx1_ASAP7_75t_L g15251 ( 
.A(n_14366),
.Y(n_15251)
);

NAND2xp5_ASAP7_75t_L g15252 ( 
.A(n_15052),
.B(n_13340),
.Y(n_15252)
);

OR2x2_ASAP7_75t_L g15253 ( 
.A(n_14522),
.B(n_13813),
.Y(n_15253)
);

INVx2_ASAP7_75t_L g15254 ( 
.A(n_14502),
.Y(n_15254)
);

AND2x2_ASAP7_75t_L g15255 ( 
.A(n_14554),
.B(n_14009),
.Y(n_15255)
);

INVx2_ASAP7_75t_L g15256 ( 
.A(n_14486),
.Y(n_15256)
);

AND2x4_ASAP7_75t_L g15257 ( 
.A(n_14599),
.B(n_14077),
.Y(n_15257)
);

INVx2_ASAP7_75t_L g15258 ( 
.A(n_15092),
.Y(n_15258)
);

INVx1_ASAP7_75t_L g15259 ( 
.A(n_14314),
.Y(n_15259)
);

OR2x2_ASAP7_75t_L g15260 ( 
.A(n_14474),
.B(n_13843),
.Y(n_15260)
);

NAND2x1p5_ASAP7_75t_SL g15261 ( 
.A(n_15067),
.B(n_13543),
.Y(n_15261)
);

INVx1_ASAP7_75t_SL g15262 ( 
.A(n_15130),
.Y(n_15262)
);

AND2x2_ASAP7_75t_L g15263 ( 
.A(n_14419),
.B(n_14031),
.Y(n_15263)
);

AO21x2_ASAP7_75t_L g15264 ( 
.A1(n_14645),
.A2(n_14022),
.B(n_13963),
.Y(n_15264)
);

INVx2_ASAP7_75t_L g15265 ( 
.A(n_15016),
.Y(n_15265)
);

HB1xp67_ASAP7_75t_L g15266 ( 
.A(n_14792),
.Y(n_15266)
);

INVx2_ASAP7_75t_L g15267 ( 
.A(n_15050),
.Y(n_15267)
);

BUFx3_ASAP7_75t_L g15268 ( 
.A(n_14727),
.Y(n_15268)
);

INVx2_ASAP7_75t_L g15269 ( 
.A(n_14323),
.Y(n_15269)
);

AOI33xp33_ASAP7_75t_L g15270 ( 
.A1(n_14309),
.A2(n_13602),
.A3(n_14218),
.B1(n_13810),
.B2(n_14002),
.B3(n_13334),
.Y(n_15270)
);

AND2x2_ASAP7_75t_L g15271 ( 
.A(n_14639),
.B(n_14299),
.Y(n_15271)
);

HB1xp67_ASAP7_75t_L g15272 ( 
.A(n_14828),
.Y(n_15272)
);

AND2x2_ASAP7_75t_L g15273 ( 
.A(n_14442),
.B(n_14053),
.Y(n_15273)
);

HB1xp67_ASAP7_75t_L g15274 ( 
.A(n_14439),
.Y(n_15274)
);

AND2x2_ASAP7_75t_L g15275 ( 
.A(n_14408),
.B(n_14169),
.Y(n_15275)
);

BUFx3_ASAP7_75t_L g15276 ( 
.A(n_14727),
.Y(n_15276)
);

INVx1_ASAP7_75t_L g15277 ( 
.A(n_15053),
.Y(n_15277)
);

INVxp67_ASAP7_75t_L g15278 ( 
.A(n_14826),
.Y(n_15278)
);

INVx4_ASAP7_75t_L g15279 ( 
.A(n_14885),
.Y(n_15279)
);

CKINVDCx20_ASAP7_75t_R g15280 ( 
.A(n_14477),
.Y(n_15280)
);

INVx1_ASAP7_75t_L g15281 ( 
.A(n_15054),
.Y(n_15281)
);

AND2x2_ASAP7_75t_L g15282 ( 
.A(n_15103),
.B(n_13941),
.Y(n_15282)
);

AND2x2_ASAP7_75t_L g15283 ( 
.A(n_14351),
.B(n_14039),
.Y(n_15283)
);

AND2x2_ASAP7_75t_L g15284 ( 
.A(n_14371),
.B(n_13566),
.Y(n_15284)
);

OR2x2_ASAP7_75t_L g15285 ( 
.A(n_14831),
.B(n_14168),
.Y(n_15285)
);

INVx1_ASAP7_75t_SL g15286 ( 
.A(n_15005),
.Y(n_15286)
);

BUFx6f_ASAP7_75t_L g15287 ( 
.A(n_14674),
.Y(n_15287)
);

INVx1_ASAP7_75t_L g15288 ( 
.A(n_15058),
.Y(n_15288)
);

OR2x2_ASAP7_75t_L g15289 ( 
.A(n_14835),
.B(n_14282),
.Y(n_15289)
);

INVx2_ASAP7_75t_L g15290 ( 
.A(n_14326),
.Y(n_15290)
);

INVx5_ASAP7_75t_SL g15291 ( 
.A(n_14472),
.Y(n_15291)
);

NAND2xp5_ASAP7_75t_L g15292 ( 
.A(n_14561),
.B(n_13991),
.Y(n_15292)
);

INVx1_ASAP7_75t_L g15293 ( 
.A(n_15098),
.Y(n_15293)
);

HB1xp67_ASAP7_75t_L g15294 ( 
.A(n_14535),
.Y(n_15294)
);

INVx2_ASAP7_75t_L g15295 ( 
.A(n_14370),
.Y(n_15295)
);

NAND4xp25_ASAP7_75t_L g15296 ( 
.A(n_15102),
.B(n_14170),
.C(n_13929),
.D(n_13539),
.Y(n_15296)
);

OR2x2_ASAP7_75t_L g15297 ( 
.A(n_14685),
.B(n_13865),
.Y(n_15297)
);

INVx1_ASAP7_75t_L g15298 ( 
.A(n_15099),
.Y(n_15298)
);

INVxp67_ASAP7_75t_SL g15299 ( 
.A(n_14693),
.Y(n_15299)
);

AND2x4_ASAP7_75t_L g15300 ( 
.A(n_14437),
.B(n_14078),
.Y(n_15300)
);

AND2x2_ASAP7_75t_L g15301 ( 
.A(n_15071),
.B(n_14080),
.Y(n_15301)
);

INVx2_ASAP7_75t_L g15302 ( 
.A(n_15133),
.Y(n_15302)
);

HB1xp67_ASAP7_75t_L g15303 ( 
.A(n_14569),
.Y(n_15303)
);

INVx2_ASAP7_75t_L g15304 ( 
.A(n_15133),
.Y(n_15304)
);

AND2x2_ASAP7_75t_L g15305 ( 
.A(n_14413),
.B(n_14201),
.Y(n_15305)
);

INVx3_ASAP7_75t_L g15306 ( 
.A(n_14606),
.Y(n_15306)
);

NAND2xp5_ASAP7_75t_L g15307 ( 
.A(n_15015),
.B(n_13352),
.Y(n_15307)
);

AOI221xp5_ASAP7_75t_L g15308 ( 
.A1(n_14302),
.A2(n_13540),
.B1(n_14040),
.B2(n_13551),
.C(n_14166),
.Y(n_15308)
);

INVx1_ASAP7_75t_L g15309 ( 
.A(n_14505),
.Y(n_15309)
);

AOI221xp5_ASAP7_75t_L g15310 ( 
.A1(n_14375),
.A2(n_13735),
.B1(n_14290),
.B2(n_13844),
.C(n_14225),
.Y(n_15310)
);

INVx1_ASAP7_75t_L g15311 ( 
.A(n_14511),
.Y(n_15311)
);

HB1xp67_ASAP7_75t_L g15312 ( 
.A(n_14576),
.Y(n_15312)
);

INVx1_ASAP7_75t_L g15313 ( 
.A(n_14514),
.Y(n_15313)
);

INVx1_ASAP7_75t_L g15314 ( 
.A(n_14517),
.Y(n_15314)
);

AND2x2_ASAP7_75t_L g15315 ( 
.A(n_14417),
.B(n_14240),
.Y(n_15315)
);

AND2x2_ASAP7_75t_L g15316 ( 
.A(n_14418),
.B(n_13888),
.Y(n_15316)
);

AND2x2_ASAP7_75t_L g15317 ( 
.A(n_14741),
.B(n_14244),
.Y(n_15317)
);

INVx1_ASAP7_75t_L g15318 ( 
.A(n_14367),
.Y(n_15318)
);

OR2x2_ASAP7_75t_L g15319 ( 
.A(n_14685),
.B(n_14156),
.Y(n_15319)
);

INVx4_ASAP7_75t_L g15320 ( 
.A(n_14978),
.Y(n_15320)
);

INVx2_ASAP7_75t_L g15321 ( 
.A(n_14316),
.Y(n_15321)
);

AO22x1_ASAP7_75t_L g15322 ( 
.A1(n_14589),
.A2(n_14608),
.B1(n_15117),
.B2(n_14785),
.Y(n_15322)
);

INVx1_ASAP7_75t_L g15323 ( 
.A(n_14380),
.Y(n_15323)
);

AND2x2_ASAP7_75t_L g15324 ( 
.A(n_14591),
.B(n_14108),
.Y(n_15324)
);

AND2x2_ASAP7_75t_L g15325 ( 
.A(n_14308),
.B(n_14183),
.Y(n_15325)
);

AND2x2_ASAP7_75t_L g15326 ( 
.A(n_14453),
.B(n_14096),
.Y(n_15326)
);

OAI22xp5_ASAP7_75t_L g15327 ( 
.A1(n_14476),
.A2(n_13502),
.B1(n_14249),
.B2(n_14296),
.Y(n_15327)
);

INVx1_ASAP7_75t_L g15328 ( 
.A(n_14393),
.Y(n_15328)
);

INVx2_ASAP7_75t_L g15329 ( 
.A(n_15089),
.Y(n_15329)
);

INVx5_ASAP7_75t_L g15330 ( 
.A(n_14734),
.Y(n_15330)
);

AO21x2_ASAP7_75t_L g15331 ( 
.A1(n_14871),
.A2(n_13973),
.B(n_13958),
.Y(n_15331)
);

NAND2xp5_ASAP7_75t_L g15332 ( 
.A(n_14465),
.B(n_14691),
.Y(n_15332)
);

INVx2_ASAP7_75t_L g15333 ( 
.A(n_15113),
.Y(n_15333)
);

INVx2_ASAP7_75t_L g15334 ( 
.A(n_15127),
.Y(n_15334)
);

AND2x4_ASAP7_75t_L g15335 ( 
.A(n_14437),
.B(n_14456),
.Y(n_15335)
);

NOR2x1_ASAP7_75t_R g15336 ( 
.A(n_14840),
.B(n_14635),
.Y(n_15336)
);

OR2x2_ASAP7_75t_L g15337 ( 
.A(n_14721),
.B(n_14652),
.Y(n_15337)
);

INVx2_ASAP7_75t_L g15338 ( 
.A(n_14877),
.Y(n_15338)
);

NAND2xp5_ASAP7_75t_L g15339 ( 
.A(n_14738),
.B(n_14143),
.Y(n_15339)
);

INVxp67_ASAP7_75t_SL g15340 ( 
.A(n_14696),
.Y(n_15340)
);

INVx1_ASAP7_75t_L g15341 ( 
.A(n_14637),
.Y(n_15341)
);

INVx1_ASAP7_75t_L g15342 ( 
.A(n_14638),
.Y(n_15342)
);

INVx1_ASAP7_75t_L g15343 ( 
.A(n_14650),
.Y(n_15343)
);

INVx1_ASAP7_75t_L g15344 ( 
.A(n_14931),
.Y(n_15344)
);

INVx2_ASAP7_75t_L g15345 ( 
.A(n_14504),
.Y(n_15345)
);

INVx1_ASAP7_75t_L g15346 ( 
.A(n_14933),
.Y(n_15346)
);

INVx2_ASAP7_75t_L g15347 ( 
.A(n_14519),
.Y(n_15347)
);

INVx1_ASAP7_75t_L g15348 ( 
.A(n_14934),
.Y(n_15348)
);

AND2x2_ASAP7_75t_L g15349 ( 
.A(n_14461),
.B(n_14463),
.Y(n_15349)
);

INVxp67_ASAP7_75t_SL g15350 ( 
.A(n_14955),
.Y(n_15350)
);

AND2x2_ASAP7_75t_L g15351 ( 
.A(n_14422),
.B(n_14066),
.Y(n_15351)
);

INVx2_ASAP7_75t_L g15352 ( 
.A(n_14449),
.Y(n_15352)
);

INVx2_ASAP7_75t_L g15353 ( 
.A(n_15001),
.Y(n_15353)
);

INVx3_ASAP7_75t_L g15354 ( 
.A(n_14606),
.Y(n_15354)
);

INVx1_ASAP7_75t_L g15355 ( 
.A(n_14633),
.Y(n_15355)
);

INVx2_ASAP7_75t_L g15356 ( 
.A(n_14909),
.Y(n_15356)
);

INVx1_ASAP7_75t_L g15357 ( 
.A(n_14636),
.Y(n_15357)
);

HB1xp67_ASAP7_75t_L g15358 ( 
.A(n_14944),
.Y(n_15358)
);

AND2x2_ASAP7_75t_L g15359 ( 
.A(n_14423),
.B(n_14035),
.Y(n_15359)
);

INVx2_ASAP7_75t_L g15360 ( 
.A(n_14507),
.Y(n_15360)
);

INVx1_ASAP7_75t_L g15361 ( 
.A(n_14492),
.Y(n_15361)
);

NAND4xp25_ASAP7_75t_L g15362 ( 
.A(n_15003),
.B(n_14214),
.C(n_13911),
.D(n_13428),
.Y(n_15362)
);

AND2x2_ASAP7_75t_L g15363 ( 
.A(n_14412),
.B(n_14038),
.Y(n_15363)
);

AND2x4_ASAP7_75t_L g15364 ( 
.A(n_14456),
.B(n_13952),
.Y(n_15364)
);

BUFx2_ASAP7_75t_L g15365 ( 
.A(n_15038),
.Y(n_15365)
);

INVx1_ASAP7_75t_L g15366 ( 
.A(n_14498),
.Y(n_15366)
);

HB1xp67_ASAP7_75t_L g15367 ( 
.A(n_14746),
.Y(n_15367)
);

INVxp67_ASAP7_75t_L g15368 ( 
.A(n_14557),
.Y(n_15368)
);

OR2x2_ASAP7_75t_L g15369 ( 
.A(n_14444),
.B(n_13383),
.Y(n_15369)
);

INVx1_ASAP7_75t_L g15370 ( 
.A(n_15049),
.Y(n_15370)
);

AND2x2_ASAP7_75t_L g15371 ( 
.A(n_14556),
.B(n_14042),
.Y(n_15371)
);

INVx2_ASAP7_75t_L g15372 ( 
.A(n_14565),
.Y(n_15372)
);

AOI22xp5_ASAP7_75t_L g15373 ( 
.A1(n_14487),
.A2(n_14204),
.B1(n_14110),
.B2(n_14135),
.Y(n_15373)
);

INVxp67_ASAP7_75t_SL g15374 ( 
.A(n_14382),
.Y(n_15374)
);

INVx1_ASAP7_75t_L g15375 ( 
.A(n_14478),
.Y(n_15375)
);

BUFx2_ASAP7_75t_L g15376 ( 
.A(n_15002),
.Y(n_15376)
);

HB1xp67_ASAP7_75t_L g15377 ( 
.A(n_14853),
.Y(n_15377)
);

AOI22xp33_ASAP7_75t_L g15378 ( 
.A1(n_14390),
.A2(n_14102),
.B1(n_14148),
.B2(n_14145),
.Y(n_15378)
);

NOR2x1_ASAP7_75t_L g15379 ( 
.A(n_14525),
.B(n_13952),
.Y(n_15379)
);

AND2x2_ASAP7_75t_L g15380 ( 
.A(n_14521),
.B(n_14125),
.Y(n_15380)
);

OR2x2_ASAP7_75t_L g15381 ( 
.A(n_14586),
.B(n_14543),
.Y(n_15381)
);

INVx1_ASAP7_75t_L g15382 ( 
.A(n_14480),
.Y(n_15382)
);

INVx1_ASAP7_75t_L g15383 ( 
.A(n_14847),
.Y(n_15383)
);

INVx2_ASAP7_75t_L g15384 ( 
.A(n_14565),
.Y(n_15384)
);

OR2x2_ASAP7_75t_L g15385 ( 
.A(n_14473),
.B(n_14000),
.Y(n_15385)
);

INVx2_ASAP7_75t_L g15386 ( 
.A(n_14523),
.Y(n_15386)
);

AND2x2_ASAP7_75t_L g15387 ( 
.A(n_15129),
.B(n_14155),
.Y(n_15387)
);

INVx3_ASAP7_75t_L g15388 ( 
.A(n_14621),
.Y(n_15388)
);

INVx1_ASAP7_75t_L g15389 ( 
.A(n_15012),
.Y(n_15389)
);

AO21x2_ASAP7_75t_L g15390 ( 
.A1(n_14592),
.A2(n_14781),
.B(n_14395),
.Y(n_15390)
);

INVx1_ASAP7_75t_L g15391 ( 
.A(n_15020),
.Y(n_15391)
);

INVx1_ASAP7_75t_L g15392 ( 
.A(n_15029),
.Y(n_15392)
);

OR2x2_ASAP7_75t_L g15393 ( 
.A(n_14985),
.B(n_14003),
.Y(n_15393)
);

NAND2xp5_ASAP7_75t_L g15394 ( 
.A(n_14977),
.B(n_13630),
.Y(n_15394)
);

AND2x2_ASAP7_75t_L g15395 ( 
.A(n_14838),
.B(n_14203),
.Y(n_15395)
);

OAI32xp33_ASAP7_75t_L g15396 ( 
.A1(n_14322),
.A2(n_14241),
.A3(n_14284),
.B1(n_13423),
.B2(n_14247),
.Y(n_15396)
);

NAND2xp5_ASAP7_75t_L g15397 ( 
.A(n_14614),
.B(n_13935),
.Y(n_15397)
);

AND2x2_ASAP7_75t_L g15398 ( 
.A(n_14333),
.B(n_13981),
.Y(n_15398)
);

INVx1_ASAP7_75t_L g15399 ( 
.A(n_15035),
.Y(n_15399)
);

OR2x2_ASAP7_75t_L g15400 ( 
.A(n_14631),
.B(n_14765),
.Y(n_15400)
);

INVx1_ASAP7_75t_L g15401 ( 
.A(n_14508),
.Y(n_15401)
);

NAND2xp5_ASAP7_75t_L g15402 ( 
.A(n_14914),
.B(n_13935),
.Y(n_15402)
);

AND2x2_ASAP7_75t_L g15403 ( 
.A(n_14856),
.B(n_13981),
.Y(n_15403)
);

OR2x2_ASAP7_75t_L g15404 ( 
.A(n_14572),
.B(n_14024),
.Y(n_15404)
);

INVx1_ASAP7_75t_L g15405 ( 
.A(n_14597),
.Y(n_15405)
);

BUFx2_ASAP7_75t_L g15406 ( 
.A(n_15077),
.Y(n_15406)
);

NAND2xp5_ASAP7_75t_L g15407 ( 
.A(n_14774),
.B(n_14819),
.Y(n_15407)
);

INVxp33_ASAP7_75t_L g15408 ( 
.A(n_14996),
.Y(n_15408)
);

OR2x2_ASAP7_75t_L g15409 ( 
.A(n_15037),
.B(n_14063),
.Y(n_15409)
);

AND2x2_ASAP7_75t_L g15410 ( 
.A(n_14857),
.B(n_13999),
.Y(n_15410)
);

INVx1_ASAP7_75t_L g15411 ( 
.A(n_14441),
.Y(n_15411)
);

INVx3_ASAP7_75t_L g15412 ( 
.A(n_14621),
.Y(n_15412)
);

AND2x2_ASAP7_75t_L g15413 ( 
.A(n_14858),
.B(n_13999),
.Y(n_15413)
);

INVx2_ASAP7_75t_SL g15414 ( 
.A(n_14613),
.Y(n_15414)
);

INVx1_ASAP7_75t_L g15415 ( 
.A(n_14750),
.Y(n_15415)
);

INVx1_ASAP7_75t_L g15416 ( 
.A(n_14772),
.Y(n_15416)
);

INVx2_ASAP7_75t_L g15417 ( 
.A(n_14531),
.Y(n_15417)
);

AND2x2_ASAP7_75t_L g15418 ( 
.A(n_14873),
.B(n_14874),
.Y(n_15418)
);

BUFx2_ASAP7_75t_L g15419 ( 
.A(n_14544),
.Y(n_15419)
);

BUFx2_ASAP7_75t_L g15420 ( 
.A(n_14544),
.Y(n_15420)
);

INVx1_ASAP7_75t_L g15421 ( 
.A(n_14796),
.Y(n_15421)
);

AND2x2_ASAP7_75t_L g15422 ( 
.A(n_14879),
.B(n_14698),
.Y(n_15422)
);

HB1xp67_ASAP7_75t_L g15423 ( 
.A(n_14534),
.Y(n_15423)
);

INVx2_ASAP7_75t_L g15424 ( 
.A(n_14672),
.Y(n_15424)
);

INVx3_ASAP7_75t_L g15425 ( 
.A(n_15032),
.Y(n_15425)
);

HB1xp67_ASAP7_75t_L g15426 ( 
.A(n_14593),
.Y(n_15426)
);

AND2x2_ASAP7_75t_L g15427 ( 
.A(n_14846),
.B(n_14219),
.Y(n_15427)
);

INVx2_ASAP7_75t_L g15428 ( 
.A(n_14767),
.Y(n_15428)
);

INVx2_ASAP7_75t_L g15429 ( 
.A(n_14482),
.Y(n_15429)
);

BUFx3_ASAP7_75t_L g15430 ( 
.A(n_14802),
.Y(n_15430)
);

INVx2_ASAP7_75t_SL g15431 ( 
.A(n_15021),
.Y(n_15431)
);

AND2x4_ASAP7_75t_L g15432 ( 
.A(n_14319),
.B(n_14251),
.Y(n_15432)
);

AO21x2_ASAP7_75t_L g15433 ( 
.A1(n_14347),
.A2(n_13975),
.B(n_13886),
.Y(n_15433)
);

NOR2x1p5_ASAP7_75t_L g15434 ( 
.A(n_14604),
.B(n_13502),
.Y(n_15434)
);

OR2x2_ASAP7_75t_L g15435 ( 
.A(n_15124),
.B(n_14109),
.Y(n_15435)
);

BUFx3_ASAP7_75t_L g15436 ( 
.A(n_14827),
.Y(n_15436)
);

AND2x2_ASAP7_75t_L g15437 ( 
.A(n_14851),
.B(n_14479),
.Y(n_15437)
);

INVxp67_ASAP7_75t_SL g15438 ( 
.A(n_14538),
.Y(n_15438)
);

INVx1_ASAP7_75t_L g15439 ( 
.A(n_14883),
.Y(n_15439)
);

AOI22xp33_ASAP7_75t_L g15440 ( 
.A1(n_14526),
.A2(n_14097),
.B1(n_14195),
.B2(n_13992),
.Y(n_15440)
);

INVx1_ASAP7_75t_L g15441 ( 
.A(n_14889),
.Y(n_15441)
);

INVxp67_ASAP7_75t_L g15442 ( 
.A(n_14904),
.Y(n_15442)
);

BUFx2_ASAP7_75t_L g15443 ( 
.A(n_14319),
.Y(n_15443)
);

AND2x2_ASAP7_75t_L g15444 ( 
.A(n_14839),
.B(n_14228),
.Y(n_15444)
);

AND2x2_ASAP7_75t_L g15445 ( 
.A(n_14842),
.B(n_14233),
.Y(n_15445)
);

AO21x2_ASAP7_75t_L g15446 ( 
.A1(n_14363),
.A2(n_13445),
.B(n_13864),
.Y(n_15446)
);

INVx1_ASAP7_75t_L g15447 ( 
.A(n_14929),
.Y(n_15447)
);

HB1xp67_ASAP7_75t_L g15448 ( 
.A(n_14618),
.Y(n_15448)
);

AND2x2_ASAP7_75t_L g15449 ( 
.A(n_14643),
.B(n_14151),
.Y(n_15449)
);

AND2x2_ASAP7_75t_L g15450 ( 
.A(n_14354),
.B(n_14583),
.Y(n_15450)
);

INVx1_ASAP7_75t_L g15451 ( 
.A(n_14722),
.Y(n_15451)
);

OR2x2_ASAP7_75t_L g15452 ( 
.A(n_15047),
.B(n_14149),
.Y(n_15452)
);

AND2x4_ASAP7_75t_L g15453 ( 
.A(n_14837),
.B(n_14241),
.Y(n_15453)
);

INVx2_ASAP7_75t_L g15454 ( 
.A(n_14491),
.Y(n_15454)
);

INVx2_ASAP7_75t_L g15455 ( 
.A(n_14497),
.Y(n_15455)
);

BUFx6f_ASAP7_75t_L g15456 ( 
.A(n_14759),
.Y(n_15456)
);

AND2x2_ASAP7_75t_L g15457 ( 
.A(n_14917),
.B(n_14127),
.Y(n_15457)
);

NAND2xp5_ASAP7_75t_L g15458 ( 
.A(n_14822),
.B(n_13986),
.Y(n_15458)
);

INVx1_ASAP7_75t_L g15459 ( 
.A(n_14709),
.Y(n_15459)
);

INVx1_ASAP7_75t_L g15460 ( 
.A(n_14875),
.Y(n_15460)
);

NAND2xp5_ASAP7_75t_L g15461 ( 
.A(n_14841),
.B(n_13986),
.Y(n_15461)
);

INVx1_ASAP7_75t_L g15462 ( 
.A(n_14949),
.Y(n_15462)
);

INVx2_ASAP7_75t_SL g15463 ( 
.A(n_14661),
.Y(n_15463)
);

INVx2_ASAP7_75t_L g15464 ( 
.A(n_14499),
.Y(n_15464)
);

BUFx3_ASAP7_75t_L g15465 ( 
.A(n_14836),
.Y(n_15465)
);

AOI222xp33_ASAP7_75t_L g15466 ( 
.A1(n_14414),
.A2(n_14159),
.B1(n_14157),
.B2(n_14208),
.C1(n_14070),
.C2(n_14049),
.Y(n_15466)
);

HB1xp67_ASAP7_75t_L g15467 ( 
.A(n_14923),
.Y(n_15467)
);

INVx1_ASAP7_75t_L g15468 ( 
.A(n_14952),
.Y(n_15468)
);

INVxp67_ASAP7_75t_L g15469 ( 
.A(n_14927),
.Y(n_15469)
);

BUFx3_ASAP7_75t_L g15470 ( 
.A(n_14849),
.Y(n_15470)
);

INVx2_ASAP7_75t_L g15471 ( 
.A(n_14494),
.Y(n_15471)
);

AND2x2_ASAP7_75t_L g15472 ( 
.A(n_14888),
.B(n_14127),
.Y(n_15472)
);

AND2x2_ASAP7_75t_L g15473 ( 
.A(n_14890),
.B(n_14119),
.Y(n_15473)
);

AND2x2_ASAP7_75t_L g15474 ( 
.A(n_14896),
.B(n_14119),
.Y(n_15474)
);

AND2x2_ASAP7_75t_L g15475 ( 
.A(n_14920),
.B(n_14144),
.Y(n_15475)
);

AND2x2_ASAP7_75t_L g15476 ( 
.A(n_14661),
.B(n_14150),
.Y(n_15476)
);

INVx2_ASAP7_75t_L g15477 ( 
.A(n_14494),
.Y(n_15477)
);

NAND2xp5_ASAP7_75t_L g15478 ( 
.A(n_14932),
.B(n_13986),
.Y(n_15478)
);

OR2x2_ASAP7_75t_L g15479 ( 
.A(n_14694),
.B(n_14152),
.Y(n_15479)
);

HB1xp67_ASAP7_75t_L g15480 ( 
.A(n_14938),
.Y(n_15480)
);

AND2x2_ASAP7_75t_L g15481 ( 
.A(n_14702),
.B(n_14242),
.Y(n_15481)
);

NOR2xp67_ASAP7_75t_L g15482 ( 
.A(n_14777),
.B(n_14246),
.Y(n_15482)
);

INVx4_ASAP7_75t_L g15483 ( 
.A(n_14577),
.Y(n_15483)
);

BUFx3_ASAP7_75t_L g15484 ( 
.A(n_14580),
.Y(n_15484)
);

AND2x2_ASAP7_75t_L g15485 ( 
.A(n_14702),
.B(n_14217),
.Y(n_15485)
);

INVx1_ASAP7_75t_L g15486 ( 
.A(n_14974),
.Y(n_15486)
);

INVx2_ASAP7_75t_L g15487 ( 
.A(n_14532),
.Y(n_15487)
);

INVx2_ASAP7_75t_L g15488 ( 
.A(n_14532),
.Y(n_15488)
);

OAI22xp5_ASAP7_75t_L g15489 ( 
.A1(n_14707),
.A2(n_13457),
.B1(n_14295),
.B2(n_14087),
.Y(n_15489)
);

AND2x2_ASAP7_75t_L g15490 ( 
.A(n_14704),
.B(n_14710),
.Y(n_15490)
);

INVx1_ASAP7_75t_L g15491 ( 
.A(n_14620),
.Y(n_15491)
);

OR2x2_ASAP7_75t_L g15492 ( 
.A(n_14983),
.B(n_14163),
.Y(n_15492)
);

OR2x2_ASAP7_75t_L g15493 ( 
.A(n_14634),
.B(n_14185),
.Y(n_15493)
);

INVx3_ASAP7_75t_L g15494 ( 
.A(n_15032),
.Y(n_15494)
);

HB1xp67_ASAP7_75t_L g15495 ( 
.A(n_14954),
.Y(n_15495)
);

AOI22xp33_ASAP7_75t_L g15496 ( 
.A1(n_14539),
.A2(n_14253),
.B1(n_14061),
.B2(n_14074),
.Y(n_15496)
);

INVx2_ASAP7_75t_L g15497 ( 
.A(n_14630),
.Y(n_15497)
);

INVx2_ASAP7_75t_L g15498 ( 
.A(n_14733),
.Y(n_15498)
);

NAND2xp5_ASAP7_75t_L g15499 ( 
.A(n_14960),
.B(n_14075),
.Y(n_15499)
);

INVx1_ASAP7_75t_L g15500 ( 
.A(n_14668),
.Y(n_15500)
);

INVx1_ASAP7_75t_L g15501 ( 
.A(n_14675),
.Y(n_15501)
);

INVx1_ASAP7_75t_L g15502 ( 
.A(n_14315),
.Y(n_15502)
);

AND2x2_ASAP7_75t_L g15503 ( 
.A(n_14704),
.B(n_14212),
.Y(n_15503)
);

INVx1_ASAP7_75t_L g15504 ( 
.A(n_15045),
.Y(n_15504)
);

INVx2_ASAP7_75t_L g15505 ( 
.A(n_14733),
.Y(n_15505)
);

OR2x2_ASAP7_75t_L g15506 ( 
.A(n_14529),
.B(n_14232),
.Y(n_15506)
);

BUFx2_ASAP7_75t_L g15507 ( 
.A(n_14383),
.Y(n_15507)
);

HB1xp67_ASAP7_75t_L g15508 ( 
.A(n_14905),
.Y(n_15508)
);

INVx2_ASAP7_75t_L g15509 ( 
.A(n_14324),
.Y(n_15509)
);

INVx3_ASAP7_75t_L g15510 ( 
.A(n_15043),
.Y(n_15510)
);

INVx2_ASAP7_75t_L g15511 ( 
.A(n_14330),
.Y(n_15511)
);

BUFx6f_ASAP7_75t_L g15512 ( 
.A(n_14331),
.Y(n_15512)
);

INVxp67_ASAP7_75t_SL g15513 ( 
.A(n_14980),
.Y(n_15513)
);

INVx2_ASAP7_75t_L g15514 ( 
.A(n_14338),
.Y(n_15514)
);

INVx1_ASAP7_75t_L g15515 ( 
.A(n_14396),
.Y(n_15515)
);

AND2x2_ASAP7_75t_L g15516 ( 
.A(n_14710),
.B(n_14126),
.Y(n_15516)
);

NAND2xp5_ASAP7_75t_L g15517 ( 
.A(n_14886),
.B(n_14190),
.Y(n_15517)
);

HB1xp67_ASAP7_75t_L g15518 ( 
.A(n_14924),
.Y(n_15518)
);

BUFx2_ASAP7_75t_L g15519 ( 
.A(n_15075),
.Y(n_15519)
);

OR2x2_ASAP7_75t_L g15520 ( 
.A(n_14590),
.B(n_13467),
.Y(n_15520)
);

INVx1_ASAP7_75t_L g15521 ( 
.A(n_14399),
.Y(n_15521)
);

INVx1_ASAP7_75t_L g15522 ( 
.A(n_14409),
.Y(n_15522)
);

AND2x2_ASAP7_75t_L g15523 ( 
.A(n_14901),
.B(n_14133),
.Y(n_15523)
);

INVx3_ASAP7_75t_L g15524 ( 
.A(n_15043),
.Y(n_15524)
);

INVx4_ASAP7_75t_L g15525 ( 
.A(n_15075),
.Y(n_15525)
);

BUFx2_ASAP7_75t_L g15526 ( 
.A(n_14317),
.Y(n_15526)
);

INVx2_ASAP7_75t_SL g15527 ( 
.A(n_14464),
.Y(n_15527)
);

INVx2_ASAP7_75t_L g15528 ( 
.A(n_14345),
.Y(n_15528)
);

INVx2_ASAP7_75t_L g15529 ( 
.A(n_14353),
.Y(n_15529)
);

AND2x2_ASAP7_75t_L g15530 ( 
.A(n_14815),
.B(n_14138),
.Y(n_15530)
);

AND2x2_ASAP7_75t_L g15531 ( 
.A(n_14829),
.B(n_14141),
.Y(n_15531)
);

INVx1_ASAP7_75t_L g15532 ( 
.A(n_14410),
.Y(n_15532)
);

NAND2xp5_ASAP7_75t_L g15533 ( 
.A(n_15059),
.B(n_14171),
.Y(n_15533)
);

INVx1_ASAP7_75t_L g15534 ( 
.A(n_14425),
.Y(n_15534)
);

INVx1_ASAP7_75t_L g15535 ( 
.A(n_14426),
.Y(n_15535)
);

INVx2_ASAP7_75t_L g15536 ( 
.A(n_14356),
.Y(n_15536)
);

BUFx2_ASAP7_75t_L g15537 ( 
.A(n_15111),
.Y(n_15537)
);

INVx1_ASAP7_75t_L g15538 ( 
.A(n_14427),
.Y(n_15538)
);

INVx1_ASAP7_75t_L g15539 ( 
.A(n_14428),
.Y(n_15539)
);

INVx3_ASAP7_75t_L g15540 ( 
.A(n_15018),
.Y(n_15540)
);

INVx1_ASAP7_75t_L g15541 ( 
.A(n_14429),
.Y(n_15541)
);

INVxp67_ASAP7_75t_SL g15542 ( 
.A(n_14717),
.Y(n_15542)
);

INVx2_ASAP7_75t_L g15543 ( 
.A(n_14365),
.Y(n_15543)
);

AND2x2_ASAP7_75t_L g15544 ( 
.A(n_14718),
.B(n_14142),
.Y(n_15544)
);

INVx2_ASAP7_75t_L g15545 ( 
.A(n_14372),
.Y(n_15545)
);

AND2x2_ASAP7_75t_L g15546 ( 
.A(n_14718),
.B(n_14114),
.Y(n_15546)
);

AND2x2_ASAP7_75t_L g15547 ( 
.A(n_14859),
.B(n_14114),
.Y(n_15547)
);

INVx3_ASAP7_75t_L g15548 ( 
.A(n_15018),
.Y(n_15548)
);

INVx1_ASAP7_75t_L g15549 ( 
.A(n_14432),
.Y(n_15549)
);

HB1xp67_ASAP7_75t_L g15550 ( 
.A(n_14458),
.Y(n_15550)
);

OR2x2_ASAP7_75t_L g15551 ( 
.A(n_15061),
.B(n_13492),
.Y(n_15551)
);

AND2x2_ASAP7_75t_L g15552 ( 
.A(n_14864),
.B(n_14268),
.Y(n_15552)
);

HB1xp67_ASAP7_75t_L g15553 ( 
.A(n_14462),
.Y(n_15553)
);

INVx1_ASAP7_75t_L g15554 ( 
.A(n_14438),
.Y(n_15554)
);

INVx2_ASAP7_75t_L g15555 ( 
.A(n_14405),
.Y(n_15555)
);

AND2x4_ASAP7_75t_SL g15556 ( 
.A(n_14868),
.B(n_14392),
.Y(n_15556)
);

AND2x4_ASAP7_75t_L g15557 ( 
.A(n_15086),
.B(n_14887),
.Y(n_15557)
);

HB1xp67_ASAP7_75t_L g15558 ( 
.A(n_14467),
.Y(n_15558)
);

INVx1_ASAP7_75t_L g15559 ( 
.A(n_14440),
.Y(n_15559)
);

INVx3_ASAP7_75t_L g15560 ( 
.A(n_15008),
.Y(n_15560)
);

INVx2_ASAP7_75t_L g15561 ( 
.A(n_14415),
.Y(n_15561)
);

AND2x2_ASAP7_75t_L g15562 ( 
.A(n_14464),
.B(n_14259),
.Y(n_15562)
);

AO21x2_ASAP7_75t_L g15563 ( 
.A1(n_14910),
.A2(n_13684),
.B(n_14088),
.Y(n_15563)
);

AND2x2_ASAP7_75t_L g15564 ( 
.A(n_14967),
.B(n_14213),
.Y(n_15564)
);

NAND2xp5_ASAP7_75t_L g15565 ( 
.A(n_14918),
.B(n_14122),
.Y(n_15565)
);

AND2x4_ASAP7_75t_L g15566 ( 
.A(n_14401),
.B(n_14269),
.Y(n_15566)
);

INVxp33_ASAP7_75t_L g15567 ( 
.A(n_14421),
.Y(n_15567)
);

INVx1_ASAP7_75t_L g15568 ( 
.A(n_14445),
.Y(n_15568)
);

INVx1_ASAP7_75t_L g15569 ( 
.A(n_14446),
.Y(n_15569)
);

HB1xp67_ASAP7_75t_L g15570 ( 
.A(n_14468),
.Y(n_15570)
);

AND2x2_ASAP7_75t_L g15571 ( 
.A(n_14967),
.B(n_14222),
.Y(n_15571)
);

NAND2xp5_ASAP7_75t_L g15572 ( 
.A(n_14834),
.B(n_14026),
.Y(n_15572)
);

NAND2xp5_ASAP7_75t_L g15573 ( 
.A(n_14843),
.B(n_14030),
.Y(n_15573)
);

INVx2_ASAP7_75t_L g15574 ( 
.A(n_14420),
.Y(n_15574)
);

INVx1_ASAP7_75t_L g15575 ( 
.A(n_14451),
.Y(n_15575)
);

AND2x2_ASAP7_75t_L g15576 ( 
.A(n_15008),
.B(n_13545),
.Y(n_15576)
);

INVx2_ASAP7_75t_SL g15577 ( 
.A(n_14899),
.Y(n_15577)
);

INVx1_ASAP7_75t_L g15578 ( 
.A(n_14455),
.Y(n_15578)
);

AND2x2_ASAP7_75t_L g15579 ( 
.A(n_15009),
.B(n_14130),
.Y(n_15579)
);

INVx1_ASAP7_75t_L g15580 ( 
.A(n_14457),
.Y(n_15580)
);

INVx2_ASAP7_75t_L g15581 ( 
.A(n_14430),
.Y(n_15581)
);

INVxp67_ASAP7_75t_SL g15582 ( 
.A(n_14404),
.Y(n_15582)
);

NAND2xp5_ASAP7_75t_L g15583 ( 
.A(n_14852),
.B(n_14043),
.Y(n_15583)
);

INVx1_ASAP7_75t_L g15584 ( 
.A(n_14459),
.Y(n_15584)
);

OR2x2_ASAP7_75t_L g15585 ( 
.A(n_15042),
.B(n_14286),
.Y(n_15585)
);

INVx1_ASAP7_75t_L g15586 ( 
.A(n_14466),
.Y(n_15586)
);

NAND2xp5_ASAP7_75t_L g15587 ( 
.A(n_14854),
.B(n_14124),
.Y(n_15587)
);

NOR2xp33_ASAP7_75t_SL g15588 ( 
.A(n_14509),
.B(n_10486),
.Y(n_15588)
);

AND2x2_ASAP7_75t_L g15589 ( 
.A(n_15009),
.B(n_14130),
.Y(n_15589)
);

BUFx2_ASAP7_75t_L g15590 ( 
.A(n_14895),
.Y(n_15590)
);

INVx4_ASAP7_75t_L g15591 ( 
.A(n_14431),
.Y(n_15591)
);

INVx1_ASAP7_75t_L g15592 ( 
.A(n_14469),
.Y(n_15592)
);

INVx2_ASAP7_75t_SL g15593 ( 
.A(n_14998),
.Y(n_15593)
);

INVx3_ASAP7_75t_L g15594 ( 
.A(n_14848),
.Y(n_15594)
);

AND2x2_ASAP7_75t_L g15595 ( 
.A(n_14998),
.B(n_14276),
.Y(n_15595)
);

AND2x4_ASAP7_75t_L g15596 ( 
.A(n_14624),
.B(n_14269),
.Y(n_15596)
);

AOI21xp33_ASAP7_75t_L g15597 ( 
.A1(n_14542),
.A2(n_14186),
.B(n_14059),
.Y(n_15597)
);

INVx1_ASAP7_75t_L g15598 ( 
.A(n_14527),
.Y(n_15598)
);

AND2x2_ASAP7_75t_L g15599 ( 
.A(n_15004),
.B(n_14277),
.Y(n_15599)
);

INVx2_ASAP7_75t_L g15600 ( 
.A(n_14433),
.Y(n_15600)
);

AND2x2_ASAP7_75t_L g15601 ( 
.A(n_15004),
.B(n_14271),
.Y(n_15601)
);

HB1xp67_ASAP7_75t_L g15602 ( 
.A(n_14493),
.Y(n_15602)
);

INVx2_ASAP7_75t_L g15603 ( 
.A(n_15138),
.Y(n_15603)
);

INVx1_ASAP7_75t_L g15604 ( 
.A(n_14528),
.Y(n_15604)
);

INVx3_ASAP7_75t_L g15605 ( 
.A(n_14848),
.Y(n_15605)
);

INVx2_ASAP7_75t_L g15606 ( 
.A(n_14682),
.Y(n_15606)
);

INVxp67_ASAP7_75t_L g15607 ( 
.A(n_14775),
.Y(n_15607)
);

INVx1_ASAP7_75t_L g15608 ( 
.A(n_14500),
.Y(n_15608)
);

AO21x2_ASAP7_75t_L g15609 ( 
.A1(n_14749),
.A2(n_14058),
.B(n_14055),
.Y(n_15609)
);

OR2x2_ASAP7_75t_L g15610 ( 
.A(n_15084),
.B(n_14008),
.Y(n_15610)
);

AND2x2_ASAP7_75t_L g15611 ( 
.A(n_14655),
.B(n_14297),
.Y(n_15611)
);

AND2x2_ASAP7_75t_L g15612 ( 
.A(n_14867),
.B(n_13919),
.Y(n_15612)
);

NOR2x1_ASAP7_75t_SL g15613 ( 
.A(n_14496),
.B(n_13736),
.Y(n_15613)
);

INVx1_ASAP7_75t_L g15614 ( 
.A(n_14811),
.Y(n_15614)
);

INVx1_ASAP7_75t_L g15615 ( 
.A(n_14818),
.Y(n_15615)
);

INVx2_ASAP7_75t_L g15616 ( 
.A(n_15112),
.Y(n_15616)
);

INVx2_ASAP7_75t_L g15617 ( 
.A(n_14720),
.Y(n_15617)
);

INVx2_ASAP7_75t_L g15618 ( 
.A(n_14595),
.Y(n_15618)
);

NAND2xp5_ASAP7_75t_L g15619 ( 
.A(n_14855),
.B(n_14140),
.Y(n_15619)
);

AND2x2_ASAP7_75t_L g15620 ( 
.A(n_14867),
.B(n_13921),
.Y(n_15620)
);

INVx2_ASAP7_75t_L g15621 ( 
.A(n_14559),
.Y(n_15621)
);

NAND2xp5_ASAP7_75t_L g15622 ( 
.A(n_14861),
.B(n_14262),
.Y(n_15622)
);

AND2x2_ASAP7_75t_L g15623 ( 
.A(n_14913),
.B(n_14946),
.Y(n_15623)
);

INVx1_ASAP7_75t_L g15624 ( 
.A(n_14830),
.Y(n_15624)
);

AND2x2_ASAP7_75t_L g15625 ( 
.A(n_14913),
.B(n_13922),
.Y(n_15625)
);

INVxp67_ASAP7_75t_SL g15626 ( 
.A(n_14435),
.Y(n_15626)
);

OR2x6_ASAP7_75t_L g15627 ( 
.A(n_14706),
.B(n_14188),
.Y(n_15627)
);

INVx1_ASAP7_75t_L g15628 ( 
.A(n_14866),
.Y(n_15628)
);

AND2x2_ASAP7_75t_L g15629 ( 
.A(n_14946),
.B(n_13995),
.Y(n_15629)
);

HB1xp67_ASAP7_75t_L g15630 ( 
.A(n_14627),
.Y(n_15630)
);

INVx2_ASAP7_75t_L g15631 ( 
.A(n_14562),
.Y(n_15631)
);

INVx1_ASAP7_75t_L g15632 ( 
.A(n_14880),
.Y(n_15632)
);

AND2x4_ASAP7_75t_L g15633 ( 
.A(n_14642),
.B(n_14234),
.Y(n_15633)
);

NAND2xp5_ASAP7_75t_L g15634 ( 
.A(n_14862),
.B(n_14281),
.Y(n_15634)
);

NAND2xp5_ASAP7_75t_L g15635 ( 
.A(n_14869),
.B(n_14257),
.Y(n_15635)
);

INVx2_ASAP7_75t_L g15636 ( 
.A(n_14564),
.Y(n_15636)
);

INVx2_ASAP7_75t_R g15637 ( 
.A(n_14318),
.Y(n_15637)
);

AND2x4_ASAP7_75t_L g15638 ( 
.A(n_14647),
.B(n_14246),
.Y(n_15638)
);

INVx2_ASAP7_75t_L g15639 ( 
.A(n_15048),
.Y(n_15639)
);

AND2x2_ASAP7_75t_L g15640 ( 
.A(n_14953),
.B(n_14966),
.Y(n_15640)
);

INVxp67_ASAP7_75t_SL g15641 ( 
.A(n_14516),
.Y(n_15641)
);

HB1xp67_ASAP7_75t_L g15642 ( 
.A(n_14656),
.Y(n_15642)
);

INVx1_ASAP7_75t_L g15643 ( 
.A(n_14700),
.Y(n_15643)
);

OAI322xp33_ASAP7_75t_L g15644 ( 
.A1(n_14321),
.A2(n_14128),
.A3(n_14060),
.B1(n_14064),
.B2(n_13601),
.C1(n_13580),
.C2(n_13598),
.Y(n_15644)
);

INVx1_ASAP7_75t_L g15645 ( 
.A(n_14703),
.Y(n_15645)
);

INVx1_ASAP7_75t_L g15646 ( 
.A(n_14705),
.Y(n_15646)
);

AND2x2_ASAP7_75t_L g15647 ( 
.A(n_14953),
.B(n_14270),
.Y(n_15647)
);

OR2x2_ASAP7_75t_L g15648 ( 
.A(n_14550),
.B(n_13957),
.Y(n_15648)
);

INVx3_ASAP7_75t_L g15649 ( 
.A(n_14966),
.Y(n_15649)
);

AND2x2_ASAP7_75t_L g15650 ( 
.A(n_15118),
.B(n_14263),
.Y(n_15650)
);

INVx1_ASAP7_75t_L g15651 ( 
.A(n_14725),
.Y(n_15651)
);

BUFx2_ASAP7_75t_L g15652 ( 
.A(n_14443),
.Y(n_15652)
);

AO21x2_ASAP7_75t_L g15653 ( 
.A1(n_14540),
.A2(n_14090),
.B(n_14081),
.Y(n_15653)
);

INVx2_ASAP7_75t_L g15654 ( 
.A(n_15057),
.Y(n_15654)
);

HB1xp67_ASAP7_75t_L g15655 ( 
.A(n_14659),
.Y(n_15655)
);

INVx5_ASAP7_75t_SL g15656 ( 
.A(n_14667),
.Y(n_15656)
);

AOI22xp33_ASAP7_75t_L g15657 ( 
.A1(n_14541),
.A2(n_14010),
.B1(n_14091),
.B2(n_14089),
.Y(n_15657)
);

INVx2_ASAP7_75t_L g15658 ( 
.A(n_15065),
.Y(n_15658)
);

AND2x4_ASAP7_75t_L g15659 ( 
.A(n_14673),
.B(n_14252),
.Y(n_15659)
);

INVx1_ASAP7_75t_L g15660 ( 
.A(n_14769),
.Y(n_15660)
);

NOR2x1p5_ASAP7_75t_L g15661 ( 
.A(n_14665),
.B(n_14252),
.Y(n_15661)
);

OR2x6_ASAP7_75t_L g15662 ( 
.A(n_14736),
.B(n_14737),
.Y(n_15662)
);

NAND2xp5_ASAP7_75t_SL g15663 ( 
.A(n_14654),
.B(n_14295),
.Y(n_15663)
);

INVx2_ASAP7_75t_L g15664 ( 
.A(n_15072),
.Y(n_15664)
);

NAND2xp5_ASAP7_75t_L g15665 ( 
.A(n_14876),
.B(n_14205),
.Y(n_15665)
);

INVx3_ASAP7_75t_L g15666 ( 
.A(n_14771),
.Y(n_15666)
);

AND2x2_ASAP7_75t_L g15667 ( 
.A(n_14907),
.B(n_14037),
.Y(n_15667)
);

BUFx3_ASAP7_75t_L g15668 ( 
.A(n_14381),
.Y(n_15668)
);

INVx1_ASAP7_75t_L g15669 ( 
.A(n_14320),
.Y(n_15669)
);

INVx1_ASAP7_75t_L g15670 ( 
.A(n_14325),
.Y(n_15670)
);

INVx3_ASAP7_75t_L g15671 ( 
.A(n_14771),
.Y(n_15671)
);

INVx1_ASAP7_75t_L g15672 ( 
.A(n_14332),
.Y(n_15672)
);

HB1xp67_ASAP7_75t_L g15673 ( 
.A(n_15055),
.Y(n_15673)
);

INVx2_ASAP7_75t_L g15674 ( 
.A(n_15082),
.Y(n_15674)
);

AND2x2_ASAP7_75t_L g15675 ( 
.A(n_14911),
.B(n_14065),
.Y(n_15675)
);

INVx2_ASAP7_75t_L g15676 ( 
.A(n_15085),
.Y(n_15676)
);

INVx1_ASAP7_75t_L g15677 ( 
.A(n_14334),
.Y(n_15677)
);

INVx1_ASAP7_75t_L g15678 ( 
.A(n_14335),
.Y(n_15678)
);

AND2x2_ASAP7_75t_L g15679 ( 
.A(n_14915),
.B(n_14068),
.Y(n_15679)
);

AND2x2_ASAP7_75t_L g15680 ( 
.A(n_14916),
.B(n_14076),
.Y(n_15680)
);

INVx1_ASAP7_75t_L g15681 ( 
.A(n_14336),
.Y(n_15681)
);

BUFx3_ASAP7_75t_L g15682 ( 
.A(n_14739),
.Y(n_15682)
);

INVx3_ASAP7_75t_L g15683 ( 
.A(n_14803),
.Y(n_15683)
);

AND2x2_ASAP7_75t_L g15684 ( 
.A(n_15132),
.B(n_14261),
.Y(n_15684)
);

INVx2_ASAP7_75t_L g15685 ( 
.A(n_15088),
.Y(n_15685)
);

OR2x2_ASAP7_75t_L g15686 ( 
.A(n_15031),
.B(n_14016),
.Y(n_15686)
);

INVx2_ASAP7_75t_L g15687 ( 
.A(n_15090),
.Y(n_15687)
);

NOR2x1_ASAP7_75t_SL g15688 ( 
.A(n_14969),
.B(n_10602),
.Y(n_15688)
);

AND2x2_ASAP7_75t_L g15689 ( 
.A(n_14817),
.B(n_14261),
.Y(n_15689)
);

HB1xp67_ASAP7_75t_L g15690 ( 
.A(n_15062),
.Y(n_15690)
);

NOR2xp33_ASAP7_75t_SL g15691 ( 
.A(n_14616),
.B(n_10602),
.Y(n_15691)
);

AND2x2_ASAP7_75t_L g15692 ( 
.A(n_14804),
.B(n_13893),
.Y(n_15692)
);

AND2x2_ASAP7_75t_L g15693 ( 
.A(n_14600),
.B(n_13903),
.Y(n_15693)
);

INVx3_ASAP7_75t_L g15694 ( 
.A(n_14803),
.Y(n_15694)
);

INVx1_ASAP7_75t_L g15695 ( 
.A(n_14339),
.Y(n_15695)
);

INVx1_ASAP7_75t_SL g15696 ( 
.A(n_14513),
.Y(n_15696)
);

AND2x2_ASAP7_75t_L g15697 ( 
.A(n_14602),
.B(n_13874),
.Y(n_15697)
);

AND2x2_ASAP7_75t_L g15698 ( 
.A(n_14603),
.B(n_14288),
.Y(n_15698)
);

INVx2_ASAP7_75t_L g15699 ( 
.A(n_15104),
.Y(n_15699)
);

AO21x2_ASAP7_75t_L g15700 ( 
.A1(n_14701),
.A2(n_14079),
.B(n_13552),
.Y(n_15700)
);

INVx2_ASAP7_75t_L g15701 ( 
.A(n_14768),
.Y(n_15701)
);

INVx1_ASAP7_75t_L g15702 ( 
.A(n_14352),
.Y(n_15702)
);

AND2x2_ASAP7_75t_L g15703 ( 
.A(n_14605),
.B(n_14051),
.Y(n_15703)
);

INVx2_ASAP7_75t_L g15704 ( 
.A(n_14713),
.Y(n_15704)
);

INVx2_ASAP7_75t_L g15705 ( 
.A(n_15122),
.Y(n_15705)
);

AND2x2_ASAP7_75t_L g15706 ( 
.A(n_14622),
.B(n_14051),
.Y(n_15706)
);

AOI221xp5_ASAP7_75t_L g15707 ( 
.A1(n_14460),
.A2(n_14052),
.B1(n_14089),
.B2(n_14091),
.C(n_13778),
.Y(n_15707)
);

INVx1_ASAP7_75t_L g15708 ( 
.A(n_14358),
.Y(n_15708)
);

AND2x2_ASAP7_75t_L g15709 ( 
.A(n_15017),
.B(n_13647),
.Y(n_15709)
);

INVx1_ASAP7_75t_L g15710 ( 
.A(n_15060),
.Y(n_15710)
);

INVx4_ASAP7_75t_L g15711 ( 
.A(n_14751),
.Y(n_15711)
);

AND2x2_ASAP7_75t_L g15712 ( 
.A(n_14687),
.B(n_14274),
.Y(n_15712)
);

BUFx3_ASAP7_75t_L g15713 ( 
.A(n_14878),
.Y(n_15713)
);

INVx2_ASAP7_75t_SL g15714 ( 
.A(n_15013),
.Y(n_15714)
);

AND2x2_ASAP7_75t_L g15715 ( 
.A(n_14690),
.B(n_14274),
.Y(n_15715)
);

AND2x4_ASAP7_75t_L g15716 ( 
.A(n_14881),
.B(n_10396),
.Y(n_15716)
);

OR2x2_ASAP7_75t_L g15717 ( 
.A(n_15126),
.B(n_14023),
.Y(n_15717)
);

INVx1_ASAP7_75t_L g15718 ( 
.A(n_15063),
.Y(n_15718)
);

OR2x2_ASAP7_75t_L g15719 ( 
.A(n_14520),
.B(n_14029),
.Y(n_15719)
);

INVx1_ASAP7_75t_L g15720 ( 
.A(n_15064),
.Y(n_15720)
);

CKINVDCx16_ASAP7_75t_R g15721 ( 
.A(n_14628),
.Y(n_15721)
);

OR2x2_ASAP7_75t_L g15722 ( 
.A(n_14524),
.B(n_14034),
.Y(n_15722)
);

OR2x2_ASAP7_75t_L g15723 ( 
.A(n_15056),
.B(n_14547),
.Y(n_15723)
);

OR2x2_ASAP7_75t_L g15724 ( 
.A(n_14377),
.B(n_13896),
.Y(n_15724)
);

INVx3_ASAP7_75t_L g15725 ( 
.A(n_14742),
.Y(n_15725)
);

OR2x2_ASAP7_75t_L g15726 ( 
.A(n_14484),
.B(n_13914),
.Y(n_15726)
);

AND2x2_ASAP7_75t_L g15727 ( 
.A(n_14708),
.B(n_13851),
.Y(n_15727)
);

INVxp67_ASAP7_75t_SL g15728 ( 
.A(n_14779),
.Y(n_15728)
);

BUFx2_ASAP7_75t_L g15729 ( 
.A(n_14386),
.Y(n_15729)
);

INVx1_ASAP7_75t_L g15730 ( 
.A(n_15068),
.Y(n_15730)
);

AND2x2_ASAP7_75t_L g15731 ( 
.A(n_14760),
.B(n_13866),
.Y(n_15731)
);

INVx2_ASAP7_75t_L g15732 ( 
.A(n_15125),
.Y(n_15732)
);

AND2x4_ASAP7_75t_L g15733 ( 
.A(n_14882),
.B(n_10396),
.Y(n_15733)
);

INVx1_ASAP7_75t_L g15734 ( 
.A(n_15069),
.Y(n_15734)
);

AND2x2_ASAP7_75t_SL g15735 ( 
.A(n_14355),
.B(n_14348),
.Y(n_15735)
);

AND2x2_ASAP7_75t_L g15736 ( 
.A(n_14664),
.B(n_13875),
.Y(n_15736)
);

INVx1_ASAP7_75t_L g15737 ( 
.A(n_15070),
.Y(n_15737)
);

NAND2xp5_ASAP7_75t_L g15738 ( 
.A(n_14903),
.B(n_14104),
.Y(n_15738)
);

AND2x2_ASAP7_75t_L g15739 ( 
.A(n_14666),
.B(n_13839),
.Y(n_15739)
);

AND2x2_ASAP7_75t_L g15740 ( 
.A(n_14678),
.B(n_11774),
.Y(n_15740)
);

INVx1_ASAP7_75t_L g15741 ( 
.A(n_15074),
.Y(n_15741)
);

BUFx2_ASAP7_75t_L g15742 ( 
.A(n_14391),
.Y(n_15742)
);

AO21x2_ASAP7_75t_L g15743 ( 
.A1(n_15134),
.A2(n_14113),
.B(n_14103),
.Y(n_15743)
);

AND2x2_ASAP7_75t_L g15744 ( 
.A(n_14754),
.B(n_11776),
.Y(n_15744)
);

OR2x2_ASAP7_75t_L g15745 ( 
.A(n_14533),
.B(n_14104),
.Y(n_15745)
);

INVx2_ASAP7_75t_L g15746 ( 
.A(n_14801),
.Y(n_15746)
);

INVx1_ASAP7_75t_L g15747 ( 
.A(n_15080),
.Y(n_15747)
);

AND2x4_ASAP7_75t_L g15748 ( 
.A(n_14937),
.B(n_14940),
.Y(n_15748)
);

INVx3_ASAP7_75t_L g15749 ( 
.A(n_14648),
.Y(n_15749)
);

INVx2_ASAP7_75t_L g15750 ( 
.A(n_14807),
.Y(n_15750)
);

AND2x2_ASAP7_75t_L g15751 ( 
.A(n_14763),
.B(n_11780),
.Y(n_15751)
);

INVx1_ASAP7_75t_L g15752 ( 
.A(n_15081),
.Y(n_15752)
);

INVx2_ASAP7_75t_L g15753 ( 
.A(n_14809),
.Y(n_15753)
);

INVx1_ASAP7_75t_L g15754 ( 
.A(n_15083),
.Y(n_15754)
);

INVx2_ASAP7_75t_SL g15755 ( 
.A(n_15023),
.Y(n_15755)
);

AND2x4_ASAP7_75t_L g15756 ( 
.A(n_14959),
.B(n_10583),
.Y(n_15756)
);

INVx1_ASAP7_75t_L g15757 ( 
.A(n_14306),
.Y(n_15757)
);

INVx1_ASAP7_75t_SL g15758 ( 
.A(n_14384),
.Y(n_15758)
);

AND2x2_ASAP7_75t_L g15759 ( 
.A(n_14764),
.B(n_11785),
.Y(n_15759)
);

AND2x2_ASAP7_75t_L g15760 ( 
.A(n_14784),
.B(n_11787),
.Y(n_15760)
);

INVx3_ASAP7_75t_L g15761 ( 
.A(n_14653),
.Y(n_15761)
);

AND2x4_ASAP7_75t_SL g15762 ( 
.A(n_14789),
.B(n_8072),
.Y(n_15762)
);

INVxp67_ASAP7_75t_L g15763 ( 
.A(n_14402),
.Y(n_15763)
);

HB1xp67_ASAP7_75t_L g15764 ( 
.A(n_14988),
.Y(n_15764)
);

INVx1_ASAP7_75t_L g15765 ( 
.A(n_14313),
.Y(n_15765)
);

INVx2_ASAP7_75t_L g15766 ( 
.A(n_14812),
.Y(n_15766)
);

INVx2_ASAP7_75t_L g15767 ( 
.A(n_14816),
.Y(n_15767)
);

OR2x2_ASAP7_75t_L g15768 ( 
.A(n_14537),
.B(n_14115),
.Y(n_15768)
);

NOR2x1_ASAP7_75t_SL g15769 ( 
.A(n_14632),
.B(n_10602),
.Y(n_15769)
);

INVx2_ASAP7_75t_L g15770 ( 
.A(n_14584),
.Y(n_15770)
);

AND2x4_ASAP7_75t_L g15771 ( 
.A(n_14545),
.B(n_10583),
.Y(n_15771)
);

INVx1_ASAP7_75t_SL g15772 ( 
.A(n_14376),
.Y(n_15772)
);

INVx1_ASAP7_75t_L g15773 ( 
.A(n_14548),
.Y(n_15773)
);

OR2x2_ASAP7_75t_L g15774 ( 
.A(n_14898),
.B(n_14115),
.Y(n_15774)
);

AND2x4_ASAP7_75t_L g15775 ( 
.A(n_14810),
.B(n_10583),
.Y(n_15775)
);

OAI22xp5_ASAP7_75t_L g15776 ( 
.A1(n_14503),
.A2(n_14279),
.B1(n_10622),
.B2(n_8728),
.Y(n_15776)
);

AOI22xp33_ASAP7_75t_L g15777 ( 
.A1(n_14369),
.A2(n_11448),
.B1(n_11455),
.B2(n_11451),
.Y(n_15777)
);

INVx4_ASAP7_75t_L g15778 ( 
.A(n_14814),
.Y(n_15778)
);

AND2x2_ASAP7_75t_L g15779 ( 
.A(n_15137),
.B(n_11792),
.Y(n_15779)
);

INVx1_ASAP7_75t_L g15780 ( 
.A(n_14558),
.Y(n_15780)
);

AND2x2_ASAP7_75t_L g15781 ( 
.A(n_14681),
.B(n_11793),
.Y(n_15781)
);

NOR2x1_ASAP7_75t_SL g15782 ( 
.A(n_14448),
.B(n_10613),
.Y(n_15782)
);

BUFx2_ASAP7_75t_L g15783 ( 
.A(n_14416),
.Y(n_15783)
);

INVx2_ASAP7_75t_SL g15784 ( 
.A(n_15024),
.Y(n_15784)
);

AND2x2_ASAP7_75t_L g15785 ( 
.A(n_15093),
.B(n_11795),
.Y(n_15785)
);

BUFx2_ASAP7_75t_L g15786 ( 
.A(n_14450),
.Y(n_15786)
);

INVx2_ASAP7_75t_SL g15787 ( 
.A(n_14506),
.Y(n_15787)
);

OR2x6_ASAP7_75t_SL g15788 ( 
.A(n_14657),
.B(n_13977),
.Y(n_15788)
);

HB1xp67_ASAP7_75t_L g15789 ( 
.A(n_14997),
.Y(n_15789)
);

INVx1_ASAP7_75t_L g15790 ( 
.A(n_14567),
.Y(n_15790)
);

INVx2_ASAP7_75t_L g15791 ( 
.A(n_14588),
.Y(n_15791)
);

INVx2_ASAP7_75t_L g15792 ( 
.A(n_14743),
.Y(n_15792)
);

AOI22xp33_ASAP7_75t_L g15793 ( 
.A1(n_14357),
.A2(n_11448),
.B1(n_11478),
.B2(n_11466),
.Y(n_15793)
);

INVx1_ASAP7_75t_L g15794 ( 
.A(n_14570),
.Y(n_15794)
);

INVx1_ASAP7_75t_L g15795 ( 
.A(n_14573),
.Y(n_15795)
);

INVx2_ASAP7_75t_L g15796 ( 
.A(n_14744),
.Y(n_15796)
);

OR2x2_ASAP7_75t_L g15797 ( 
.A(n_14398),
.B(n_14239),
.Y(n_15797)
);

AND2x2_ASAP7_75t_L g15798 ( 
.A(n_15094),
.B(n_11799),
.Y(n_15798)
);

BUFx2_ASAP7_75t_L g15799 ( 
.A(n_14579),
.Y(n_15799)
);

INVx1_ASAP7_75t_L g15800 ( 
.A(n_14609),
.Y(n_15800)
);

NOR2xp33_ASAP7_75t_L g15801 ( 
.A(n_14770),
.B(n_14790),
.Y(n_15801)
);

NOR2xp33_ASAP7_75t_L g15802 ( 
.A(n_15025),
.B(n_15027),
.Y(n_15802)
);

INVx2_ASAP7_75t_L g15803 ( 
.A(n_14594),
.Y(n_15803)
);

AND2x2_ASAP7_75t_L g15804 ( 
.A(n_14574),
.B(n_11812),
.Y(n_15804)
);

AND2x2_ASAP7_75t_L g15805 ( 
.A(n_14578),
.B(n_11820),
.Y(n_15805)
);

AND2x2_ASAP7_75t_L g15806 ( 
.A(n_14798),
.B(n_11821),
.Y(n_15806)
);

INVx2_ASAP7_75t_L g15807 ( 
.A(n_14729),
.Y(n_15807)
);

INVx1_ASAP7_75t_L g15808 ( 
.A(n_14611),
.Y(n_15808)
);

NOR3xp33_ASAP7_75t_L g15809 ( 
.A(n_15014),
.B(n_13316),
.C(n_13261),
.Y(n_15809)
);

HB1xp67_ASAP7_75t_L g15810 ( 
.A(n_15006),
.Y(n_15810)
);

INVx2_ASAP7_75t_L g15811 ( 
.A(n_15036),
.Y(n_15811)
);

INVx4_ASAP7_75t_L g15812 ( 
.A(n_14481),
.Y(n_15812)
);

INVx1_ASAP7_75t_L g15813 ( 
.A(n_15051),
.Y(n_15813)
);

NAND2xp5_ASAP7_75t_L g15814 ( 
.A(n_15028),
.B(n_14239),
.Y(n_15814)
);

INVx1_ASAP7_75t_L g15815 ( 
.A(n_14928),
.Y(n_15815)
);

INVx1_ASAP7_75t_L g15816 ( 
.A(n_14795),
.Y(n_15816)
);

AND2x2_ASAP7_75t_L g15817 ( 
.A(n_15041),
.B(n_11827),
.Y(n_15817)
);

AND2x2_ASAP7_75t_L g15818 ( 
.A(n_14596),
.B(n_11828),
.Y(n_15818)
);

INVx1_ASAP7_75t_L g15819 ( 
.A(n_14897),
.Y(n_15819)
);

INVx1_ASAP7_75t_L g15820 ( 
.A(n_14761),
.Y(n_15820)
);

INVxp67_ASAP7_75t_L g15821 ( 
.A(n_14470),
.Y(n_15821)
);

INVx1_ASAP7_75t_L g15822 ( 
.A(n_14778),
.Y(n_15822)
);

INVx2_ASAP7_75t_L g15823 ( 
.A(n_14957),
.Y(n_15823)
);

AOI22xp33_ASAP7_75t_L g15824 ( 
.A1(n_14303),
.A2(n_11466),
.B1(n_11479),
.B2(n_11478),
.Y(n_15824)
);

AND2x2_ASAP7_75t_L g15825 ( 
.A(n_14780),
.B(n_11834),
.Y(n_15825)
);

INVx1_ASAP7_75t_SL g15826 ( 
.A(n_15078),
.Y(n_15826)
);

AND2x2_ASAP7_75t_L g15827 ( 
.A(n_14787),
.B(n_11835),
.Y(n_15827)
);

INVx1_ASAP7_75t_L g15828 ( 
.A(n_14782),
.Y(n_15828)
);

INVx1_ASAP7_75t_L g15829 ( 
.A(n_14786),
.Y(n_15829)
);

NAND2xp5_ASAP7_75t_L g15830 ( 
.A(n_14941),
.B(n_14239),
.Y(n_15830)
);

OR2x2_ASAP7_75t_L g15831 ( 
.A(n_14726),
.B(n_11840),
.Y(n_15831)
);

INVxp67_ASAP7_75t_SL g15832 ( 
.A(n_14679),
.Y(n_15832)
);

INVx3_ASAP7_75t_L g15833 ( 
.A(n_14791),
.Y(n_15833)
);

AND2x2_ASAP7_75t_L g15834 ( 
.A(n_14546),
.B(n_11850),
.Y(n_15834)
);

AOI22xp33_ASAP7_75t_L g15835 ( 
.A1(n_14598),
.A2(n_11479),
.B1(n_11494),
.B2(n_11489),
.Y(n_15835)
);

AND2x2_ASAP7_75t_L g15836 ( 
.A(n_14961),
.B(n_11855),
.Y(n_15836)
);

NAND2xp5_ASAP7_75t_L g15837 ( 
.A(n_14942),
.B(n_8313),
.Y(n_15837)
);

AND2x2_ASAP7_75t_L g15838 ( 
.A(n_14989),
.B(n_11859),
.Y(n_15838)
);

INVx2_ASAP7_75t_L g15839 ( 
.A(n_14958),
.Y(n_15839)
);

INVxp67_ASAP7_75t_SL g15840 ( 
.A(n_14732),
.Y(n_15840)
);

INVx2_ASAP7_75t_L g15841 ( 
.A(n_14757),
.Y(n_15841)
);

INVx2_ASAP7_75t_L g15842 ( 
.A(n_15076),
.Y(n_15842)
);

INVx2_ASAP7_75t_L g15843 ( 
.A(n_15079),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_14993),
.B(n_11864),
.Y(n_15844)
);

AND2x2_ASAP7_75t_L g15845 ( 
.A(n_14995),
.B(n_11872),
.Y(n_15845)
);

INVx2_ASAP7_75t_L g15846 ( 
.A(n_15091),
.Y(n_15846)
);

INVx1_ASAP7_75t_L g15847 ( 
.A(n_14788),
.Y(n_15847)
);

AND2x2_ASAP7_75t_L g15848 ( 
.A(n_14483),
.B(n_11875),
.Y(n_15848)
);

INVx1_ASAP7_75t_L g15849 ( 
.A(n_14793),
.Y(n_15849)
);

AND2x2_ASAP7_75t_L g15850 ( 
.A(n_14490),
.B(n_14971),
.Y(n_15850)
);

INVx1_ASAP7_75t_L g15851 ( 
.A(n_14794),
.Y(n_15851)
);

AOI22xp33_ASAP7_75t_L g15852 ( 
.A1(n_14397),
.A2(n_11489),
.B1(n_11495),
.B2(n_11494),
.Y(n_15852)
);

OR2x2_ASAP7_75t_L g15853 ( 
.A(n_14762),
.B(n_11876),
.Y(n_15853)
);

OAI21xp5_ASAP7_75t_L g15854 ( 
.A1(n_14452),
.A2(n_11741),
.B(n_11740),
.Y(n_15854)
);

INVx2_ASAP7_75t_L g15855 ( 
.A(n_15096),
.Y(n_15855)
);

HB1xp67_ASAP7_75t_L g15856 ( 
.A(n_15116),
.Y(n_15856)
);

AND2x2_ASAP7_75t_L g15857 ( 
.A(n_14973),
.B(n_11878),
.Y(n_15857)
);

OR2x2_ASAP7_75t_L g15858 ( 
.A(n_15131),
.B(n_11881),
.Y(n_15858)
);

AND2x4_ASAP7_75t_SL g15859 ( 
.A(n_14651),
.B(n_8072),
.Y(n_15859)
);

INVx5_ASAP7_75t_SL g15860 ( 
.A(n_15120),
.Y(n_15860)
);

OR2x2_ASAP7_75t_L g15861 ( 
.A(n_14979),
.B(n_11888),
.Y(n_15861)
);

INVx1_ASAP7_75t_L g15862 ( 
.A(n_14797),
.Y(n_15862)
);

INVx4_ASAP7_75t_L g15863 ( 
.A(n_15135),
.Y(n_15863)
);

AND2x2_ASAP7_75t_L g15864 ( 
.A(n_14964),
.B(n_11895),
.Y(n_15864)
);

INVx1_ASAP7_75t_L g15865 ( 
.A(n_14800),
.Y(n_15865)
);

AND2x4_ASAP7_75t_L g15866 ( 
.A(n_14943),
.B(n_10583),
.Y(n_15866)
);

OAI22xp5_ASAP7_75t_L g15867 ( 
.A1(n_14337),
.A2(n_8775),
.B1(n_8579),
.B2(n_8401),
.Y(n_15867)
);

AND2x2_ASAP7_75t_L g15868 ( 
.A(n_14930),
.B(n_11901),
.Y(n_15868)
);

BUFx3_ASAP7_75t_L g15869 ( 
.A(n_14962),
.Y(n_15869)
);

AND2x2_ASAP7_75t_L g15870 ( 
.A(n_15139),
.B(n_14658),
.Y(n_15870)
);

INVx1_ASAP7_75t_L g15871 ( 
.A(n_15274),
.Y(n_15871)
);

AND2x4_ASAP7_75t_L g15872 ( 
.A(n_15268),
.B(n_14660),
.Y(n_15872)
);

OR2x2_ASAP7_75t_L g15873 ( 
.A(n_15319),
.B(n_14956),
.Y(n_15873)
);

OR2x2_ASAP7_75t_L g15874 ( 
.A(n_15186),
.B(n_15087),
.Y(n_15874)
);

INVx2_ASAP7_75t_L g15875 ( 
.A(n_15276),
.Y(n_15875)
);

OR2x2_ASAP7_75t_L g15876 ( 
.A(n_15154),
.B(n_15107),
.Y(n_15876)
);

NAND2xp5_ASAP7_75t_L g15877 ( 
.A(n_15141),
.B(n_15438),
.Y(n_15877)
);

NAND2xp5_ASAP7_75t_L g15878 ( 
.A(n_15204),
.B(n_14965),
.Y(n_15878)
);

AND2x4_ASAP7_75t_L g15879 ( 
.A(n_15431),
.B(n_15217),
.Y(n_15879)
);

INVx2_ASAP7_75t_SL g15880 ( 
.A(n_15173),
.Y(n_15880)
);

OA211x2_ASAP7_75t_L g15881 ( 
.A1(n_15588),
.A2(n_14870),
.B(n_14551),
.C(n_15097),
.Y(n_15881)
);

INVx1_ASAP7_75t_L g15882 ( 
.A(n_15219),
.Y(n_15882)
);

INVx2_ASAP7_75t_L g15883 ( 
.A(n_15519),
.Y(n_15883)
);

AND2x2_ASAP7_75t_L g15884 ( 
.A(n_15199),
.B(n_14662),
.Y(n_15884)
);

AND2x2_ASAP7_75t_L g15885 ( 
.A(n_15199),
.B(n_14669),
.Y(n_15885)
);

NAND2xp5_ASAP7_75t_L g15886 ( 
.A(n_15229),
.B(n_15175),
.Y(n_15886)
);

OR2x2_ASAP7_75t_L g15887 ( 
.A(n_15286),
.B(n_14805),
.Y(n_15887)
);

AND2x2_ASAP7_75t_L g15888 ( 
.A(n_15167),
.B(n_14671),
.Y(n_15888)
);

AND2x4_ASAP7_75t_L g15889 ( 
.A(n_15210),
.B(n_14676),
.Y(n_15889)
);

AND2x2_ASAP7_75t_L g15890 ( 
.A(n_15159),
.B(n_14677),
.Y(n_15890)
);

INVx1_ASAP7_75t_L g15891 ( 
.A(n_15219),
.Y(n_15891)
);

INVx1_ASAP7_75t_L g15892 ( 
.A(n_15367),
.Y(n_15892)
);

AND2x2_ASAP7_75t_L g15893 ( 
.A(n_15148),
.B(n_14680),
.Y(n_15893)
);

NAND2xp5_ASAP7_75t_L g15894 ( 
.A(n_15519),
.B(n_14970),
.Y(n_15894)
);

OR2x2_ASAP7_75t_L g15895 ( 
.A(n_15381),
.B(n_14808),
.Y(n_15895)
);

AND2x2_ASAP7_75t_L g15896 ( 
.A(n_15168),
.B(n_14683),
.Y(n_15896)
);

AND2x2_ASAP7_75t_L g15897 ( 
.A(n_15275),
.B(n_14686),
.Y(n_15897)
);

INVx1_ASAP7_75t_L g15898 ( 
.A(n_15467),
.Y(n_15898)
);

NOR2x1p5_ASAP7_75t_L g15899 ( 
.A(n_15241),
.B(n_14813),
.Y(n_15899)
);

AND2x2_ASAP7_75t_L g15900 ( 
.A(n_15212),
.B(n_14688),
.Y(n_15900)
);

AND2x2_ASAP7_75t_L g15901 ( 
.A(n_15262),
.B(n_14689),
.Y(n_15901)
);

NAND2xp5_ASAP7_75t_L g15902 ( 
.A(n_15200),
.B(n_14972),
.Y(n_15902)
);

AND2x2_ASAP7_75t_L g15903 ( 
.A(n_15142),
.B(n_14692),
.Y(n_15903)
);

AND2x2_ASAP7_75t_L g15904 ( 
.A(n_15145),
.B(n_14697),
.Y(n_15904)
);

INVx2_ASAP7_75t_L g15905 ( 
.A(n_15203),
.Y(n_15905)
);

INVx2_ASAP7_75t_L g15906 ( 
.A(n_15203),
.Y(n_15906)
);

AND2x2_ASAP7_75t_L g15907 ( 
.A(n_15231),
.B(n_14711),
.Y(n_15907)
);

OR2x2_ASAP7_75t_L g15908 ( 
.A(n_15180),
.B(n_15723),
.Y(n_15908)
);

AND2x2_ASAP7_75t_L g15909 ( 
.A(n_15184),
.B(n_14712),
.Y(n_15909)
);

AND2x2_ASAP7_75t_L g15910 ( 
.A(n_15194),
.B(n_14714),
.Y(n_15910)
);

NOR3xp33_ASAP7_75t_L g15911 ( 
.A(n_15322),
.B(n_15123),
.C(n_15095),
.Y(n_15911)
);

OR2x2_ASAP7_75t_L g15912 ( 
.A(n_15143),
.B(n_14820),
.Y(n_15912)
);

OR2x2_ASAP7_75t_L g15913 ( 
.A(n_15332),
.B(n_14821),
.Y(n_15913)
);

AND2x2_ASAP7_75t_L g15914 ( 
.A(n_15230),
.B(n_14715),
.Y(n_15914)
);

NAND2xp5_ASAP7_75t_L g15915 ( 
.A(n_15301),
.B(n_14975),
.Y(n_15915)
);

INVxp67_ASAP7_75t_SL g15916 ( 
.A(n_15297),
.Y(n_15916)
);

NAND2xp5_ASAP7_75t_L g15917 ( 
.A(n_15283),
.B(n_14976),
.Y(n_15917)
);

NAND2xp5_ASAP7_75t_L g15918 ( 
.A(n_15735),
.B(n_14982),
.Y(n_15918)
);

INVx1_ASAP7_75t_L g15919 ( 
.A(n_15480),
.Y(n_15919)
);

NAND2xp5_ASAP7_75t_L g15920 ( 
.A(n_15826),
.B(n_14986),
.Y(n_15920)
);

INVx1_ASAP7_75t_L g15921 ( 
.A(n_15495),
.Y(n_15921)
);

NAND2xp5_ASAP7_75t_L g15922 ( 
.A(n_15406),
.B(n_14990),
.Y(n_15922)
);

INVx1_ASAP7_75t_L g15923 ( 
.A(n_15266),
.Y(n_15923)
);

OR2x2_ASAP7_75t_L g15924 ( 
.A(n_15652),
.B(n_14824),
.Y(n_15924)
);

INVx1_ASAP7_75t_L g15925 ( 
.A(n_15272),
.Y(n_15925)
);

AND2x2_ASAP7_75t_L g15926 ( 
.A(n_15525),
.B(n_14716),
.Y(n_15926)
);

INVx4_ASAP7_75t_L g15927 ( 
.A(n_15173),
.Y(n_15927)
);

INVx1_ASAP7_75t_L g15928 ( 
.A(n_15161),
.Y(n_15928)
);

INVx1_ASAP7_75t_L g15929 ( 
.A(n_15161),
.Y(n_15929)
);

AND2x2_ASAP7_75t_L g15930 ( 
.A(n_15177),
.B(n_14719),
.Y(n_15930)
);

AND2x4_ASAP7_75t_L g15931 ( 
.A(n_15157),
.B(n_14723),
.Y(n_15931)
);

AND2x4_ASAP7_75t_L g15932 ( 
.A(n_15218),
.B(n_14728),
.Y(n_15932)
);

INVx1_ASAP7_75t_L g15933 ( 
.A(n_15376),
.Y(n_15933)
);

INVx4_ASAP7_75t_L g15934 ( 
.A(n_15173),
.Y(n_15934)
);

INVx1_ASAP7_75t_L g15935 ( 
.A(n_15376),
.Y(n_15935)
);

NOR2xp33_ASAP7_75t_SL g15936 ( 
.A(n_15320),
.B(n_10613),
.Y(n_15936)
);

NAND2xp5_ASAP7_75t_L g15937 ( 
.A(n_15406),
.B(n_14991),
.Y(n_15937)
);

AND2x2_ASAP7_75t_L g15938 ( 
.A(n_15472),
.B(n_14730),
.Y(n_15938)
);

NAND2xp5_ASAP7_75t_L g15939 ( 
.A(n_15537),
.B(n_14994),
.Y(n_15939)
);

INVx1_ASAP7_75t_L g15940 ( 
.A(n_15294),
.Y(n_15940)
);

NAND2xp5_ASAP7_75t_L g15941 ( 
.A(n_15537),
.B(n_14999),
.Y(n_15941)
);

AND2x2_ASAP7_75t_L g15942 ( 
.A(n_15271),
.B(n_14731),
.Y(n_15942)
);

INVx1_ASAP7_75t_L g15943 ( 
.A(n_15303),
.Y(n_15943)
);

INVx2_ASAP7_75t_L g15944 ( 
.A(n_15365),
.Y(n_15944)
);

AND2x2_ASAP7_75t_L g15945 ( 
.A(n_15473),
.B(n_14735),
.Y(n_15945)
);

NOR2x1_ASAP7_75t_L g15946 ( 
.A(n_15234),
.B(n_14833),
.Y(n_15946)
);

NAND2xp5_ASAP7_75t_L g15947 ( 
.A(n_15729),
.B(n_15000),
.Y(n_15947)
);

INVx1_ASAP7_75t_L g15948 ( 
.A(n_15312),
.Y(n_15948)
);

OR2x2_ASAP7_75t_L g15949 ( 
.A(n_15652),
.B(n_14844),
.Y(n_15949)
);

NAND2xp5_ASAP7_75t_L g15950 ( 
.A(n_15729),
.B(n_15007),
.Y(n_15950)
);

AND2x4_ASAP7_75t_L g15951 ( 
.A(n_15430),
.B(n_14740),
.Y(n_15951)
);

NOR3xp33_ASAP7_75t_L g15952 ( 
.A(n_15526),
.B(n_15101),
.C(n_15100),
.Y(n_15952)
);

A2O1A1Ixp33_ASAP7_75t_SL g15953 ( 
.A1(n_15153),
.A2(n_15254),
.B(n_15248),
.C(n_15243),
.Y(n_15953)
);

AND2x4_ASAP7_75t_L g15954 ( 
.A(n_15436),
.B(n_14747),
.Y(n_15954)
);

INVx1_ASAP7_75t_L g15955 ( 
.A(n_15426),
.Y(n_15955)
);

INVx1_ASAP7_75t_L g15956 ( 
.A(n_15448),
.Y(n_15956)
);

INVx2_ASAP7_75t_L g15957 ( 
.A(n_15365),
.Y(n_15957)
);

NAND2xp5_ASAP7_75t_L g15958 ( 
.A(n_15742),
.B(n_15019),
.Y(n_15958)
);

AND2x2_ASAP7_75t_L g15959 ( 
.A(n_15474),
.B(n_15457),
.Y(n_15959)
);

INVx1_ASAP7_75t_SL g15960 ( 
.A(n_15240),
.Y(n_15960)
);

INVx1_ASAP7_75t_L g15961 ( 
.A(n_15158),
.Y(n_15961)
);

OR2x2_ASAP7_75t_L g15962 ( 
.A(n_15400),
.B(n_14850),
.Y(n_15962)
);

AND2x4_ASAP7_75t_L g15963 ( 
.A(n_15465),
.B(n_14752),
.Y(n_15963)
);

AND2x2_ASAP7_75t_L g15964 ( 
.A(n_15206),
.B(n_14753),
.Y(n_15964)
);

AND2x2_ASAP7_75t_L g15965 ( 
.A(n_15387),
.B(n_14755),
.Y(n_15965)
);

INVx1_ASAP7_75t_L g15966 ( 
.A(n_15185),
.Y(n_15966)
);

NAND3xp33_ASAP7_75t_L g15967 ( 
.A(n_15260),
.B(n_14912),
.C(n_14663),
.Y(n_15967)
);

NAND2xp5_ASAP7_75t_L g15968 ( 
.A(n_15742),
.B(n_15022),
.Y(n_15968)
);

NAND3xp33_ASAP7_75t_L g15969 ( 
.A(n_15234),
.B(n_14823),
.C(n_14623),
.Y(n_15969)
);

INVx1_ASAP7_75t_L g15970 ( 
.A(n_15195),
.Y(n_15970)
);

AND2x2_ASAP7_75t_L g15971 ( 
.A(n_15156),
.B(n_14756),
.Y(n_15971)
);

OR2x2_ASAP7_75t_L g15972 ( 
.A(n_15783),
.B(n_14863),
.Y(n_15972)
);

INVx1_ASAP7_75t_L g15973 ( 
.A(n_15227),
.Y(n_15973)
);

AND2x2_ASAP7_75t_L g15974 ( 
.A(n_15190),
.B(n_14758),
.Y(n_15974)
);

INVx1_ASAP7_75t_L g15975 ( 
.A(n_15508),
.Y(n_15975)
);

INVx2_ASAP7_75t_L g15976 ( 
.A(n_15242),
.Y(n_15976)
);

AND2x2_ASAP7_75t_L g15977 ( 
.A(n_15398),
.B(n_14865),
.Y(n_15977)
);

AND2x2_ASAP7_75t_L g15978 ( 
.A(n_15656),
.B(n_14891),
.Y(n_15978)
);

AND2x2_ASAP7_75t_L g15979 ( 
.A(n_15656),
.B(n_14892),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15518),
.Y(n_15980)
);

INVx2_ASAP7_75t_L g15981 ( 
.A(n_15242),
.Y(n_15981)
);

AND2x2_ASAP7_75t_L g15982 ( 
.A(n_15380),
.B(n_15443),
.Y(n_15982)
);

HB1xp67_ASAP7_75t_L g15983 ( 
.A(n_15192),
.Y(n_15983)
);

HB1xp67_ASAP7_75t_L g15984 ( 
.A(n_15192),
.Y(n_15984)
);

AND2x2_ASAP7_75t_L g15985 ( 
.A(n_15443),
.B(n_14893),
.Y(n_15985)
);

NAND2xp5_ASAP7_75t_L g15986 ( 
.A(n_15783),
.B(n_14902),
.Y(n_15986)
);

INVx1_ASAP7_75t_L g15987 ( 
.A(n_15786),
.Y(n_15987)
);

HB1xp67_ASAP7_75t_L g15988 ( 
.A(n_15482),
.Y(n_15988)
);

NAND2xp5_ASAP7_75t_L g15989 ( 
.A(n_15786),
.B(n_14908),
.Y(n_15989)
);

HB1xp67_ASAP7_75t_L g15990 ( 
.A(n_15331),
.Y(n_15990)
);

AND2x2_ASAP7_75t_L g15991 ( 
.A(n_15282),
.B(n_14919),
.Y(n_15991)
);

INVx1_ASAP7_75t_L g15992 ( 
.A(n_15358),
.Y(n_15992)
);

INVx2_ASAP7_75t_L g15993 ( 
.A(n_15189),
.Y(n_15993)
);

INVx1_ASAP7_75t_L g15994 ( 
.A(n_15226),
.Y(n_15994)
);

AND2x4_ASAP7_75t_SL g15995 ( 
.A(n_15432),
.B(n_14921),
.Y(n_15995)
);

NAND2xp5_ASAP7_75t_L g15996 ( 
.A(n_15295),
.B(n_14925),
.Y(n_15996)
);

INVx2_ASAP7_75t_L g15997 ( 
.A(n_15257),
.Y(n_15997)
);

AND2x2_ASAP7_75t_L g15998 ( 
.A(n_15225),
.B(n_14926),
.Y(n_15998)
);

OR2x2_ASAP7_75t_L g15999 ( 
.A(n_15285),
.B(n_14471),
.Y(n_15999)
);

AND2x4_ASAP7_75t_L g16000 ( 
.A(n_15470),
.B(n_14935),
.Y(n_16000)
);

INVx1_ASAP7_75t_L g16001 ( 
.A(n_15377),
.Y(n_16001)
);

NAND2x1p5_ASAP7_75t_L g16002 ( 
.A(n_15191),
.B(n_15106),
.Y(n_16002)
);

AND2x2_ASAP7_75t_L g16003 ( 
.A(n_15324),
.B(n_14936),
.Y(n_16003)
);

INVx1_ASAP7_75t_L g16004 ( 
.A(n_15799),
.Y(n_16004)
);

AND2x2_ASAP7_75t_L g16005 ( 
.A(n_15490),
.B(n_14939),
.Y(n_16005)
);

NAND4xp25_ASAP7_75t_L g16006 ( 
.A(n_15188),
.B(n_14644),
.C(n_14640),
.D(n_14832),
.Y(n_16006)
);

AND2x2_ASAP7_75t_L g16007 ( 
.A(n_15450),
.B(n_14947),
.Y(n_16007)
);

AND2x2_ASAP7_75t_L g16008 ( 
.A(n_15223),
.B(n_14951),
.Y(n_16008)
);

AND2x2_ASAP7_75t_L g16009 ( 
.A(n_15562),
.B(n_14922),
.Y(n_16009)
);

INVx1_ASAP7_75t_L g16010 ( 
.A(n_15799),
.Y(n_16010)
);

INVx2_ASAP7_75t_L g16011 ( 
.A(n_15280),
.Y(n_16011)
);

NAND2xp67_ASAP7_75t_L g16012 ( 
.A(n_15151),
.B(n_14945),
.Y(n_16012)
);

NAND2xp5_ASAP7_75t_SL g16013 ( 
.A(n_15453),
.B(n_14724),
.Y(n_16013)
);

AND2x2_ASAP7_75t_L g16014 ( 
.A(n_15255),
.B(n_15026),
.Y(n_16014)
);

INVx2_ASAP7_75t_L g16015 ( 
.A(n_15698),
.Y(n_16015)
);

AND2x2_ASAP7_75t_L g16016 ( 
.A(n_15273),
.B(n_15108),
.Y(n_16016)
);

NAND2xp5_ASAP7_75t_L g16017 ( 
.A(n_15840),
.B(n_15128),
.Y(n_16017)
);

INVx2_ASAP7_75t_L g16018 ( 
.A(n_15662),
.Y(n_16018)
);

INVx1_ASAP7_75t_L g16019 ( 
.A(n_15499),
.Y(n_16019)
);

OR2x2_ASAP7_75t_L g16020 ( 
.A(n_15164),
.B(n_15066),
.Y(n_16020)
);

INVx2_ASAP7_75t_L g16021 ( 
.A(n_15662),
.Y(n_16021)
);

AND2x2_ASAP7_75t_L g16022 ( 
.A(n_15371),
.B(n_15205),
.Y(n_16022)
);

INVx1_ASAP7_75t_L g16023 ( 
.A(n_15686),
.Y(n_16023)
);

INVx1_ASAP7_75t_L g16024 ( 
.A(n_15165),
.Y(n_16024)
);

INVx1_ASAP7_75t_L g16025 ( 
.A(n_15407),
.Y(n_16025)
);

INVx1_ASAP7_75t_L g16026 ( 
.A(n_15299),
.Y(n_16026)
);

INVx1_ASAP7_75t_L g16027 ( 
.A(n_15340),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15166),
.Y(n_16028)
);

INVx1_ASAP7_75t_L g16029 ( 
.A(n_15179),
.Y(n_16029)
);

AND2x2_ASAP7_75t_L g16030 ( 
.A(n_15317),
.B(n_15110),
.Y(n_16030)
);

INVx1_ASAP7_75t_L g16031 ( 
.A(n_15717),
.Y(n_16031)
);

NAND2xp5_ASAP7_75t_L g16032 ( 
.A(n_15507),
.B(n_15136),
.Y(n_16032)
);

NAND2xp5_ASAP7_75t_L g16033 ( 
.A(n_15507),
.B(n_14950),
.Y(n_16033)
);

NAND2xp5_ASAP7_75t_L g16034 ( 
.A(n_15483),
.B(n_15115),
.Y(n_16034)
);

INVx2_ASAP7_75t_L g16035 ( 
.A(n_15627),
.Y(n_16035)
);

INVx1_ASAP7_75t_SL g16036 ( 
.A(n_15140),
.Y(n_16036)
);

OR2x2_ASAP7_75t_L g16037 ( 
.A(n_15452),
.B(n_14695),
.Y(n_16037)
);

INVx1_ASAP7_75t_SL g16038 ( 
.A(n_15638),
.Y(n_16038)
);

AOI21xp33_ASAP7_75t_SL g16039 ( 
.A1(n_15261),
.A2(n_15327),
.B(n_15458),
.Y(n_16039)
);

INVx2_ASAP7_75t_L g16040 ( 
.A(n_15627),
.Y(n_16040)
);

NAND2xp5_ASAP7_75t_L g16041 ( 
.A(n_15801),
.B(n_15121),
.Y(n_16041)
);

INVx2_ASAP7_75t_L g16042 ( 
.A(n_15425),
.Y(n_16042)
);

INVx2_ASAP7_75t_L g16043 ( 
.A(n_15494),
.Y(n_16043)
);

INVx1_ASAP7_75t_L g16044 ( 
.A(n_15542),
.Y(n_16044)
);

NAND2xp5_ASAP7_75t_L g16045 ( 
.A(n_15711),
.B(n_14501),
.Y(n_16045)
);

INVx1_ASAP7_75t_L g16046 ( 
.A(n_15648),
.Y(n_16046)
);

NAND2xp5_ASAP7_75t_L g16047 ( 
.A(n_15778),
.B(n_14968),
.Y(n_16047)
);

INVx1_ASAP7_75t_L g16048 ( 
.A(n_15610),
.Y(n_16048)
);

NAND2xp5_ASAP7_75t_L g16049 ( 
.A(n_15748),
.B(n_14825),
.Y(n_16049)
);

NOR2xp33_ASAP7_75t_L g16050 ( 
.A(n_15147),
.B(n_14745),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15239),
.B(n_15010),
.Y(n_16051)
);

INVx2_ASAP7_75t_L g16052 ( 
.A(n_15510),
.Y(n_16052)
);

INVx1_ASAP7_75t_L g16053 ( 
.A(n_15176),
.Y(n_16053)
);

NAND2xp33_ASAP7_75t_R g16054 ( 
.A(n_15526),
.B(n_15046),
.Y(n_16054)
);

OR2x2_ASAP7_75t_L g16055 ( 
.A(n_15492),
.B(n_15073),
.Y(n_16055)
);

AND2x2_ASAP7_75t_L g16056 ( 
.A(n_15523),
.B(n_14553),
.Y(n_16056)
);

BUFx2_ASAP7_75t_L g16057 ( 
.A(n_15245),
.Y(n_16057)
);

INVx1_ASAP7_75t_L g16058 ( 
.A(n_15181),
.Y(n_16058)
);

AND2x2_ASAP7_75t_L g16059 ( 
.A(n_15579),
.B(n_14560),
.Y(n_16059)
);

AND2x2_ASAP7_75t_L g16060 ( 
.A(n_15589),
.B(n_14566),
.Y(n_16060)
);

NOR2xp33_ASAP7_75t_L g16061 ( 
.A(n_15336),
.B(n_14984),
.Y(n_16061)
);

NAND2xp5_ASAP7_75t_L g16062 ( 
.A(n_15350),
.B(n_15475),
.Y(n_16062)
);

NAND2xp5_ASAP7_75t_L g16063 ( 
.A(n_15454),
.B(n_15030),
.Y(n_16063)
);

OR2x2_ASAP7_75t_L g16064 ( 
.A(n_15393),
.B(n_14845),
.Y(n_16064)
);

AND2x2_ASAP7_75t_L g16065 ( 
.A(n_15516),
.B(n_14568),
.Y(n_16065)
);

AND2x2_ASAP7_75t_L g16066 ( 
.A(n_15263),
.B(n_14582),
.Y(n_16066)
);

INVx2_ASAP7_75t_L g16067 ( 
.A(n_15524),
.Y(n_16067)
);

INVx2_ASAP7_75t_L g16068 ( 
.A(n_15484),
.Y(n_16068)
);

OR2x2_ASAP7_75t_L g16069 ( 
.A(n_15233),
.B(n_15289),
.Y(n_16069)
);

NAND2xp5_ASAP7_75t_L g16070 ( 
.A(n_15455),
.B(n_14612),
.Y(n_16070)
);

AND2x2_ASAP7_75t_L g16071 ( 
.A(n_15623),
.B(n_14617),
.Y(n_16071)
);

INVx1_ASAP7_75t_L g16072 ( 
.A(n_15187),
.Y(n_16072)
);

INVx1_ASAP7_75t_L g16073 ( 
.A(n_15196),
.Y(n_16073)
);

AND2x2_ASAP7_75t_L g16074 ( 
.A(n_15640),
.B(n_11903),
.Y(n_16074)
);

OR2x2_ASAP7_75t_L g16075 ( 
.A(n_15152),
.B(n_14515),
.Y(n_16075)
);

INVx1_ASAP7_75t_L g16076 ( 
.A(n_15207),
.Y(n_16076)
);

INVx1_ASAP7_75t_L g16077 ( 
.A(n_15209),
.Y(n_16077)
);

OAI21xp33_ASAP7_75t_L g16078 ( 
.A1(n_15362),
.A2(n_14343),
.B(n_14783),
.Y(n_16078)
);

OR2x2_ASAP7_75t_L g16079 ( 
.A(n_15235),
.B(n_11910),
.Y(n_16079)
);

INVx1_ASAP7_75t_L g16080 ( 
.A(n_15423),
.Y(n_16080)
);

AND2x6_ASAP7_75t_SL g16081 ( 
.A(n_15339),
.B(n_9434),
.Y(n_16081)
);

AND2x2_ASAP7_75t_L g16082 ( 
.A(n_15485),
.B(n_11912),
.Y(n_16082)
);

INVx1_ASAP7_75t_L g16083 ( 
.A(n_15724),
.Y(n_16083)
);

AND2x2_ASAP7_75t_L g16084 ( 
.A(n_15215),
.B(n_11915),
.Y(n_16084)
);

AND2x4_ASAP7_75t_L g16085 ( 
.A(n_15160),
.B(n_9165),
.Y(n_16085)
);

INVx2_ASAP7_75t_L g16086 ( 
.A(n_15666),
.Y(n_16086)
);

INVx1_ASAP7_75t_L g16087 ( 
.A(n_15630),
.Y(n_16087)
);

AND2x2_ASAP7_75t_L g16088 ( 
.A(n_15238),
.B(n_11918),
.Y(n_16088)
);

INVx1_ASAP7_75t_L g16089 ( 
.A(n_15642),
.Y(n_16089)
);

AND2x2_ASAP7_75t_L g16090 ( 
.A(n_15359),
.B(n_11919),
.Y(n_16090)
);

NAND2xp5_ASAP7_75t_L g16091 ( 
.A(n_15464),
.B(n_14963),
.Y(n_16091)
);

AND2x2_ASAP7_75t_L g16092 ( 
.A(n_15363),
.B(n_11923),
.Y(n_16092)
);

NOR3xp33_ASAP7_75t_SL g16093 ( 
.A(n_15721),
.B(n_14906),
.C(n_9470),
.Y(n_16093)
);

AOI22xp5_ASAP7_75t_L g16094 ( 
.A1(n_15609),
.A2(n_14948),
.B1(n_15044),
.B2(n_10759),
.Y(n_16094)
);

OR2x2_ASAP7_75t_L g16095 ( 
.A(n_15404),
.B(n_11928),
.Y(n_16095)
);

INVx1_ASAP7_75t_L g16096 ( 
.A(n_15655),
.Y(n_16096)
);

AND2x2_ASAP7_75t_L g16097 ( 
.A(n_15351),
.B(n_11930),
.Y(n_16097)
);

INVx1_ASAP7_75t_SL g16098 ( 
.A(n_15659),
.Y(n_16098)
);

AND2x4_ASAP7_75t_L g16099 ( 
.A(n_15527),
.B(n_9165),
.Y(n_16099)
);

INVx1_ASAP7_75t_L g16100 ( 
.A(n_15764),
.Y(n_16100)
);

AND2x2_ASAP7_75t_L g16101 ( 
.A(n_15571),
.B(n_15544),
.Y(n_16101)
);

INVx3_ASAP7_75t_L g16102 ( 
.A(n_15364),
.Y(n_16102)
);

NAND2xp5_ASAP7_75t_L g16103 ( 
.A(n_15593),
.B(n_8520),
.Y(n_16103)
);

NAND2xp5_ASAP7_75t_L g16104 ( 
.A(n_15641),
.B(n_8532),
.Y(n_16104)
);

HB1xp67_ASAP7_75t_L g16105 ( 
.A(n_15433),
.Y(n_16105)
);

NAND2xp5_ASAP7_75t_SL g16106 ( 
.A(n_15150),
.B(n_10538),
.Y(n_16106)
);

AND2x2_ASAP7_75t_L g16107 ( 
.A(n_15476),
.B(n_15540),
.Y(n_16107)
);

INVx2_ASAP7_75t_L g16108 ( 
.A(n_15671),
.Y(n_16108)
);

INVx2_ASAP7_75t_L g16109 ( 
.A(n_15683),
.Y(n_16109)
);

NAND2xp5_ASAP7_75t_L g16110 ( 
.A(n_15374),
.B(n_8532),
.Y(n_16110)
);

AND2x4_ASAP7_75t_L g16111 ( 
.A(n_15300),
.B(n_9165),
.Y(n_16111)
);

NAND3xp33_ASAP7_75t_L g16112 ( 
.A(n_15461),
.B(n_11263),
.C(n_11252),
.Y(n_16112)
);

INVx2_ASAP7_75t_L g16113 ( 
.A(n_15694),
.Y(n_16113)
);

INVx1_ASAP7_75t_L g16114 ( 
.A(n_15789),
.Y(n_16114)
);

AND2x2_ASAP7_75t_L g16115 ( 
.A(n_15548),
.B(n_11932),
.Y(n_16115)
);

AND2x2_ASAP7_75t_L g16116 ( 
.A(n_15560),
.B(n_11935),
.Y(n_16116)
);

AND2x2_ASAP7_75t_L g16117 ( 
.A(n_15595),
.B(n_11938),
.Y(n_16117)
);

INVx2_ASAP7_75t_L g16118 ( 
.A(n_15689),
.Y(n_16118)
);

OR2x2_ASAP7_75t_L g16119 ( 
.A(n_15493),
.B(n_11941),
.Y(n_16119)
);

AND2x2_ASAP7_75t_L g16120 ( 
.A(n_15599),
.B(n_11944),
.Y(n_16120)
);

INVx2_ASAP7_75t_L g16121 ( 
.A(n_15682),
.Y(n_16121)
);

INVxp33_ASAP7_75t_L g16122 ( 
.A(n_15292),
.Y(n_16122)
);

NAND2xp33_ASAP7_75t_SL g16123 ( 
.A(n_15434),
.B(n_10759),
.Y(n_16123)
);

NAND2xp5_ASAP7_75t_L g16124 ( 
.A(n_15429),
.B(n_8966),
.Y(n_16124)
);

INVx1_ASAP7_75t_L g16125 ( 
.A(n_15810),
.Y(n_16125)
);

NOR2xp33_ASAP7_75t_L g16126 ( 
.A(n_15591),
.B(n_10759),
.Y(n_16126)
);

AND2x2_ASAP7_75t_L g16127 ( 
.A(n_15601),
.B(n_11947),
.Y(n_16127)
);

NAND2x1_ASAP7_75t_L g16128 ( 
.A(n_15594),
.B(n_11495),
.Y(n_16128)
);

INVx2_ASAP7_75t_L g16129 ( 
.A(n_15605),
.Y(n_16129)
);

INVx1_ASAP7_75t_SL g16130 ( 
.A(n_15590),
.Y(n_16130)
);

AND2x2_ASAP7_75t_L g16131 ( 
.A(n_15395),
.B(n_11951),
.Y(n_16131)
);

INVx2_ASAP7_75t_L g16132 ( 
.A(n_15649),
.Y(n_16132)
);

AND2x2_ASAP7_75t_L g16133 ( 
.A(n_15503),
.B(n_11954),
.Y(n_16133)
);

NAND2xp5_ASAP7_75t_L g16134 ( 
.A(n_15360),
.B(n_8966),
.Y(n_16134)
);

NAND2xp5_ASAP7_75t_L g16135 ( 
.A(n_15386),
.B(n_11956),
.Y(n_16135)
);

INVx2_ASAP7_75t_L g16136 ( 
.A(n_15306),
.Y(n_16136)
);

OR2x2_ASAP7_75t_L g16137 ( 
.A(n_15337),
.B(n_11957),
.Y(n_16137)
);

OAI21xp5_ASAP7_75t_L g16138 ( 
.A1(n_15478),
.A2(n_12062),
.B(n_11447),
.Y(n_16138)
);

INVx1_ASAP7_75t_L g16139 ( 
.A(n_15856),
.Y(n_16139)
);

AND2x2_ASAP7_75t_L g16140 ( 
.A(n_15329),
.B(n_15333),
.Y(n_16140)
);

INVx2_ASAP7_75t_L g16141 ( 
.A(n_15354),
.Y(n_16141)
);

AND2x2_ASAP7_75t_L g16142 ( 
.A(n_15334),
.B(n_11958),
.Y(n_16142)
);

AND2x2_ASAP7_75t_L g16143 ( 
.A(n_15372),
.B(n_11963),
.Y(n_16143)
);

OR2x2_ASAP7_75t_L g16144 ( 
.A(n_15442),
.B(n_15469),
.Y(n_16144)
);

OR2x2_ASAP7_75t_L g16145 ( 
.A(n_15435),
.B(n_11968),
.Y(n_16145)
);

AND2x4_ASAP7_75t_L g16146 ( 
.A(n_15463),
.B(n_8469),
.Y(n_16146)
);

AND2x4_ASAP7_75t_L g16147 ( 
.A(n_15335),
.B(n_8469),
.Y(n_16147)
);

NOR2xp67_ASAP7_75t_L g16148 ( 
.A(n_15178),
.B(n_10613),
.Y(n_16148)
);

INVx2_ASAP7_75t_L g16149 ( 
.A(n_15388),
.Y(n_16149)
);

HB1xp67_ASAP7_75t_L g16150 ( 
.A(n_15563),
.Y(n_16150)
);

INVxp67_ASAP7_75t_SL g16151 ( 
.A(n_15797),
.Y(n_16151)
);

INVx1_ASAP7_75t_L g16152 ( 
.A(n_15673),
.Y(n_16152)
);

INVx1_ASAP7_75t_L g16153 ( 
.A(n_15690),
.Y(n_16153)
);

AND2x2_ASAP7_75t_L g16154 ( 
.A(n_15384),
.B(n_11971),
.Y(n_16154)
);

INVx1_ASAP7_75t_L g16155 ( 
.A(n_15550),
.Y(n_16155)
);

AND2x2_ASAP7_75t_L g16156 ( 
.A(n_15291),
.B(n_11973),
.Y(n_16156)
);

NAND2xp5_ASAP7_75t_L g16157 ( 
.A(n_15832),
.B(n_15860),
.Y(n_16157)
);

AND2x2_ASAP7_75t_L g16158 ( 
.A(n_15291),
.B(n_11975),
.Y(n_16158)
);

AND2x2_ASAP7_75t_L g16159 ( 
.A(n_15530),
.B(n_11976),
.Y(n_16159)
);

INVx2_ASAP7_75t_L g16160 ( 
.A(n_15412),
.Y(n_16160)
);

HB1xp67_ASAP7_75t_L g16161 ( 
.A(n_15637),
.Y(n_16161)
);

AOI211xp5_ASAP7_75t_L g16162 ( 
.A1(n_15489),
.A2(n_11266),
.B(n_11535),
.C(n_12062),
.Y(n_16162)
);

INVx1_ASAP7_75t_L g16163 ( 
.A(n_15553),
.Y(n_16163)
);

INVx2_ASAP7_75t_L g16164 ( 
.A(n_15713),
.Y(n_16164)
);

INVx2_ASAP7_75t_L g16165 ( 
.A(n_15456),
.Y(n_16165)
);

INVx1_ASAP7_75t_L g16166 ( 
.A(n_15558),
.Y(n_16166)
);

HB1xp67_ASAP7_75t_L g16167 ( 
.A(n_15258),
.Y(n_16167)
);

NAND2xp5_ASAP7_75t_L g16168 ( 
.A(n_15860),
.B(n_11978),
.Y(n_16168)
);

NAND2xp5_ASAP7_75t_L g16169 ( 
.A(n_15582),
.B(n_11984),
.Y(n_16169)
);

INVx1_ASAP7_75t_L g16170 ( 
.A(n_15570),
.Y(n_16170)
);

AND2x4_ASAP7_75t_L g16171 ( 
.A(n_15213),
.B(n_8469),
.Y(n_16171)
);

BUFx2_ASAP7_75t_SL g16172 ( 
.A(n_15356),
.Y(n_16172)
);

INVx1_ASAP7_75t_L g16173 ( 
.A(n_15602),
.Y(n_16173)
);

HB1xp67_ASAP7_75t_L g16174 ( 
.A(n_15267),
.Y(n_16174)
);

INVx1_ASAP7_75t_L g16175 ( 
.A(n_15172),
.Y(n_16175)
);

INVx4_ASAP7_75t_L g16176 ( 
.A(n_15456),
.Y(n_16176)
);

INVx1_ASAP7_75t_L g16177 ( 
.A(n_15174),
.Y(n_16177)
);

INVx2_ASAP7_75t_L g16178 ( 
.A(n_15613),
.Y(n_16178)
);

AND2x2_ASAP7_75t_L g16179 ( 
.A(n_15531),
.B(n_11989),
.Y(n_16179)
);

NAND2x1p5_ASAP7_75t_L g16180 ( 
.A(n_15419),
.B(n_9329),
.Y(n_16180)
);

INVx1_ASAP7_75t_L g16181 ( 
.A(n_15214),
.Y(n_16181)
);

OR2x2_ASAP7_75t_L g16182 ( 
.A(n_15269),
.B(n_11994),
.Y(n_16182)
);

INVx2_ASAP7_75t_SL g16183 ( 
.A(n_15178),
.Y(n_16183)
);

AND2x2_ASAP7_75t_L g16184 ( 
.A(n_15315),
.B(n_12000),
.Y(n_16184)
);

BUFx2_ASAP7_75t_SL g16185 ( 
.A(n_15178),
.Y(n_16185)
);

NAND2x1p5_ASAP7_75t_L g16186 ( 
.A(n_15419),
.B(n_9329),
.Y(n_16186)
);

BUFx2_ASAP7_75t_L g16187 ( 
.A(n_15264),
.Y(n_16187)
);

HB1xp67_ASAP7_75t_L g16188 ( 
.A(n_15661),
.Y(n_16188)
);

INVx2_ASAP7_75t_L g16189 ( 
.A(n_15330),
.Y(n_16189)
);

AND2x2_ASAP7_75t_L g16190 ( 
.A(n_15481),
.B(n_12006),
.Y(n_16190)
);

NAND2xp5_ASAP7_75t_L g16191 ( 
.A(n_15626),
.B(n_15290),
.Y(n_16191)
);

AND2x2_ASAP7_75t_L g16192 ( 
.A(n_15647),
.B(n_12008),
.Y(n_16192)
);

NAND3xp33_ASAP7_75t_L g16193 ( 
.A(n_15466),
.B(n_11263),
.C(n_11252),
.Y(n_16193)
);

INVx1_ASAP7_75t_L g16194 ( 
.A(n_15155),
.Y(n_16194)
);

AND2x2_ASAP7_75t_L g16195 ( 
.A(n_15564),
.B(n_12009),
.Y(n_16195)
);

INVx2_ASAP7_75t_L g16196 ( 
.A(n_15330),
.Y(n_16196)
);

AND2x2_ASAP7_75t_L g16197 ( 
.A(n_15403),
.B(n_12010),
.Y(n_16197)
);

OR2x2_ASAP7_75t_L g16198 ( 
.A(n_15479),
.B(n_12013),
.Y(n_16198)
);

HB1xp67_ASAP7_75t_L g16199 ( 
.A(n_15338),
.Y(n_16199)
);

NAND3xp33_ASAP7_75t_L g16200 ( 
.A(n_15496),
.B(n_11268),
.C(n_11265),
.Y(n_16200)
);

INVx1_ASAP7_75t_L g16201 ( 
.A(n_15162),
.Y(n_16201)
);

INVx2_ASAP7_75t_L g16202 ( 
.A(n_15330),
.Y(n_16202)
);

NAND2xp5_ASAP7_75t_L g16203 ( 
.A(n_15863),
.B(n_12014),
.Y(n_16203)
);

AND2x2_ASAP7_75t_L g16204 ( 
.A(n_15410),
.B(n_12015),
.Y(n_16204)
);

NOR2xp33_ASAP7_75t_L g16205 ( 
.A(n_15279),
.B(n_10759),
.Y(n_16205)
);

OR2x2_ASAP7_75t_L g16206 ( 
.A(n_15224),
.B(n_12018),
.Y(n_16206)
);

INVx1_ASAP7_75t_L g16207 ( 
.A(n_15163),
.Y(n_16207)
);

INVx3_ASAP7_75t_L g16208 ( 
.A(n_15596),
.Y(n_16208)
);

AND2x2_ASAP7_75t_L g16209 ( 
.A(n_15413),
.B(n_12019),
.Y(n_16209)
);

AND2x2_ASAP7_75t_L g16210 ( 
.A(n_15305),
.B(n_12020),
.Y(n_16210)
);

NAND2xp5_ASAP7_75t_L g16211 ( 
.A(n_15608),
.B(n_12024),
.Y(n_16211)
);

BUFx2_ASAP7_75t_SL g16212 ( 
.A(n_15182),
.Y(n_16212)
);

BUFx2_ASAP7_75t_L g16213 ( 
.A(n_15830),
.Y(n_16213)
);

AND2x2_ASAP7_75t_L g16214 ( 
.A(n_15552),
.B(n_12026),
.Y(n_16214)
);

AND2x4_ASAP7_75t_L g16215 ( 
.A(n_15424),
.B(n_8469),
.Y(n_16215)
);

INVx1_ASAP7_75t_L g16216 ( 
.A(n_15169),
.Y(n_16216)
);

AND2x4_ASAP7_75t_L g16217 ( 
.A(n_15428),
.B(n_8469),
.Y(n_16217)
);

AND2x2_ASAP7_75t_L g16218 ( 
.A(n_15349),
.B(n_12029),
.Y(n_16218)
);

INVx1_ASAP7_75t_L g16219 ( 
.A(n_15170),
.Y(n_16219)
);

INVx1_ASAP7_75t_L g16220 ( 
.A(n_15399),
.Y(n_16220)
);

INVx2_ASAP7_75t_L g16221 ( 
.A(n_15712),
.Y(n_16221)
);

INVx1_ASAP7_75t_L g16222 ( 
.A(n_15533),
.Y(n_16222)
);

NAND2xp5_ASAP7_75t_L g16223 ( 
.A(n_15763),
.B(n_15460),
.Y(n_16223)
);

OR2x2_ASAP7_75t_L g16224 ( 
.A(n_15585),
.B(n_12034),
.Y(n_16224)
);

AND2x2_ASAP7_75t_L g16225 ( 
.A(n_15422),
.B(n_12035),
.Y(n_16225)
);

AND2x4_ASAP7_75t_SL g16226 ( 
.A(n_15557),
.B(n_8072),
.Y(n_16226)
);

AND2x4_ASAP7_75t_L g16227 ( 
.A(n_15246),
.B(n_15222),
.Y(n_16227)
);

AND2x2_ASAP7_75t_L g16228 ( 
.A(n_15427),
.B(n_12036),
.Y(n_16228)
);

HB1xp67_ASAP7_75t_L g16229 ( 
.A(n_15353),
.Y(n_16229)
);

INVx1_ASAP7_75t_L g16230 ( 
.A(n_15211),
.Y(n_16230)
);

NAND2xp5_ASAP7_75t_SL g16231 ( 
.A(n_15512),
.B(n_10538),
.Y(n_16231)
);

NAND2xp5_ASAP7_75t_L g16232 ( 
.A(n_15674),
.B(n_12038),
.Y(n_16232)
);

INVx2_ASAP7_75t_L g16233 ( 
.A(n_15715),
.Y(n_16233)
);

OAI21xp33_ASAP7_75t_L g16234 ( 
.A1(n_15296),
.A2(n_11268),
.B(n_11265),
.Y(n_16234)
);

NAND2xp5_ASAP7_75t_L g16235 ( 
.A(n_15676),
.B(n_12040),
.Y(n_16235)
);

INVx1_ASAP7_75t_SL g16236 ( 
.A(n_15506),
.Y(n_16236)
);

NOR2xp33_ASAP7_75t_L g16237 ( 
.A(n_15408),
.B(n_10568),
.Y(n_16237)
);

NAND2xp5_ASAP7_75t_L g16238 ( 
.A(n_15685),
.B(n_15383),
.Y(n_16238)
);

AND2x2_ASAP7_75t_L g16239 ( 
.A(n_15546),
.B(n_12045),
.Y(n_16239)
);

NAND2xp5_ASAP7_75t_L g16240 ( 
.A(n_15850),
.B(n_12048),
.Y(n_16240)
);

AND2x2_ASAP7_75t_L g16241 ( 
.A(n_15437),
.B(n_12052),
.Y(n_16241)
);

NAND2xp5_ASAP7_75t_L g16242 ( 
.A(n_15616),
.B(n_12057),
.Y(n_16242)
);

INVx2_ASAP7_75t_SL g16243 ( 
.A(n_15182),
.Y(n_16243)
);

AND2x4_ASAP7_75t_L g16244 ( 
.A(n_15611),
.B(n_8469),
.Y(n_16244)
);

NOR2xp33_ASAP7_75t_L g16245 ( 
.A(n_15182),
.B(n_10568),
.Y(n_16245)
);

NAND2xp5_ASAP7_75t_L g16246 ( 
.A(n_15654),
.B(n_12061),
.Y(n_16246)
);

INVx1_ASAP7_75t_L g16247 ( 
.A(n_15216),
.Y(n_16247)
);

INVx1_ASAP7_75t_L g16248 ( 
.A(n_15858),
.Y(n_16248)
);

AND2x2_ASAP7_75t_L g16249 ( 
.A(n_15326),
.B(n_12063),
.Y(n_16249)
);

HB1xp67_ASAP7_75t_SL g16250 ( 
.A(n_15668),
.Y(n_16250)
);

OR2x2_ASAP7_75t_L g16251 ( 
.A(n_15385),
.B(n_12066),
.Y(n_16251)
);

AND2x4_ASAP7_75t_L g16252 ( 
.A(n_15471),
.B(n_8518),
.Y(n_16252)
);

INVx1_ASAP7_75t_L g16253 ( 
.A(n_15665),
.Y(n_16253)
);

AND2x4_ASAP7_75t_SL g16254 ( 
.A(n_15418),
.B(n_8072),
.Y(n_16254)
);

INVx1_ASAP7_75t_L g16255 ( 
.A(n_15745),
.Y(n_16255)
);

BUFx2_ASAP7_75t_L g16256 ( 
.A(n_15788),
.Y(n_16256)
);

NAND2xp5_ASAP7_75t_L g16257 ( 
.A(n_15658),
.B(n_15687),
.Y(n_16257)
);

AND2x2_ASAP7_75t_L g16258 ( 
.A(n_15769),
.B(n_12067),
.Y(n_16258)
);

OR2x2_ASAP7_75t_L g16259 ( 
.A(n_15409),
.B(n_12068),
.Y(n_16259)
);

HB1xp67_ASAP7_75t_L g16260 ( 
.A(n_15653),
.Y(n_16260)
);

INVx2_ASAP7_75t_L g16261 ( 
.A(n_15512),
.Y(n_16261)
);

INVx1_ASAP7_75t_L g16262 ( 
.A(n_15768),
.Y(n_16262)
);

INVx1_ASAP7_75t_L g16263 ( 
.A(n_15622),
.Y(n_16263)
);

AND2x2_ASAP7_75t_L g16264 ( 
.A(n_15749),
.B(n_12070),
.Y(n_16264)
);

AND2x4_ASAP7_75t_L g16265 ( 
.A(n_15379),
.B(n_14082),
.Y(n_16265)
);

NAND2xp5_ASAP7_75t_L g16266 ( 
.A(n_15699),
.B(n_12071),
.Y(n_16266)
);

HB1xp67_ASAP7_75t_L g16267 ( 
.A(n_15446),
.Y(n_16267)
);

NAND2xp5_ASAP7_75t_L g16268 ( 
.A(n_15705),
.B(n_12079),
.Y(n_16268)
);

AND2x4_ASAP7_75t_L g16269 ( 
.A(n_15477),
.B(n_14082),
.Y(n_16269)
);

INVx2_ASAP7_75t_L g16270 ( 
.A(n_15265),
.Y(n_16270)
);

INVx1_ASAP7_75t_L g16271 ( 
.A(n_15744),
.Y(n_16271)
);

INVx1_ASAP7_75t_L g16272 ( 
.A(n_15751),
.Y(n_16272)
);

INVx1_ASAP7_75t_L g16273 ( 
.A(n_15759),
.Y(n_16273)
);

INVx1_ASAP7_75t_L g16274 ( 
.A(n_15760),
.Y(n_16274)
);

OR2x6_ASAP7_75t_L g16275 ( 
.A(n_15417),
.B(n_10568),
.Y(n_16275)
);

AND2x2_ASAP7_75t_L g16276 ( 
.A(n_15761),
.B(n_12080),
.Y(n_16276)
);

NAND2xp5_ASAP7_75t_L g16277 ( 
.A(n_15732),
.B(n_12083),
.Y(n_16277)
);

AND2x2_ASAP7_75t_L g16278 ( 
.A(n_15449),
.B(n_12086),
.Y(n_16278)
);

AND2x4_ASAP7_75t_L g16279 ( 
.A(n_15487),
.B(n_8518),
.Y(n_16279)
);

AND2x2_ASAP7_75t_L g16280 ( 
.A(n_15444),
.B(n_12087),
.Y(n_16280)
);

OAI221xp5_ASAP7_75t_SL g16281 ( 
.A1(n_15835),
.A2(n_11499),
.B1(n_11500),
.B2(n_11498),
.C(n_11497),
.Y(n_16281)
);

AND2x2_ASAP7_75t_L g16282 ( 
.A(n_15445),
.B(n_15325),
.Y(n_16282)
);

AND2x2_ASAP7_75t_L g16283 ( 
.A(n_15725),
.B(n_12091),
.Y(n_16283)
);

AND2x4_ASAP7_75t_L g16284 ( 
.A(n_15488),
.B(n_8518),
.Y(n_16284)
);

AND2x2_ASAP7_75t_L g16285 ( 
.A(n_15684),
.B(n_12092),
.Y(n_16285)
);

NAND2xp5_ASAP7_75t_L g16286 ( 
.A(n_15639),
.B(n_12097),
.Y(n_16286)
);

NAND2xp5_ASAP7_75t_L g16287 ( 
.A(n_15459),
.B(n_12100),
.Y(n_16287)
);

HB1xp67_ASAP7_75t_L g16288 ( 
.A(n_15345),
.Y(n_16288)
);

OR2x2_ASAP7_75t_L g16289 ( 
.A(n_15402),
.B(n_12102),
.Y(n_16289)
);

INVx1_ASAP7_75t_L g16290 ( 
.A(n_15831),
.Y(n_16290)
);

NAND2xp5_ASAP7_75t_L g16291 ( 
.A(n_15462),
.B(n_15468),
.Y(n_16291)
);

INVxp67_ASAP7_75t_L g16292 ( 
.A(n_15390),
.Y(n_16292)
);

AND2x4_ASAP7_75t_L g16293 ( 
.A(n_15232),
.B(n_8518),
.Y(n_16293)
);

NAND2xp5_ASAP7_75t_L g16294 ( 
.A(n_15486),
.B(n_12108),
.Y(n_16294)
);

AND2x2_ASAP7_75t_L g16295 ( 
.A(n_15833),
.B(n_12109),
.Y(n_16295)
);

AND2x2_ASAP7_75t_L g16296 ( 
.A(n_15612),
.B(n_15620),
.Y(n_16296)
);

NAND2xp5_ASAP7_75t_L g16297 ( 
.A(n_15603),
.B(n_12112),
.Y(n_16297)
);

OR2x2_ASAP7_75t_L g16298 ( 
.A(n_15394),
.B(n_12114),
.Y(n_16298)
);

AND2x2_ASAP7_75t_L g16299 ( 
.A(n_15625),
.B(n_12116),
.Y(n_16299)
);

NAND2xp5_ASAP7_75t_L g16300 ( 
.A(n_15667),
.B(n_12117),
.Y(n_16300)
);

AND2x2_ASAP7_75t_L g16301 ( 
.A(n_15547),
.B(n_12118),
.Y(n_16301)
);

OR2x2_ASAP7_75t_L g16302 ( 
.A(n_15401),
.B(n_12130),
.Y(n_16302)
);

INVx2_ASAP7_75t_L g16303 ( 
.A(n_15727),
.Y(n_16303)
);

INVx2_ASAP7_75t_L g16304 ( 
.A(n_15731),
.Y(n_16304)
);

BUFx2_ASAP7_75t_L g16305 ( 
.A(n_15814),
.Y(n_16305)
);

AND2x2_ASAP7_75t_L g16306 ( 
.A(n_15284),
.B(n_12134),
.Y(n_16306)
);

HB1xp67_ASAP7_75t_L g16307 ( 
.A(n_15347),
.Y(n_16307)
);

NAND2xp5_ASAP7_75t_L g16308 ( 
.A(n_15675),
.B(n_12135),
.Y(n_16308)
);

INVx1_ASAP7_75t_L g16309 ( 
.A(n_15853),
.Y(n_16309)
);

OAI21xp5_ASAP7_75t_L g16310 ( 
.A1(n_15663),
.A2(n_11266),
.B(n_11535),
.Y(n_16310)
);

NAND2xp5_ASAP7_75t_L g16311 ( 
.A(n_15504),
.B(n_12138),
.Y(n_16311)
);

AND2x4_ASAP7_75t_L g16312 ( 
.A(n_15352),
.B(n_8518),
.Y(n_16312)
);

OR2x2_ASAP7_75t_L g16313 ( 
.A(n_15405),
.B(n_12142),
.Y(n_16313)
);

INVx1_ASAP7_75t_L g16314 ( 
.A(n_15635),
.Y(n_16314)
);

INVx1_ASAP7_75t_L g16315 ( 
.A(n_15869),
.Y(n_16315)
);

INVx3_ASAP7_75t_L g16316 ( 
.A(n_15775),
.Y(n_16316)
);

AND2x4_ASAP7_75t_L g16317 ( 
.A(n_15183),
.B(n_8518),
.Y(n_16317)
);

OR2x2_ASAP7_75t_L g16318 ( 
.A(n_15411),
.B(n_12148),
.Y(n_16318)
);

INVx1_ASAP7_75t_L g16319 ( 
.A(n_15171),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_15498),
.B(n_12162),
.Y(n_16320)
);

AND2x2_ASAP7_75t_L g16321 ( 
.A(n_15505),
.B(n_12163),
.Y(n_16321)
);

INVx1_ASAP7_75t_L g16322 ( 
.A(n_15572),
.Y(n_16322)
);

NAND2xp5_ASAP7_75t_L g16323 ( 
.A(n_15728),
.B(n_12164),
.Y(n_16323)
);

INVx2_ASAP7_75t_L g16324 ( 
.A(n_15287),
.Y(n_16324)
);

INVx1_ASAP7_75t_L g16325 ( 
.A(n_15573),
.Y(n_16325)
);

BUFx2_ASAP7_75t_L g16326 ( 
.A(n_15420),
.Y(n_16326)
);

AND2x2_ASAP7_75t_L g16327 ( 
.A(n_15316),
.B(n_12165),
.Y(n_16327)
);

INVx1_ASAP7_75t_L g16328 ( 
.A(n_15583),
.Y(n_16328)
);

AND2x2_ASAP7_75t_L g16329 ( 
.A(n_15703),
.B(n_12172),
.Y(n_16329)
);

AND2x2_ASAP7_75t_L g16330 ( 
.A(n_15706),
.B(n_12178),
.Y(n_16330)
);

OR2x2_ASAP7_75t_L g16331 ( 
.A(n_15415),
.B(n_12179),
.Y(n_16331)
);

INVx1_ASAP7_75t_L g16332 ( 
.A(n_15785),
.Y(n_16332)
);

INVxp67_ASAP7_75t_SL g16333 ( 
.A(n_15149),
.Y(n_16333)
);

INVx1_ASAP7_75t_L g16334 ( 
.A(n_15798),
.Y(n_16334)
);

NAND2xp5_ASAP7_75t_L g16335 ( 
.A(n_15816),
.B(n_12183),
.Y(n_16335)
);

BUFx3_ASAP7_75t_L g16336 ( 
.A(n_15420),
.Y(n_16336)
);

INVx1_ASAP7_75t_L g16337 ( 
.A(n_15834),
.Y(n_16337)
);

BUFx2_ASAP7_75t_L g16338 ( 
.A(n_15202),
.Y(n_16338)
);

NAND2xp5_ASAP7_75t_SL g16339 ( 
.A(n_15787),
.B(n_10538),
.Y(n_16339)
);

AND2x2_ASAP7_75t_L g16340 ( 
.A(n_15650),
.B(n_12184),
.Y(n_16340)
);

HB1xp67_ASAP7_75t_L g16341 ( 
.A(n_15629),
.Y(n_16341)
);

NAND2xp5_ASAP7_75t_L g16342 ( 
.A(n_15819),
.B(n_15812),
.Y(n_16342)
);

INVx1_ASAP7_75t_L g16343 ( 
.A(n_15848),
.Y(n_16343)
);

OR2x2_ASAP7_75t_L g16344 ( 
.A(n_15416),
.B(n_12187),
.Y(n_16344)
);

INVx1_ASAP7_75t_L g16345 ( 
.A(n_15861),
.Y(n_16345)
);

INVx1_ASAP7_75t_L g16346 ( 
.A(n_15587),
.Y(n_16346)
);

AND2x2_ASAP7_75t_L g16347 ( 
.A(n_15736),
.B(n_12193),
.Y(n_16347)
);

AND2x2_ASAP7_75t_L g16348 ( 
.A(n_15193),
.B(n_12194),
.Y(n_16348)
);

INVx2_ASAP7_75t_L g16349 ( 
.A(n_15287),
.Y(n_16349)
);

AND2x4_ASAP7_75t_L g16350 ( 
.A(n_15197),
.B(n_8555),
.Y(n_16350)
);

AND2x2_ASAP7_75t_L g16351 ( 
.A(n_15201),
.B(n_12196),
.Y(n_16351)
);

INVx2_ASAP7_75t_L g16352 ( 
.A(n_15739),
.Y(n_16352)
);

AND2x2_ASAP7_75t_L g16353 ( 
.A(n_15497),
.B(n_12203),
.Y(n_16353)
);

NAND2xp5_ASAP7_75t_L g16354 ( 
.A(n_15421),
.B(n_12212),
.Y(n_16354)
);

AND2x4_ASAP7_75t_L g16355 ( 
.A(n_15144),
.B(n_8555),
.Y(n_16355)
);

INVx1_ASAP7_75t_L g16356 ( 
.A(n_15619),
.Y(n_16356)
);

OR2x2_ASAP7_75t_L g16357 ( 
.A(n_15439),
.B(n_12214),
.Y(n_16357)
);

NOR2xp67_ASAP7_75t_L g16358 ( 
.A(n_15278),
.B(n_11497),
.Y(n_16358)
);

AND2x2_ASAP7_75t_L g16359 ( 
.A(n_15146),
.B(n_12216),
.Y(n_16359)
);

INVxp67_ASAP7_75t_L g16360 ( 
.A(n_15691),
.Y(n_16360)
);

AND2x2_ASAP7_75t_L g16361 ( 
.A(n_15302),
.B(n_12217),
.Y(n_16361)
);

INVx1_ASAP7_75t_L g16362 ( 
.A(n_15441),
.Y(n_16362)
);

AND2x4_ASAP7_75t_SL g16363 ( 
.A(n_15566),
.B(n_8116),
.Y(n_16363)
);

NAND2xp5_ASAP7_75t_L g16364 ( 
.A(n_15447),
.B(n_12219),
.Y(n_16364)
);

INVx1_ASAP7_75t_L g16365 ( 
.A(n_15451),
.Y(n_16365)
);

NAND2xp5_ASAP7_75t_L g16366 ( 
.A(n_15679),
.B(n_12220),
.Y(n_16366)
);

INVx3_ASAP7_75t_L g16367 ( 
.A(n_15716),
.Y(n_16367)
);

AND2x4_ASAP7_75t_L g16368 ( 
.A(n_15304),
.B(n_15220),
.Y(n_16368)
);

OR2x2_ASAP7_75t_L g16369 ( 
.A(n_15726),
.B(n_12226),
.Y(n_16369)
);

OAI21xp5_ASAP7_75t_L g16370 ( 
.A1(n_15310),
.A2(n_11262),
.B(n_11258),
.Y(n_16370)
);

AND2x4_ASAP7_75t_SL g16371 ( 
.A(n_15633),
.B(n_8116),
.Y(n_16371)
);

INVx1_ASAP7_75t_L g16372 ( 
.A(n_15774),
.Y(n_16372)
);

INVx2_ASAP7_75t_L g16373 ( 
.A(n_15733),
.Y(n_16373)
);

AND2x4_ASAP7_75t_SL g16374 ( 
.A(n_15321),
.B(n_8116),
.Y(n_16374)
);

INVx1_ASAP7_75t_L g16375 ( 
.A(n_15565),
.Y(n_16375)
);

AND2x2_ASAP7_75t_L g16376 ( 
.A(n_15680),
.B(n_15606),
.Y(n_16376)
);

INVx1_ASAP7_75t_L g16377 ( 
.A(n_15664),
.Y(n_16377)
);

INVx1_ASAP7_75t_L g16378 ( 
.A(n_15517),
.Y(n_16378)
);

INVxp67_ASAP7_75t_L g16379 ( 
.A(n_15253),
.Y(n_16379)
);

NOR2xp33_ASAP7_75t_L g16380 ( 
.A(n_15567),
.B(n_10568),
.Y(n_16380)
);

INVx1_ASAP7_75t_L g16381 ( 
.A(n_15719),
.Y(n_16381)
);

INVx1_ASAP7_75t_L g16382 ( 
.A(n_15722),
.Y(n_16382)
);

NAND2xp5_ASAP7_75t_L g16383 ( 
.A(n_15802),
.B(n_12228),
.Y(n_16383)
);

AND2x2_ASAP7_75t_L g16384 ( 
.A(n_15617),
.B(n_12229),
.Y(n_16384)
);

BUFx3_ASAP7_75t_L g16385 ( 
.A(n_15556),
.Y(n_16385)
);

OR2x2_ASAP7_75t_L g16386 ( 
.A(n_15520),
.B(n_12234),
.Y(n_16386)
);

INVx1_ASAP7_75t_L g16387 ( 
.A(n_15247),
.Y(n_16387)
);

INVx1_ASAP7_75t_L g16388 ( 
.A(n_15249),
.Y(n_16388)
);

NAND2xp5_ASAP7_75t_L g16389 ( 
.A(n_15815),
.B(n_12239),
.Y(n_16389)
);

NAND2x1_ASAP7_75t_SL g16390 ( 
.A(n_15256),
.B(n_11498),
.Y(n_16390)
);

INVx2_ASAP7_75t_L g16391 ( 
.A(n_15756),
.Y(n_16391)
);

INVx2_ASAP7_75t_L g16392 ( 
.A(n_15866),
.Y(n_16392)
);

INVx1_ASAP7_75t_L g16393 ( 
.A(n_15250),
.Y(n_16393)
);

AND2x2_ASAP7_75t_L g16394 ( 
.A(n_15704),
.B(n_12243),
.Y(n_16394)
);

AND2x4_ASAP7_75t_L g16395 ( 
.A(n_15577),
.B(n_8555),
.Y(n_16395)
);

AND2x2_ASAP7_75t_L g16396 ( 
.A(n_15746),
.B(n_15750),
.Y(n_16396)
);

NOR2xp33_ASAP7_75t_L g16397 ( 
.A(n_15368),
.B(n_12244),
.Y(n_16397)
);

INVx1_ASAP7_75t_L g16398 ( 
.A(n_15251),
.Y(n_16398)
);

AND2x4_ASAP7_75t_SL g16399 ( 
.A(n_15414),
.B(n_8116),
.Y(n_16399)
);

OR2x2_ASAP7_75t_L g16400 ( 
.A(n_15551),
.B(n_12257),
.Y(n_16400)
);

INVx3_ASAP7_75t_SL g16401 ( 
.A(n_15202),
.Y(n_16401)
);

BUFx2_ASAP7_75t_L g16402 ( 
.A(n_15307),
.Y(n_16402)
);

INVx1_ASAP7_75t_L g16403 ( 
.A(n_15309),
.Y(n_16403)
);

BUFx2_ASAP7_75t_L g16404 ( 
.A(n_15700),
.Y(n_16404)
);

INVx1_ASAP7_75t_L g16405 ( 
.A(n_15311),
.Y(n_16405)
);

INVxp67_ASAP7_75t_SL g16406 ( 
.A(n_15252),
.Y(n_16406)
);

AND2x2_ASAP7_75t_L g16407 ( 
.A(n_15753),
.B(n_12258),
.Y(n_16407)
);

AND2x4_ASAP7_75t_L g16408 ( 
.A(n_15782),
.B(n_8555),
.Y(n_16408)
);

INVx2_ASAP7_75t_L g16409 ( 
.A(n_15771),
.Y(n_16409)
);

INVx1_ASAP7_75t_L g16410 ( 
.A(n_15313),
.Y(n_16410)
);

NAND2xp5_ASAP7_75t_L g16411 ( 
.A(n_15618),
.B(n_12260),
.Y(n_16411)
);

OR2x2_ASAP7_75t_L g16412 ( 
.A(n_15369),
.B(n_8579),
.Y(n_16412)
);

AND2x2_ASAP7_75t_L g16413 ( 
.A(n_15766),
.B(n_9540),
.Y(n_16413)
);

AND2x2_ASAP7_75t_L g16414 ( 
.A(n_15767),
.B(n_9540),
.Y(n_16414)
);

INVx2_ASAP7_75t_L g16415 ( 
.A(n_15692),
.Y(n_16415)
);

NAND2xp5_ASAP7_75t_SL g16416 ( 
.A(n_15809),
.B(n_10538),
.Y(n_16416)
);

AND2x2_ASAP7_75t_L g16417 ( 
.A(n_15701),
.B(n_9548),
.Y(n_16417)
);

AND2x2_ASAP7_75t_L g16418 ( 
.A(n_15792),
.B(n_9548),
.Y(n_16418)
);

INVx1_ASAP7_75t_L g16419 ( 
.A(n_15314),
.Y(n_16419)
);

INVx1_ASAP7_75t_L g16420 ( 
.A(n_15259),
.Y(n_16420)
);

AND2x2_ASAP7_75t_L g16421 ( 
.A(n_15796),
.B(n_9334),
.Y(n_16421)
);

NAND2xp5_ASAP7_75t_L g16422 ( 
.A(n_15807),
.B(n_15491),
.Y(n_16422)
);

AND2x2_ASAP7_75t_L g16423 ( 
.A(n_15770),
.B(n_9334),
.Y(n_16423)
);

INVx1_ASAP7_75t_L g16424 ( 
.A(n_15738),
.Y(n_16424)
);

HB1xp67_ASAP7_75t_L g16425 ( 
.A(n_15714),
.Y(n_16425)
);

AND2x2_ASAP7_75t_L g16426 ( 
.A(n_15791),
.B(n_9334),
.Y(n_16426)
);

INVx1_ASAP7_75t_L g16427 ( 
.A(n_15293),
.Y(n_16427)
);

NAND2xp5_ASAP7_75t_L g16428 ( 
.A(n_15500),
.B(n_9342),
.Y(n_16428)
);

INVx2_ASAP7_75t_L g16429 ( 
.A(n_15803),
.Y(n_16429)
);

NAND2xp5_ASAP7_75t_L g16430 ( 
.A(n_15501),
.B(n_9342),
.Y(n_16430)
);

INVxp33_ASAP7_75t_L g16431 ( 
.A(n_15688),
.Y(n_16431)
);

NAND2xp5_ASAP7_75t_L g16432 ( 
.A(n_15614),
.B(n_9342),
.Y(n_16432)
);

AND2x2_ASAP7_75t_L g16433 ( 
.A(n_15621),
.B(n_9406),
.Y(n_16433)
);

INVxp67_ASAP7_75t_SL g16434 ( 
.A(n_15513),
.Y(n_16434)
);

INVx3_ASAP7_75t_L g16435 ( 
.A(n_15762),
.Y(n_16435)
);

AND2x2_ASAP7_75t_L g16436 ( 
.A(n_15631),
.B(n_9406),
.Y(n_16436)
);

OAI221xp5_ASAP7_75t_SL g16437 ( 
.A1(n_15270),
.A2(n_11503),
.B1(n_11510),
.B2(n_11500),
.C(n_11499),
.Y(n_16437)
);

OR2x2_ASAP7_75t_L g16438 ( 
.A(n_15397),
.B(n_8775),
.Y(n_16438)
);

INVx2_ASAP7_75t_L g16439 ( 
.A(n_15818),
.Y(n_16439)
);

INVx1_ASAP7_75t_L g16440 ( 
.A(n_15298),
.Y(n_16440)
);

AND2x2_ASAP7_75t_L g16441 ( 
.A(n_15636),
.B(n_9406),
.Y(n_16441)
);

HB1xp67_ASAP7_75t_L g16442 ( 
.A(n_15755),
.Y(n_16442)
);

INVx1_ASAP7_75t_L g16443 ( 
.A(n_15355),
.Y(n_16443)
);

INVx2_ASAP7_75t_L g16444 ( 
.A(n_15779),
.Y(n_16444)
);

INVx1_ASAP7_75t_L g16445 ( 
.A(n_15357),
.Y(n_16445)
);

AND2x4_ASAP7_75t_L g16446 ( 
.A(n_15509),
.B(n_8555),
.Y(n_16446)
);

INVx1_ASAP7_75t_L g16447 ( 
.A(n_15757),
.Y(n_16447)
);

INVxp67_ASAP7_75t_L g16448 ( 
.A(n_15743),
.Y(n_16448)
);

NAND2xp5_ASAP7_75t_L g16449 ( 
.A(n_15615),
.B(n_8479),
.Y(n_16449)
);

AND2x2_ASAP7_75t_L g16450 ( 
.A(n_15693),
.B(n_8522),
.Y(n_16450)
);

INVx1_ASAP7_75t_L g16451 ( 
.A(n_15765),
.Y(n_16451)
);

AND2x2_ASAP7_75t_L g16452 ( 
.A(n_15697),
.B(n_15859),
.Y(n_16452)
);

INVx1_ASAP7_75t_L g16453 ( 
.A(n_15389),
.Y(n_16453)
);

INVx1_ASAP7_75t_L g16454 ( 
.A(n_15391),
.Y(n_16454)
);

AND2x4_ASAP7_75t_L g16455 ( 
.A(n_15511),
.B(n_8555),
.Y(n_16455)
);

OR2x2_ASAP7_75t_L g16456 ( 
.A(n_15514),
.B(n_14082),
.Y(n_16456)
);

INVx1_ASAP7_75t_L g16457 ( 
.A(n_15392),
.Y(n_16457)
);

OR2x2_ASAP7_75t_L g16458 ( 
.A(n_15528),
.B(n_9036),
.Y(n_16458)
);

AND2x2_ASAP7_75t_L g16459 ( 
.A(n_15709),
.B(n_8522),
.Y(n_16459)
);

OR2x2_ASAP7_75t_L g16460 ( 
.A(n_15529),
.B(n_9036),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_15813),
.Y(n_16461)
);

AND2x2_ASAP7_75t_L g16462 ( 
.A(n_15576),
.B(n_15823),
.Y(n_16462)
);

NAND2x1p5_ASAP7_75t_L g16463 ( 
.A(n_15536),
.B(n_8232),
.Y(n_16463)
);

AND2x2_ASAP7_75t_L g16464 ( 
.A(n_15839),
.B(n_8522),
.Y(n_16464)
);

AND2x2_ASAP7_75t_L g16465 ( 
.A(n_15781),
.B(n_8578),
.Y(n_16465)
);

XOR2xp5_ASAP7_75t_L g16466 ( 
.A(n_15373),
.B(n_8964),
.Y(n_16466)
);

INVx1_ASAP7_75t_L g16467 ( 
.A(n_15543),
.Y(n_16467)
);

INVx2_ASAP7_75t_L g16468 ( 
.A(n_15806),
.Y(n_16468)
);

AND2x2_ASAP7_75t_L g16469 ( 
.A(n_15804),
.B(n_8578),
.Y(n_16469)
);

INVx2_ASAP7_75t_L g16470 ( 
.A(n_15740),
.Y(n_16470)
);

AND2x2_ASAP7_75t_L g16471 ( 
.A(n_15805),
.B(n_8578),
.Y(n_16471)
);

INVx1_ASAP7_75t_L g16472 ( 
.A(n_15545),
.Y(n_16472)
);

OR2x2_ASAP7_75t_L g16473 ( 
.A(n_15555),
.B(n_9052),
.Y(n_16473)
);

AND2x2_ASAP7_75t_L g16474 ( 
.A(n_15825),
.B(n_15827),
.Y(n_16474)
);

INVx1_ASAP7_75t_L g16475 ( 
.A(n_15561),
.Y(n_16475)
);

NAND2xp5_ASAP7_75t_L g16476 ( 
.A(n_15624),
.B(n_8479),
.Y(n_16476)
);

NAND2xp5_ASAP7_75t_L g16477 ( 
.A(n_15628),
.B(n_8479),
.Y(n_16477)
);

INVx1_ASAP7_75t_L g16478 ( 
.A(n_15574),
.Y(n_16478)
);

INVx1_ASAP7_75t_L g16479 ( 
.A(n_15581),
.Y(n_16479)
);

NOR2xp67_ASAP7_75t_L g16480 ( 
.A(n_15784),
.B(n_11503),
.Y(n_16480)
);

INVx1_ASAP7_75t_L g16481 ( 
.A(n_15600),
.Y(n_16481)
);

AND2x2_ASAP7_75t_L g16482 ( 
.A(n_15208),
.B(n_8588),
.Y(n_16482)
);

OR2x2_ASAP7_75t_L g16483 ( 
.A(n_15632),
.B(n_15660),
.Y(n_16483)
);

OR2x2_ASAP7_75t_L g16484 ( 
.A(n_15643),
.B(n_9052),
.Y(n_16484)
);

OR2x2_ASAP7_75t_L g16485 ( 
.A(n_15645),
.B(n_15646),
.Y(n_16485)
);

AND2x4_ASAP7_75t_L g16486 ( 
.A(n_15607),
.B(n_8573),
.Y(n_16486)
);

NAND2xp5_ASAP7_75t_L g16487 ( 
.A(n_15842),
.B(n_8479),
.Y(n_16487)
);

NAND2x1p5_ASAP7_75t_L g16488 ( 
.A(n_15502),
.B(n_8232),
.Y(n_16488)
);

INVx1_ASAP7_75t_L g16489 ( 
.A(n_15228),
.Y(n_16489)
);

AND2x2_ASAP7_75t_L g16490 ( 
.A(n_15651),
.B(n_15864),
.Y(n_16490)
);

AND2x2_ASAP7_75t_L g16491 ( 
.A(n_15838),
.B(n_15844),
.Y(n_16491)
);

AND2x2_ASAP7_75t_L g16492 ( 
.A(n_15845),
.B(n_8588),
.Y(n_16492)
);

OR2x2_ASAP7_75t_L g16493 ( 
.A(n_15843),
.B(n_9061),
.Y(n_16493)
);

HB1xp67_ASAP7_75t_L g16494 ( 
.A(n_15841),
.Y(n_16494)
);

OR2x2_ASAP7_75t_L g16495 ( 
.A(n_15846),
.B(n_9061),
.Y(n_16495)
);

AND2x4_ASAP7_75t_L g16496 ( 
.A(n_15855),
.B(n_8573),
.Y(n_16496)
);

NAND2xp5_ASAP7_75t_L g16497 ( 
.A(n_15772),
.B(n_8479),
.Y(n_16497)
);

AND2x2_ASAP7_75t_L g16498 ( 
.A(n_15836),
.B(n_8588),
.Y(n_16498)
);

INVx1_ASAP7_75t_L g16499 ( 
.A(n_15237),
.Y(n_16499)
);

NAND2xp5_ASAP7_75t_L g16500 ( 
.A(n_15696),
.B(n_8479),
.Y(n_16500)
);

INVx1_ASAP7_75t_L g16501 ( 
.A(n_15244),
.Y(n_16501)
);

INVx2_ASAP7_75t_L g16502 ( 
.A(n_15868),
.Y(n_16502)
);

OR2x2_ASAP7_75t_L g16503 ( 
.A(n_15710),
.B(n_9091),
.Y(n_16503)
);

INVx2_ASAP7_75t_L g16504 ( 
.A(n_15811),
.Y(n_16504)
);

AND2x2_ASAP7_75t_L g16505 ( 
.A(n_15857),
.B(n_15817),
.Y(n_16505)
);

INVxp67_ASAP7_75t_L g16506 ( 
.A(n_15634),
.Y(n_16506)
);

INVx2_ASAP7_75t_L g16507 ( 
.A(n_15718),
.Y(n_16507)
);

AND2x2_ASAP7_75t_L g16508 ( 
.A(n_15820),
.B(n_8611),
.Y(n_16508)
);

AND2x2_ASAP7_75t_L g16509 ( 
.A(n_15822),
.B(n_15828),
.Y(n_16509)
);

NAND2xp5_ASAP7_75t_L g16510 ( 
.A(n_15758),
.B(n_8479),
.Y(n_16510)
);

INVx1_ASAP7_75t_L g16511 ( 
.A(n_15375),
.Y(n_16511)
);

INVx1_ASAP7_75t_L g16512 ( 
.A(n_15382),
.Y(n_16512)
);

AND2x2_ASAP7_75t_L g16513 ( 
.A(n_15829),
.B(n_8611),
.Y(n_16513)
);

INVx1_ASAP7_75t_L g16514 ( 
.A(n_15318),
.Y(n_16514)
);

AND2x4_ASAP7_75t_L g16515 ( 
.A(n_15847),
.B(n_8573),
.Y(n_16515)
);

INVxp67_ASAP7_75t_L g16516 ( 
.A(n_15849),
.Y(n_16516)
);

INVx1_ASAP7_75t_L g16517 ( 
.A(n_15323),
.Y(n_16517)
);

NAND2xp5_ASAP7_75t_L g16518 ( 
.A(n_15851),
.B(n_8479),
.Y(n_16518)
);

AND2x2_ASAP7_75t_L g16519 ( 
.A(n_15862),
.B(n_8611),
.Y(n_16519)
);

INVx2_ASAP7_75t_L g16520 ( 
.A(n_15720),
.Y(n_16520)
);

INVx1_ASAP7_75t_L g16521 ( 
.A(n_15328),
.Y(n_16521)
);

INVx1_ASAP7_75t_L g16522 ( 
.A(n_15341),
.Y(n_16522)
);

INVx1_ASAP7_75t_L g16523 ( 
.A(n_15342),
.Y(n_16523)
);

NAND4xp25_ASAP7_75t_L g16524 ( 
.A(n_15953),
.B(n_15308),
.C(n_15824),
.D(n_15793),
.Y(n_16524)
);

NOR2x1_ASAP7_75t_L g16525 ( 
.A(n_16187),
.B(n_15361),
.Y(n_16525)
);

AND2x2_ASAP7_75t_L g16526 ( 
.A(n_15982),
.B(n_15730),
.Y(n_16526)
);

AND2x4_ASAP7_75t_L g16527 ( 
.A(n_16385),
.B(n_16011),
.Y(n_16527)
);

INVx1_ASAP7_75t_L g16528 ( 
.A(n_16187),
.Y(n_16528)
);

INVx1_ASAP7_75t_L g16529 ( 
.A(n_15990),
.Y(n_16529)
);

AND2x4_ASAP7_75t_L g16530 ( 
.A(n_15959),
.B(n_15865),
.Y(n_16530)
);

INVx2_ASAP7_75t_L g16531 ( 
.A(n_16022),
.Y(n_16531)
);

INVx1_ASAP7_75t_L g16532 ( 
.A(n_16260),
.Y(n_16532)
);

OR2x2_ASAP7_75t_L g16533 ( 
.A(n_16069),
.B(n_15734),
.Y(n_16533)
);

AND2x2_ASAP7_75t_L g16534 ( 
.A(n_16101),
.B(n_15737),
.Y(n_16534)
);

AND2x2_ASAP7_75t_L g16535 ( 
.A(n_15995),
.B(n_15741),
.Y(n_16535)
);

AND2x2_ASAP7_75t_L g16536 ( 
.A(n_16107),
.B(n_15747),
.Y(n_16536)
);

INVx1_ASAP7_75t_L g16537 ( 
.A(n_16326),
.Y(n_16537)
);

NAND2xp5_ASAP7_75t_L g16538 ( 
.A(n_16326),
.B(n_15752),
.Y(n_16538)
);

AND2x2_ASAP7_75t_L g16539 ( 
.A(n_16282),
.B(n_15754),
.Y(n_16539)
);

AND2x2_ASAP7_75t_L g16540 ( 
.A(n_16256),
.B(n_15669),
.Y(n_16540)
);

INVx1_ASAP7_75t_L g16541 ( 
.A(n_16404),
.Y(n_16541)
);

AND2x2_ASAP7_75t_L g16542 ( 
.A(n_16256),
.B(n_15670),
.Y(n_16542)
);

INVx2_ASAP7_75t_SL g16543 ( 
.A(n_16336),
.Y(n_16543)
);

INVxp67_ASAP7_75t_L g16544 ( 
.A(n_16250),
.Y(n_16544)
);

INVx2_ASAP7_75t_L g16545 ( 
.A(n_16265),
.Y(n_16545)
);

INVx2_ASAP7_75t_L g16546 ( 
.A(n_16265),
.Y(n_16546)
);

OR2x2_ASAP7_75t_L g16547 ( 
.A(n_15883),
.B(n_15672),
.Y(n_16547)
);

AND2x2_ASAP7_75t_L g16548 ( 
.A(n_16176),
.B(n_15677),
.Y(n_16548)
);

NAND2xp5_ASAP7_75t_L g16549 ( 
.A(n_16236),
.B(n_15678),
.Y(n_16549)
);

INVx1_ASAP7_75t_L g16550 ( 
.A(n_16404),
.Y(n_16550)
);

NOR4xp25_ASAP7_75t_SL g16551 ( 
.A(n_16054),
.B(n_15707),
.C(n_15277),
.D(n_15288),
.Y(n_16551)
);

NAND2xp5_ASAP7_75t_L g16552 ( 
.A(n_16402),
.B(n_15681),
.Y(n_16552)
);

AND2x2_ASAP7_75t_L g16553 ( 
.A(n_16296),
.B(n_15695),
.Y(n_16553)
);

OR2x2_ASAP7_75t_L g16554 ( 
.A(n_16130),
.B(n_15702),
.Y(n_16554)
);

INVx2_ASAP7_75t_L g16555 ( 
.A(n_15927),
.Y(n_16555)
);

INVx2_ASAP7_75t_L g16556 ( 
.A(n_15934),
.Y(n_16556)
);

INVx1_ASAP7_75t_L g16557 ( 
.A(n_16105),
.Y(n_16557)
);

INVx1_ASAP7_75t_L g16558 ( 
.A(n_16057),
.Y(n_16558)
);

NAND2xp5_ASAP7_75t_SL g16559 ( 
.A(n_16402),
.B(n_15854),
.Y(n_16559)
);

INVx1_ASAP7_75t_SL g16560 ( 
.A(n_16401),
.Y(n_16560)
);

AND2x2_ASAP7_75t_L g16561 ( 
.A(n_16118),
.B(n_15708),
.Y(n_16561)
);

AND2x2_ASAP7_75t_L g16562 ( 
.A(n_16102),
.B(n_15773),
.Y(n_16562)
);

AND2x2_ASAP7_75t_L g16563 ( 
.A(n_16474),
.B(n_15780),
.Y(n_16563)
);

INVx1_ASAP7_75t_L g16564 ( 
.A(n_16057),
.Y(n_16564)
);

AND2x2_ASAP7_75t_L g16565 ( 
.A(n_15893),
.B(n_15790),
.Y(n_16565)
);

INVx2_ASAP7_75t_L g16566 ( 
.A(n_16338),
.Y(n_16566)
);

INVx1_ASAP7_75t_L g16567 ( 
.A(n_16288),
.Y(n_16567)
);

AND2x2_ASAP7_75t_L g16568 ( 
.A(n_16015),
.B(n_15794),
.Y(n_16568)
);

AND2x2_ASAP7_75t_L g16569 ( 
.A(n_15897),
.B(n_15795),
.Y(n_16569)
);

AND2x2_ASAP7_75t_L g16570 ( 
.A(n_16208),
.B(n_15800),
.Y(n_16570)
);

INVxp67_ASAP7_75t_L g16571 ( 
.A(n_16185),
.Y(n_16571)
);

AND2x2_ASAP7_75t_L g16572 ( 
.A(n_15879),
.B(n_15808),
.Y(n_16572)
);

AND2x2_ASAP7_75t_L g16573 ( 
.A(n_16016),
.B(n_15515),
.Y(n_16573)
);

HB1xp67_ASAP7_75t_L g16574 ( 
.A(n_16161),
.Y(n_16574)
);

INVx1_ASAP7_75t_SL g16575 ( 
.A(n_16038),
.Y(n_16575)
);

INVx2_ASAP7_75t_L g16576 ( 
.A(n_16338),
.Y(n_16576)
);

NAND2xp5_ASAP7_75t_L g16577 ( 
.A(n_16098),
.B(n_15281),
.Y(n_16577)
);

NAND2xp5_ASAP7_75t_L g16578 ( 
.A(n_15983),
.B(n_15370),
.Y(n_16578)
);

NAND2xp5_ASAP7_75t_L g16579 ( 
.A(n_15984),
.B(n_15521),
.Y(n_16579)
);

INVx1_ASAP7_75t_L g16580 ( 
.A(n_16307),
.Y(n_16580)
);

INVx1_ASAP7_75t_L g16581 ( 
.A(n_16199),
.Y(n_16581)
);

INVx1_ASAP7_75t_L g16582 ( 
.A(n_16150),
.Y(n_16582)
);

AND2x2_ASAP7_75t_L g16583 ( 
.A(n_15974),
.B(n_15522),
.Y(n_16583)
);

HB1xp67_ASAP7_75t_L g16584 ( 
.A(n_16267),
.Y(n_16584)
);

INVx4_ASAP7_75t_L g16585 ( 
.A(n_16227),
.Y(n_16585)
);

INVx2_ASAP7_75t_L g16586 ( 
.A(n_16390),
.Y(n_16586)
);

NAND2xp5_ASAP7_75t_L g16587 ( 
.A(n_15964),
.B(n_15532),
.Y(n_16587)
);

AND2x4_ASAP7_75t_L g16588 ( 
.A(n_16221),
.B(n_15534),
.Y(n_16588)
);

NAND2xp5_ASAP7_75t_L g16589 ( 
.A(n_15914),
.B(n_15535),
.Y(n_16589)
);

INVx1_ASAP7_75t_L g16590 ( 
.A(n_16341),
.Y(n_16590)
);

OR2x2_ASAP7_75t_L g16591 ( 
.A(n_15874),
.B(n_15538),
.Y(n_16591)
);

INVx2_ASAP7_75t_L g16592 ( 
.A(n_16002),
.Y(n_16592)
);

INVx1_ASAP7_75t_L g16593 ( 
.A(n_15985),
.Y(n_16593)
);

INVx3_ASAP7_75t_L g16594 ( 
.A(n_15931),
.Y(n_16594)
);

NAND2xp5_ASAP7_75t_L g16595 ( 
.A(n_15909),
.B(n_15539),
.Y(n_16595)
);

NOR2xp33_ASAP7_75t_L g16596 ( 
.A(n_16122),
.B(n_15396),
.Y(n_16596)
);

INVx1_ASAP7_75t_L g16597 ( 
.A(n_16167),
.Y(n_16597)
);

BUFx2_ASAP7_75t_L g16598 ( 
.A(n_15988),
.Y(n_16598)
);

OR2x2_ASAP7_75t_L g16599 ( 
.A(n_15908),
.B(n_15541),
.Y(n_16599)
);

INVx3_ASAP7_75t_L g16600 ( 
.A(n_16000),
.Y(n_16600)
);

AOI21xp5_ASAP7_75t_L g16601 ( 
.A1(n_16292),
.A2(n_15644),
.B(n_15597),
.Y(n_16601)
);

OR2x2_ASAP7_75t_L g16602 ( 
.A(n_15877),
.B(n_15549),
.Y(n_16602)
);

AND2x2_ASAP7_75t_L g16603 ( 
.A(n_16030),
.B(n_15554),
.Y(n_16603)
);

AND2x2_ASAP7_75t_L g16604 ( 
.A(n_15910),
.B(n_15559),
.Y(n_16604)
);

AND2x4_ASAP7_75t_L g16605 ( 
.A(n_16233),
.B(n_15568),
.Y(n_16605)
);

INVx1_ASAP7_75t_L g16606 ( 
.A(n_16174),
.Y(n_16606)
);

NAND2xp5_ASAP7_75t_L g16607 ( 
.A(n_16505),
.B(n_15569),
.Y(n_16607)
);

AND2x2_ASAP7_75t_L g16608 ( 
.A(n_15888),
.B(n_15575),
.Y(n_16608)
);

AOI22xp33_ASAP7_75t_L g16609 ( 
.A1(n_15967),
.A2(n_15198),
.B1(n_15657),
.B2(n_15852),
.Y(n_16609)
);

OR2x2_ASAP7_75t_L g16610 ( 
.A(n_15944),
.B(n_15578),
.Y(n_16610)
);

OR2x2_ASAP7_75t_L g16611 ( 
.A(n_15957),
.B(n_15580),
.Y(n_16611)
);

INVx1_ASAP7_75t_L g16612 ( 
.A(n_16229),
.Y(n_16612)
);

AND2x2_ASAP7_75t_L g16613 ( 
.A(n_16303),
.B(n_15584),
.Y(n_16613)
);

NOR2x1_ASAP7_75t_L g16614 ( 
.A(n_16212),
.B(n_15366),
.Y(n_16614)
);

INVx2_ASAP7_75t_L g16615 ( 
.A(n_16269),
.Y(n_16615)
);

INVxp67_ASAP7_75t_SL g16616 ( 
.A(n_15886),
.Y(n_16616)
);

INVx1_ASAP7_75t_L g16617 ( 
.A(n_15942),
.Y(n_16617)
);

NAND2xp5_ASAP7_75t_L g16618 ( 
.A(n_15965),
.B(n_15586),
.Y(n_16618)
);

AND2x2_ASAP7_75t_L g16619 ( 
.A(n_16304),
.B(n_15592),
.Y(n_16619)
);

NAND2xp5_ASAP7_75t_L g16620 ( 
.A(n_16406),
.B(n_15598),
.Y(n_16620)
);

INVx1_ASAP7_75t_L g16621 ( 
.A(n_16434),
.Y(n_16621)
);

AND2x2_ASAP7_75t_L g16622 ( 
.A(n_16008),
.B(n_15604),
.Y(n_16622)
);

AND2x2_ASAP7_75t_L g16623 ( 
.A(n_16003),
.B(n_15343),
.Y(n_16623)
);

NAND2xp5_ASAP7_75t_L g16624 ( 
.A(n_16381),
.B(n_15777),
.Y(n_16624)
);

INVx2_ASAP7_75t_L g16625 ( 
.A(n_16269),
.Y(n_16625)
);

INVx2_ASAP7_75t_L g16626 ( 
.A(n_16491),
.Y(n_16626)
);

AND2x2_ASAP7_75t_L g16627 ( 
.A(n_15998),
.B(n_15344),
.Y(n_16627)
);

AND2x4_ASAP7_75t_SL g16628 ( 
.A(n_15905),
.B(n_15346),
.Y(n_16628)
);

AND2x2_ASAP7_75t_L g16629 ( 
.A(n_15930),
.B(n_15896),
.Y(n_16629)
);

AND2x4_ASAP7_75t_L g16630 ( 
.A(n_15875),
.B(n_15348),
.Y(n_16630)
);

NAND2xp5_ASAP7_75t_L g16631 ( 
.A(n_16382),
.B(n_15821),
.Y(n_16631)
);

INVx1_ASAP7_75t_L g16632 ( 
.A(n_15972),
.Y(n_16632)
);

INVx1_ASAP7_75t_L g16633 ( 
.A(n_15924),
.Y(n_16633)
);

AND2x4_ASAP7_75t_L g16634 ( 
.A(n_16140),
.B(n_15837),
.Y(n_16634)
);

NOR2xp67_ASAP7_75t_L g16635 ( 
.A(n_16379),
.B(n_15867),
.Y(n_16635)
);

INVx4_ASAP7_75t_SL g16636 ( 
.A(n_15880),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_15949),
.Y(n_16637)
);

NOR2x1_ASAP7_75t_L g16638 ( 
.A(n_15946),
.B(n_15776),
.Y(n_16638)
);

AND2x2_ASAP7_75t_L g16639 ( 
.A(n_15938),
.B(n_15440),
.Y(n_16639)
);

INVx1_ASAP7_75t_L g16640 ( 
.A(n_15987),
.Y(n_16640)
);

AND2x2_ASAP7_75t_L g16641 ( 
.A(n_15945),
.B(n_16352),
.Y(n_16641)
);

NOR2xp33_ASAP7_75t_SL g16642 ( 
.A(n_16036),
.B(n_8260),
.Y(n_16642)
);

INVx1_ASAP7_75t_L g16643 ( 
.A(n_15882),
.Y(n_16643)
);

INVx2_ASAP7_75t_L g16644 ( 
.A(n_15870),
.Y(n_16644)
);

OR2x2_ASAP7_75t_L g16645 ( 
.A(n_15975),
.B(n_15378),
.Y(n_16645)
);

AND2x2_ASAP7_75t_L g16646 ( 
.A(n_16462),
.B(n_15221),
.Y(n_16646)
);

AND2x2_ASAP7_75t_L g16647 ( 
.A(n_15991),
.B(n_15236),
.Y(n_16647)
);

INVx1_ASAP7_75t_L g16648 ( 
.A(n_15891),
.Y(n_16648)
);

NOR2xp33_ASAP7_75t_L g16649 ( 
.A(n_15936),
.B(n_11271),
.Y(n_16649)
);

AND2x2_ASAP7_75t_L g16650 ( 
.A(n_15907),
.B(n_11271),
.Y(n_16650)
);

AND2x2_ASAP7_75t_L g16651 ( 
.A(n_15890),
.B(n_11277),
.Y(n_16651)
);

INVx2_ASAP7_75t_L g16652 ( 
.A(n_16180),
.Y(n_16652)
);

INVx2_ASAP7_75t_L g16653 ( 
.A(n_16186),
.Y(n_16653)
);

OR2x2_ASAP7_75t_L g16654 ( 
.A(n_15980),
.B(n_15962),
.Y(n_16654)
);

NAND2xp5_ASAP7_75t_L g16655 ( 
.A(n_16333),
.B(n_8505),
.Y(n_16655)
);

AND2x2_ASAP7_75t_L g16656 ( 
.A(n_15900),
.B(n_11277),
.Y(n_16656)
);

INVx1_ASAP7_75t_L g16657 ( 
.A(n_15901),
.Y(n_16657)
);

AND2x2_ASAP7_75t_L g16658 ( 
.A(n_16172),
.B(n_11286),
.Y(n_16658)
);

AND2x2_ASAP7_75t_L g16659 ( 
.A(n_16007),
.B(n_11286),
.Y(n_16659)
);

BUFx4f_ASAP7_75t_L g16660 ( 
.A(n_15906),
.Y(n_16660)
);

AND2x2_ASAP7_75t_L g16661 ( 
.A(n_15977),
.B(n_11290),
.Y(n_16661)
);

INVx1_ASAP7_75t_L g16662 ( 
.A(n_16032),
.Y(n_16662)
);

AND2x2_ASAP7_75t_L g16663 ( 
.A(n_16005),
.B(n_11290),
.Y(n_16663)
);

INVx1_ASAP7_75t_L g16664 ( 
.A(n_15894),
.Y(n_16664)
);

INVx1_ASAP7_75t_L g16665 ( 
.A(n_16004),
.Y(n_16665)
);

OR2x2_ASAP7_75t_L g16666 ( 
.A(n_15918),
.B(n_11294),
.Y(n_16666)
);

AND2x4_ASAP7_75t_L g16667 ( 
.A(n_16068),
.B(n_8626),
.Y(n_16667)
);

INVx2_ASAP7_75t_L g16668 ( 
.A(n_16183),
.Y(n_16668)
);

AND2x2_ASAP7_75t_L g16669 ( 
.A(n_16376),
.B(n_11294),
.Y(n_16669)
);

INVx1_ASAP7_75t_L g16670 ( 
.A(n_16010),
.Y(n_16670)
);

HB1xp67_ASAP7_75t_L g16671 ( 
.A(n_16358),
.Y(n_16671)
);

INVx2_ASAP7_75t_L g16672 ( 
.A(n_16243),
.Y(n_16672)
);

INVx4_ASAP7_75t_L g16673 ( 
.A(n_15932),
.Y(n_16673)
);

NAND2xp5_ASAP7_75t_L g16674 ( 
.A(n_16131),
.B(n_8505),
.Y(n_16674)
);

HB1xp67_ASAP7_75t_L g16675 ( 
.A(n_16188),
.Y(n_16675)
);

BUFx2_ASAP7_75t_L g16676 ( 
.A(n_15872),
.Y(n_16676)
);

OR2x2_ASAP7_75t_L g16677 ( 
.A(n_16048),
.B(n_11299),
.Y(n_16677)
);

HB1xp67_ASAP7_75t_L g16678 ( 
.A(n_16062),
.Y(n_16678)
);

AND2x2_ASAP7_75t_L g16679 ( 
.A(n_16121),
.B(n_11299),
.Y(n_16679)
);

AND2x4_ASAP7_75t_SL g16680 ( 
.A(n_16164),
.B(n_7076),
.Y(n_16680)
);

AND2x2_ASAP7_75t_L g16681 ( 
.A(n_15903),
.B(n_11300),
.Y(n_16681)
);

HB1xp67_ASAP7_75t_L g16682 ( 
.A(n_16415),
.Y(n_16682)
);

AND2x2_ASAP7_75t_L g16683 ( 
.A(n_15904),
.B(n_11300),
.Y(n_16683)
);

INVx1_ASAP7_75t_L g16684 ( 
.A(n_15887),
.Y(n_16684)
);

INVx1_ASAP7_75t_SL g16685 ( 
.A(n_16064),
.Y(n_16685)
);

INVx1_ASAP7_75t_L g16686 ( 
.A(n_16494),
.Y(n_16686)
);

OR2x2_ASAP7_75t_L g16687 ( 
.A(n_15940),
.B(n_11301),
.Y(n_16687)
);

INVx1_ASAP7_75t_L g16688 ( 
.A(n_15943),
.Y(n_16688)
);

NOR2xp67_ASAP7_75t_L g16689 ( 
.A(n_16316),
.B(n_11510),
.Y(n_16689)
);

INVx1_ASAP7_75t_L g16690 ( 
.A(n_15948),
.Y(n_16690)
);

INVxp67_ASAP7_75t_L g16691 ( 
.A(n_16050),
.Y(n_16691)
);

OR2x2_ASAP7_75t_L g16692 ( 
.A(n_15895),
.B(n_11301),
.Y(n_16692)
);

OR2x2_ASAP7_75t_L g16693 ( 
.A(n_15960),
.B(n_11302),
.Y(n_16693)
);

INVx1_ASAP7_75t_L g16694 ( 
.A(n_15933),
.Y(n_16694)
);

AND2x2_ASAP7_75t_L g16695 ( 
.A(n_15884),
.B(n_11302),
.Y(n_16695)
);

AOI22xp33_ASAP7_75t_L g16696 ( 
.A1(n_15881),
.A2(n_11523),
.B1(n_11527),
.B2(n_11522),
.Y(n_16696)
);

OAI22xp5_ASAP7_75t_L g16697 ( 
.A1(n_15969),
.A2(n_11308),
.B1(n_11310),
.B2(n_11307),
.Y(n_16697)
);

BUFx2_ASAP7_75t_L g16698 ( 
.A(n_15951),
.Y(n_16698)
);

AND2x2_ASAP7_75t_L g16699 ( 
.A(n_15885),
.B(n_11307),
.Y(n_16699)
);

AND2x4_ASAP7_75t_L g16700 ( 
.A(n_15997),
.B(n_16129),
.Y(n_16700)
);

AND2x2_ASAP7_75t_L g16701 ( 
.A(n_16452),
.B(n_16490),
.Y(n_16701)
);

AOI22xp33_ASAP7_75t_SL g16702 ( 
.A1(n_16014),
.A2(n_11523),
.B1(n_11527),
.B2(n_11522),
.Y(n_16702)
);

INVx1_ASAP7_75t_L g16703 ( 
.A(n_15935),
.Y(n_16703)
);

HB1xp67_ASAP7_75t_L g16704 ( 
.A(n_16480),
.Y(n_16704)
);

OR2x2_ASAP7_75t_L g16705 ( 
.A(n_16080),
.B(n_16191),
.Y(n_16705)
);

INVx2_ASAP7_75t_SL g16706 ( 
.A(n_15899),
.Y(n_16706)
);

AND2x2_ASAP7_75t_L g16707 ( 
.A(n_16226),
.B(n_11308),
.Y(n_16707)
);

INVx2_ASAP7_75t_SL g16708 ( 
.A(n_16371),
.Y(n_16708)
);

AND2x2_ASAP7_75t_L g16709 ( 
.A(n_16023),
.B(n_16046),
.Y(n_16709)
);

INVx2_ASAP7_75t_L g16710 ( 
.A(n_16035),
.Y(n_16710)
);

AND2x4_ASAP7_75t_L g16711 ( 
.A(n_16132),
.B(n_8626),
.Y(n_16711)
);

BUFx4f_ASAP7_75t_SL g16712 ( 
.A(n_16165),
.Y(n_16712)
);

AND2x2_ASAP7_75t_L g16713 ( 
.A(n_16031),
.B(n_11310),
.Y(n_16713)
);

INVx1_ASAP7_75t_L g16714 ( 
.A(n_15947),
.Y(n_16714)
);

AND2x2_ASAP7_75t_L g16715 ( 
.A(n_16009),
.B(n_11311),
.Y(n_16715)
);

NAND2xp5_ASAP7_75t_L g16716 ( 
.A(n_16332),
.B(n_8505),
.Y(n_16716)
);

INVx3_ASAP7_75t_L g16717 ( 
.A(n_15954),
.Y(n_16717)
);

INVx2_ASAP7_75t_L g16718 ( 
.A(n_16040),
.Y(n_16718)
);

OR2x6_ASAP7_75t_L g16719 ( 
.A(n_16157),
.B(n_10424),
.Y(n_16719)
);

INVx3_ASAP7_75t_L g16720 ( 
.A(n_15963),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_15950),
.Y(n_16721)
);

AND2x2_ASAP7_75t_L g16722 ( 
.A(n_16042),
.B(n_11311),
.Y(n_16722)
);

INVx4_ASAP7_75t_L g16723 ( 
.A(n_16368),
.Y(n_16723)
);

INVxp67_ASAP7_75t_L g16724 ( 
.A(n_15999),
.Y(n_16724)
);

INVx1_ASAP7_75t_L g16725 ( 
.A(n_15958),
.Y(n_16725)
);

OR2x2_ASAP7_75t_L g16726 ( 
.A(n_15915),
.B(n_15917),
.Y(n_16726)
);

AOI21xp5_ASAP7_75t_L g16727 ( 
.A1(n_16013),
.A2(n_16448),
.B(n_16151),
.Y(n_16727)
);

NAND2xp5_ASAP7_75t_L g16728 ( 
.A(n_16334),
.B(n_8505),
.Y(n_16728)
);

AND2x4_ASAP7_75t_SL g16729 ( 
.A(n_16435),
.B(n_7076),
.Y(n_16729)
);

AND2x2_ASAP7_75t_L g16730 ( 
.A(n_16043),
.B(n_11315),
.Y(n_16730)
);

NAND2xp5_ASAP7_75t_L g16731 ( 
.A(n_16225),
.B(n_8505),
.Y(n_16731)
);

INVx2_ASAP7_75t_L g16732 ( 
.A(n_16018),
.Y(n_16732)
);

INVx2_ASAP7_75t_L g16733 ( 
.A(n_16021),
.Y(n_16733)
);

HB1xp67_ASAP7_75t_L g16734 ( 
.A(n_16128),
.Y(n_16734)
);

HB1xp67_ASAP7_75t_L g16735 ( 
.A(n_16189),
.Y(n_16735)
);

AND2x2_ASAP7_75t_L g16736 ( 
.A(n_16052),
.B(n_11315),
.Y(n_16736)
);

AND2x2_ASAP7_75t_L g16737 ( 
.A(n_16067),
.B(n_11316),
.Y(n_16737)
);

INVx1_ASAP7_75t_L g16738 ( 
.A(n_15968),
.Y(n_16738)
);

INVx1_ASAP7_75t_L g16739 ( 
.A(n_15973),
.Y(n_16739)
);

AND2x2_ASAP7_75t_L g16740 ( 
.A(n_16136),
.B(n_16141),
.Y(n_16740)
);

INVx1_ASAP7_75t_L g16741 ( 
.A(n_15986),
.Y(n_16741)
);

INVx2_ASAP7_75t_SL g16742 ( 
.A(n_16254),
.Y(n_16742)
);

INVx1_ASAP7_75t_SL g16743 ( 
.A(n_16037),
.Y(n_16743)
);

AND2x2_ASAP7_75t_L g16744 ( 
.A(n_16149),
.B(n_11316),
.Y(n_16744)
);

INVx1_ASAP7_75t_L g16745 ( 
.A(n_15989),
.Y(n_16745)
);

AND2x2_ASAP7_75t_L g16746 ( 
.A(n_16160),
.B(n_11318),
.Y(n_16746)
);

AND2x2_ASAP7_75t_L g16747 ( 
.A(n_16083),
.B(n_11318),
.Y(n_16747)
);

AND2x2_ASAP7_75t_L g16748 ( 
.A(n_16439),
.B(n_11321),
.Y(n_16748)
);

AND2x2_ASAP7_75t_L g16749 ( 
.A(n_16444),
.B(n_11321),
.Y(n_16749)
);

AND2x2_ASAP7_75t_L g16750 ( 
.A(n_16468),
.B(n_11322),
.Y(n_16750)
);

INVx1_ASAP7_75t_L g16751 ( 
.A(n_15955),
.Y(n_16751)
);

NAND2xp5_ASAP7_75t_L g16752 ( 
.A(n_16470),
.B(n_8505),
.Y(n_16752)
);

NAND2xp5_ASAP7_75t_L g16753 ( 
.A(n_16337),
.B(n_8505),
.Y(n_16753)
);

NAND2xp5_ASAP7_75t_L g16754 ( 
.A(n_16343),
.B(n_8505),
.Y(n_16754)
);

INVx2_ASAP7_75t_L g16755 ( 
.A(n_16459),
.Y(n_16755)
);

INVx2_ASAP7_75t_L g16756 ( 
.A(n_16196),
.Y(n_16756)
);

AND2x2_ASAP7_75t_L g16757 ( 
.A(n_16367),
.B(n_11322),
.Y(n_16757)
);

AND2x2_ASAP7_75t_L g16758 ( 
.A(n_15926),
.B(n_11328),
.Y(n_16758)
);

AND2x4_ASAP7_75t_L g16759 ( 
.A(n_16396),
.B(n_8626),
.Y(n_16759)
);

NAND2xp5_ASAP7_75t_L g16760 ( 
.A(n_16271),
.B(n_11328),
.Y(n_16760)
);

OR2x2_ASAP7_75t_L g16761 ( 
.A(n_15956),
.B(n_11337),
.Y(n_16761)
);

AND2x2_ASAP7_75t_L g16762 ( 
.A(n_15978),
.B(n_11337),
.Y(n_16762)
);

AND2x2_ASAP7_75t_L g16763 ( 
.A(n_15979),
.B(n_11338),
.Y(n_16763)
);

INVxp67_ASAP7_75t_L g16764 ( 
.A(n_16049),
.Y(n_16764)
);

AND2x2_ASAP7_75t_L g16765 ( 
.A(n_16363),
.B(n_11338),
.Y(n_16765)
);

AND2x2_ASAP7_75t_L g16766 ( 
.A(n_16261),
.B(n_11341),
.Y(n_16766)
);

INVxp67_ASAP7_75t_L g16767 ( 
.A(n_16425),
.Y(n_16767)
);

INVx1_ASAP7_75t_SL g16768 ( 
.A(n_15971),
.Y(n_16768)
);

INVx1_ASAP7_75t_L g16769 ( 
.A(n_16100),
.Y(n_16769)
);

INVx4_ASAP7_75t_L g16770 ( 
.A(n_15889),
.Y(n_16770)
);

NAND2xp5_ASAP7_75t_L g16771 ( 
.A(n_16272),
.B(n_11341),
.Y(n_16771)
);

AND2x4_ASAP7_75t_L g16772 ( 
.A(n_16086),
.B(n_8654),
.Y(n_16772)
);

OR2x2_ASAP7_75t_L g16773 ( 
.A(n_16114),
.B(n_11344),
.Y(n_16773)
);

OR2x2_ASAP7_75t_L g16774 ( 
.A(n_16125),
.B(n_11344),
.Y(n_16774)
);

INVx2_ASAP7_75t_SL g16775 ( 
.A(n_16399),
.Y(n_16775)
);

OR2x2_ASAP7_75t_L g16776 ( 
.A(n_16087),
.B(n_11345),
.Y(n_16776)
);

INVx1_ASAP7_75t_L g16777 ( 
.A(n_15939),
.Y(n_16777)
);

INVx1_ASAP7_75t_L g16778 ( 
.A(n_15941),
.Y(n_16778)
);

AND2x2_ASAP7_75t_L g16779 ( 
.A(n_16108),
.B(n_11345),
.Y(n_16779)
);

INVx1_ASAP7_75t_L g16780 ( 
.A(n_15922),
.Y(n_16780)
);

INVxp67_ASAP7_75t_SL g16781 ( 
.A(n_16148),
.Y(n_16781)
);

AND2x2_ASAP7_75t_L g16782 ( 
.A(n_16109),
.B(n_11347),
.Y(n_16782)
);

BUFx2_ASAP7_75t_L g16783 ( 
.A(n_16456),
.Y(n_16783)
);

AND2x2_ASAP7_75t_L g16784 ( 
.A(n_16113),
.B(n_11347),
.Y(n_16784)
);

AND2x2_ASAP7_75t_L g16785 ( 
.A(n_16502),
.B(n_11353),
.Y(n_16785)
);

NAND2xp5_ASAP7_75t_SL g16786 ( 
.A(n_16039),
.B(n_10538),
.Y(n_16786)
);

AND2x2_ASAP7_75t_L g16787 ( 
.A(n_16285),
.B(n_11353),
.Y(n_16787)
);

AND2x2_ASAP7_75t_L g16788 ( 
.A(n_16244),
.B(n_16066),
.Y(n_16788)
);

NAND2xp33_ASAP7_75t_SL g16789 ( 
.A(n_16431),
.B(n_15912),
.Y(n_16789)
);

INVx3_ASAP7_75t_L g16790 ( 
.A(n_16146),
.Y(n_16790)
);

BUFx3_ASAP7_75t_L g16791 ( 
.A(n_16089),
.Y(n_16791)
);

AND2x2_ASAP7_75t_L g16792 ( 
.A(n_16301),
.B(n_11369),
.Y(n_16792)
);

AND2x4_ASAP7_75t_L g16793 ( 
.A(n_16392),
.B(n_8654),
.Y(n_16793)
);

NAND2xp5_ASAP7_75t_L g16794 ( 
.A(n_16273),
.B(n_11369),
.Y(n_16794)
);

INVx1_ASAP7_75t_L g16795 ( 
.A(n_15937),
.Y(n_16795)
);

NAND2xp5_ASAP7_75t_L g16796 ( 
.A(n_16274),
.B(n_16214),
.Y(n_16796)
);

INVx1_ASAP7_75t_SL g16797 ( 
.A(n_16075),
.Y(n_16797)
);

OR2x2_ASAP7_75t_L g16798 ( 
.A(n_16096),
.B(n_11370),
.Y(n_16798)
);

NAND2xp5_ASAP7_75t_L g16799 ( 
.A(n_16228),
.B(n_11370),
.Y(n_16799)
);

INVx2_ASAP7_75t_L g16800 ( 
.A(n_16202),
.Y(n_16800)
);

NAND2xp5_ASAP7_75t_L g16801 ( 
.A(n_16280),
.B(n_11385),
.Y(n_16801)
);

AND2x2_ASAP7_75t_L g16802 ( 
.A(n_16090),
.B(n_11385),
.Y(n_16802)
);

NAND2xp5_ASAP7_75t_L g16803 ( 
.A(n_16092),
.B(n_11388),
.Y(n_16803)
);

AND2x2_ASAP7_75t_L g16804 ( 
.A(n_16097),
.B(n_11388),
.Y(n_16804)
);

NAND2xp5_ASAP7_75t_L g16805 ( 
.A(n_16088),
.B(n_16241),
.Y(n_16805)
);

AND2x2_ASAP7_75t_L g16806 ( 
.A(n_16409),
.B(n_11393),
.Y(n_16806)
);

INVx1_ASAP7_75t_L g16807 ( 
.A(n_15928),
.Y(n_16807)
);

OR2x2_ASAP7_75t_L g16808 ( 
.A(n_16152),
.B(n_11393),
.Y(n_16808)
);

AND2x2_ASAP7_75t_L g16809 ( 
.A(n_16275),
.B(n_11398),
.Y(n_16809)
);

HB1xp67_ASAP7_75t_L g16810 ( 
.A(n_16442),
.Y(n_16810)
);

AND2x2_ASAP7_75t_L g16811 ( 
.A(n_16275),
.B(n_11398),
.Y(n_16811)
);

INVx2_ASAP7_75t_L g16812 ( 
.A(n_16224),
.Y(n_16812)
);

OR2x6_ASAP7_75t_L g16813 ( 
.A(n_16026),
.B(n_10424),
.Y(n_16813)
);

NAND2xp5_ASAP7_75t_L g16814 ( 
.A(n_16159),
.B(n_11400),
.Y(n_16814)
);

AND2x2_ASAP7_75t_L g16815 ( 
.A(n_16056),
.B(n_11400),
.Y(n_16815)
);

AND2x2_ASAP7_75t_L g16816 ( 
.A(n_16429),
.B(n_11404),
.Y(n_16816)
);

INVx1_ASAP7_75t_L g16817 ( 
.A(n_15929),
.Y(n_16817)
);

INVx1_ASAP7_75t_L g16818 ( 
.A(n_16153),
.Y(n_16818)
);

HB1xp67_ASAP7_75t_L g16819 ( 
.A(n_16155),
.Y(n_16819)
);

OR2x2_ASAP7_75t_L g16820 ( 
.A(n_16163),
.B(n_11404),
.Y(n_16820)
);

NAND2xp5_ASAP7_75t_L g16821 ( 
.A(n_16179),
.B(n_11413),
.Y(n_16821)
);

AND2x2_ASAP7_75t_L g16822 ( 
.A(n_16184),
.B(n_11413),
.Y(n_16822)
);

BUFx2_ASAP7_75t_L g16823 ( 
.A(n_16123),
.Y(n_16823)
);

INVx1_ASAP7_75t_L g16824 ( 
.A(n_16166),
.Y(n_16824)
);

NAND2xp5_ASAP7_75t_L g16825 ( 
.A(n_15952),
.B(n_11415),
.Y(n_16825)
);

NAND2xp5_ASAP7_75t_L g16826 ( 
.A(n_16347),
.B(n_11415),
.Y(n_16826)
);

OR2x2_ASAP7_75t_L g16827 ( 
.A(n_16170),
.B(n_11420),
.Y(n_16827)
);

INVx1_ASAP7_75t_SL g16828 ( 
.A(n_16156),
.Y(n_16828)
);

INVx1_ASAP7_75t_L g16829 ( 
.A(n_16173),
.Y(n_16829)
);

INVx5_ASAP7_75t_L g16830 ( 
.A(n_15976),
.Y(n_16830)
);

INVx1_ASAP7_75t_L g16831 ( 
.A(n_16278),
.Y(n_16831)
);

INVx2_ASAP7_75t_L g16832 ( 
.A(n_16369),
.Y(n_16832)
);

OR2x2_ASAP7_75t_L g16833 ( 
.A(n_16139),
.B(n_11420),
.Y(n_16833)
);

NOR2x1_ASAP7_75t_L g16834 ( 
.A(n_16178),
.B(n_11534),
.Y(n_16834)
);

AND2x2_ASAP7_75t_L g16835 ( 
.A(n_16084),
.B(n_16025),
.Y(n_16835)
);

AND2x2_ASAP7_75t_L g16836 ( 
.A(n_16065),
.B(n_16024),
.Y(n_16836)
);

NAND2xp5_ASAP7_75t_L g16837 ( 
.A(n_16218),
.B(n_11423),
.Y(n_16837)
);

AND2x4_ASAP7_75t_L g16838 ( 
.A(n_16373),
.B(n_8654),
.Y(n_16838)
);

AND2x2_ASAP7_75t_L g16839 ( 
.A(n_16028),
.B(n_11423),
.Y(n_16839)
);

AND2x2_ASAP7_75t_L g16840 ( 
.A(n_16029),
.B(n_11424),
.Y(n_16840)
);

NAND2xp5_ASAP7_75t_L g16841 ( 
.A(n_16249),
.B(n_11424),
.Y(n_16841)
);

INVx2_ASAP7_75t_L g16842 ( 
.A(n_16111),
.Y(n_16842)
);

INVx1_ASAP7_75t_L g16843 ( 
.A(n_16095),
.Y(n_16843)
);

INVx1_ASAP7_75t_L g16844 ( 
.A(n_16119),
.Y(n_16844)
);

INVx1_ASAP7_75t_SL g16845 ( 
.A(n_16158),
.Y(n_16845)
);

NAND2xp5_ASAP7_75t_L g16846 ( 
.A(n_16210),
.B(n_11430),
.Y(n_16846)
);

AND2x2_ASAP7_75t_L g16847 ( 
.A(n_16315),
.B(n_11430),
.Y(n_16847)
);

INVx2_ASAP7_75t_SL g16848 ( 
.A(n_16374),
.Y(n_16848)
);

AND2x2_ASAP7_75t_L g16849 ( 
.A(n_16082),
.B(n_11431),
.Y(n_16849)
);

INVx1_ASAP7_75t_L g16850 ( 
.A(n_16198),
.Y(n_16850)
);

OR2x2_ASAP7_75t_L g16851 ( 
.A(n_15873),
.B(n_11431),
.Y(n_16851)
);

INVx1_ASAP7_75t_L g16852 ( 
.A(n_15992),
.Y(n_16852)
);

HB1xp67_ASAP7_75t_L g16853 ( 
.A(n_16270),
.Y(n_16853)
);

HB1xp67_ASAP7_75t_L g16854 ( 
.A(n_15993),
.Y(n_16854)
);

AND2x2_ASAP7_75t_SL g16855 ( 
.A(n_15911),
.B(n_10539),
.Y(n_16855)
);

NAND2xp5_ASAP7_75t_L g16856 ( 
.A(n_16506),
.B(n_11432),
.Y(n_16856)
);

AND2x2_ASAP7_75t_L g16857 ( 
.A(n_16192),
.B(n_11432),
.Y(n_16857)
);

INVx2_ASAP7_75t_L g16858 ( 
.A(n_16147),
.Y(n_16858)
);

INVx2_ASAP7_75t_L g16859 ( 
.A(n_16145),
.Y(n_16859)
);

NAND2x1p5_ASAP7_75t_L g16860 ( 
.A(n_16027),
.B(n_8232),
.Y(n_16860)
);

INVx1_ASAP7_75t_L g16861 ( 
.A(n_16251),
.Y(n_16861)
);

AND2x2_ASAP7_75t_L g16862 ( 
.A(n_16133),
.B(n_11434),
.Y(n_16862)
);

NOR2x1p5_ASAP7_75t_L g16863 ( 
.A(n_16257),
.B(n_11434),
.Y(n_16863)
);

NAND2xp5_ASAP7_75t_L g16864 ( 
.A(n_16290),
.B(n_11444),
.Y(n_16864)
);

AND2x2_ASAP7_75t_L g16865 ( 
.A(n_16340),
.B(n_11444),
.Y(n_16865)
);

INVx1_ASAP7_75t_L g16866 ( 
.A(n_16483),
.Y(n_16866)
);

NAND2xp5_ASAP7_75t_L g16867 ( 
.A(n_16309),
.B(n_9228),
.Y(n_16867)
);

INVx2_ASAP7_75t_L g16868 ( 
.A(n_16137),
.Y(n_16868)
);

AND2x2_ASAP7_75t_SL g16869 ( 
.A(n_16041),
.B(n_10539),
.Y(n_16869)
);

AND2x2_ASAP7_75t_L g16870 ( 
.A(n_16195),
.B(n_8805),
.Y(n_16870)
);

INVx2_ASAP7_75t_L g16871 ( 
.A(n_16488),
.Y(n_16871)
);

NAND2xp5_ASAP7_75t_L g16872 ( 
.A(n_16197),
.B(n_16204),
.Y(n_16872)
);

NOR2xp67_ASAP7_75t_L g16873 ( 
.A(n_16200),
.B(n_11534),
.Y(n_16873)
);

INVx2_ASAP7_75t_SL g16874 ( 
.A(n_16144),
.Y(n_16874)
);

AOI22xp33_ASAP7_75t_SL g16875 ( 
.A1(n_16370),
.A2(n_11544),
.B1(n_11545),
.B2(n_11543),
.Y(n_16875)
);

AND2x2_ASAP7_75t_L g16876 ( 
.A(n_16044),
.B(n_8805),
.Y(n_16876)
);

AND2x2_ASAP7_75t_L g16877 ( 
.A(n_16071),
.B(n_8805),
.Y(n_16877)
);

INVx3_ASAP7_75t_L g16878 ( 
.A(n_16099),
.Y(n_16878)
);

AND2x2_ASAP7_75t_L g16879 ( 
.A(n_16117),
.B(n_8877),
.Y(n_16879)
);

INVx1_ASAP7_75t_L g16880 ( 
.A(n_16034),
.Y(n_16880)
);

INVx2_ASAP7_75t_L g16881 ( 
.A(n_16312),
.Y(n_16881)
);

NAND2xp5_ASAP7_75t_L g16882 ( 
.A(n_16209),
.B(n_9228),
.Y(n_16882)
);

AND2x2_ASAP7_75t_L g16883 ( 
.A(n_16120),
.B(n_8877),
.Y(n_16883)
);

INVx1_ASAP7_75t_L g16884 ( 
.A(n_15920),
.Y(n_16884)
);

AND2x2_ASAP7_75t_L g16885 ( 
.A(n_16127),
.B(n_16051),
.Y(n_16885)
);

HB1xp67_ASAP7_75t_L g16886 ( 
.A(n_15981),
.Y(n_16886)
);

NAND2xp5_ASAP7_75t_L g16887 ( 
.A(n_16019),
.B(n_9228),
.Y(n_16887)
);

NAND2xp5_ASAP7_75t_L g16888 ( 
.A(n_16375),
.B(n_9228),
.Y(n_16888)
);

INVx2_ASAP7_75t_L g16889 ( 
.A(n_16465),
.Y(n_16889)
);

AOI21xp5_ASAP7_75t_L g16890 ( 
.A1(n_16006),
.A2(n_11544),
.B(n_11543),
.Y(n_16890)
);

INVx2_ASAP7_75t_L g16891 ( 
.A(n_16446),
.Y(n_16891)
);

NAND2xp5_ASAP7_75t_L g16892 ( 
.A(n_16378),
.B(n_9228),
.Y(n_16892)
);

NAND2xp5_ASAP7_75t_L g16893 ( 
.A(n_16253),
.B(n_9228),
.Y(n_16893)
);

AND2x2_ASAP7_75t_L g16894 ( 
.A(n_15994),
.B(n_8877),
.Y(n_16894)
);

NAND2xp5_ASAP7_75t_L g16895 ( 
.A(n_16222),
.B(n_16248),
.Y(n_16895)
);

INVxp67_ASAP7_75t_L g16896 ( 
.A(n_16245),
.Y(n_16896)
);

INVx1_ASAP7_75t_L g16897 ( 
.A(n_15871),
.Y(n_16897)
);

INVx2_ASAP7_75t_L g16898 ( 
.A(n_16455),
.Y(n_16898)
);

AND2x2_ASAP7_75t_L g16899 ( 
.A(n_16001),
.B(n_8895),
.Y(n_16899)
);

AND2x2_ASAP7_75t_L g16900 ( 
.A(n_16190),
.B(n_8895),
.Y(n_16900)
);

OR2x2_ASAP7_75t_L g16901 ( 
.A(n_16238),
.B(n_9091),
.Y(n_16901)
);

AND2x2_ASAP7_75t_L g16902 ( 
.A(n_16324),
.B(n_8895),
.Y(n_16902)
);

NAND2xp5_ASAP7_75t_L g16903 ( 
.A(n_16509),
.B(n_9228),
.Y(n_16903)
);

AND2x2_ASAP7_75t_L g16904 ( 
.A(n_16349),
.B(n_8910),
.Y(n_16904)
);

AND2x2_ASAP7_75t_L g16905 ( 
.A(n_16239),
.B(n_8910),
.Y(n_16905)
);

NAND2xp5_ASAP7_75t_L g16906 ( 
.A(n_16413),
.B(n_9228),
.Y(n_16906)
);

INVx1_ASAP7_75t_L g16907 ( 
.A(n_15892),
.Y(n_16907)
);

BUFx2_ASAP7_75t_SL g16908 ( 
.A(n_15898),
.Y(n_16908)
);

BUFx2_ASAP7_75t_L g16909 ( 
.A(n_16081),
.Y(n_16909)
);

INVx1_ASAP7_75t_L g16910 ( 
.A(n_15919),
.Y(n_16910)
);

INVx1_ASAP7_75t_L g16911 ( 
.A(n_15921),
.Y(n_16911)
);

AND2x2_ASAP7_75t_L g16912 ( 
.A(n_16360),
.B(n_8910),
.Y(n_16912)
);

HB1xp67_ASAP7_75t_L g16913 ( 
.A(n_16391),
.Y(n_16913)
);

AND2x2_ASAP7_75t_L g16914 ( 
.A(n_16414),
.B(n_8949),
.Y(n_16914)
);

AND2x2_ASAP7_75t_L g16915 ( 
.A(n_16417),
.B(n_8949),
.Y(n_16915)
);

INVx1_ASAP7_75t_L g16916 ( 
.A(n_15923),
.Y(n_16916)
);

INVx1_ASAP7_75t_L g16917 ( 
.A(n_15925),
.Y(n_16917)
);

INVx6_ASAP7_75t_L g16918 ( 
.A(n_15913),
.Y(n_16918)
);

NAND2xp5_ASAP7_75t_L g16919 ( 
.A(n_16418),
.B(n_9400),
.Y(n_16919)
);

AND2x2_ASAP7_75t_L g16920 ( 
.A(n_16074),
.B(n_8949),
.Y(n_16920)
);

OR2x2_ASAP7_75t_L g16921 ( 
.A(n_16291),
.B(n_9140),
.Y(n_16921)
);

AND2x2_ASAP7_75t_L g16922 ( 
.A(n_16372),
.B(n_9020),
.Y(n_16922)
);

INVx1_ASAP7_75t_L g16923 ( 
.A(n_16485),
.Y(n_16923)
);

INVx2_ASAP7_75t_L g16924 ( 
.A(n_16450),
.Y(n_16924)
);

OR2x2_ASAP7_75t_L g16925 ( 
.A(n_15902),
.B(n_9140),
.Y(n_16925)
);

AND2x2_ASAP7_75t_L g16926 ( 
.A(n_16327),
.B(n_9020),
.Y(n_16926)
);

INVx1_ASAP7_75t_L g16927 ( 
.A(n_15878),
.Y(n_16927)
);

INVx1_ASAP7_75t_L g16928 ( 
.A(n_16259),
.Y(n_16928)
);

INVx2_ASAP7_75t_L g16929 ( 
.A(n_16469),
.Y(n_16929)
);

AND2x2_ASAP7_75t_L g16930 ( 
.A(n_16293),
.B(n_9020),
.Y(n_16930)
);

INVx1_ASAP7_75t_L g16931 ( 
.A(n_15961),
.Y(n_16931)
);

OR2x2_ASAP7_75t_L g16932 ( 
.A(n_15996),
.B(n_9104),
.Y(n_16932)
);

AND2x4_ASAP7_75t_L g16933 ( 
.A(n_16255),
.B(n_9085),
.Y(n_16933)
);

BUFx2_ASAP7_75t_L g16934 ( 
.A(n_16467),
.Y(n_16934)
);

NAND2xp5_ASAP7_75t_L g16935 ( 
.A(n_16263),
.B(n_16314),
.Y(n_16935)
);

INVx3_ASAP7_75t_L g16936 ( 
.A(n_16085),
.Y(n_16936)
);

BUFx3_ASAP7_75t_L g16937 ( 
.A(n_16262),
.Y(n_16937)
);

INVx1_ASAP7_75t_L g16938 ( 
.A(n_15966),
.Y(n_16938)
);

INVx1_ASAP7_75t_L g16939 ( 
.A(n_15970),
.Y(n_16939)
);

AND2x2_ASAP7_75t_L g16940 ( 
.A(n_16306),
.B(n_9085),
.Y(n_16940)
);

OR2x2_ASAP7_75t_L g16941 ( 
.A(n_15876),
.B(n_9104),
.Y(n_16941)
);

AND2x2_ASAP7_75t_L g16942 ( 
.A(n_16059),
.B(n_9085),
.Y(n_16942)
);

AND2x2_ASAP7_75t_L g16943 ( 
.A(n_16060),
.B(n_16299),
.Y(n_16943)
);

NAND2xp5_ASAP7_75t_L g16944 ( 
.A(n_16346),
.B(n_9428),
.Y(n_16944)
);

AND2x2_ASAP7_75t_L g16945 ( 
.A(n_16319),
.B(n_9137),
.Y(n_16945)
);

INVxp67_ASAP7_75t_L g16946 ( 
.A(n_16033),
.Y(n_16946)
);

INVx1_ASAP7_75t_L g16947 ( 
.A(n_16017),
.Y(n_16947)
);

OR2x2_ASAP7_75t_L g16948 ( 
.A(n_16472),
.B(n_16475),
.Y(n_16948)
);

INVx1_ASAP7_75t_L g16949 ( 
.A(n_16240),
.Y(n_16949)
);

INVx1_ASAP7_75t_L g16950 ( 
.A(n_16298),
.Y(n_16950)
);

INVxp67_ASAP7_75t_L g16951 ( 
.A(n_16126),
.Y(n_16951)
);

INVx1_ASAP7_75t_L g16952 ( 
.A(n_16213),
.Y(n_16952)
);

AND2x2_ASAP7_75t_L g16953 ( 
.A(n_16423),
.B(n_9137),
.Y(n_16953)
);

INVx1_ASAP7_75t_L g16954 ( 
.A(n_16213),
.Y(n_16954)
);

NAND2xp5_ASAP7_75t_L g16955 ( 
.A(n_16356),
.B(n_9449),
.Y(n_16955)
);

OR2x2_ASAP7_75t_L g16956 ( 
.A(n_16478),
.B(n_9104),
.Y(n_16956)
);

NAND2x1p5_ASAP7_75t_L g16957 ( 
.A(n_16479),
.B(n_16481),
.Y(n_16957)
);

AND2x2_ASAP7_75t_L g16958 ( 
.A(n_16426),
.B(n_9137),
.Y(n_16958)
);

AND2x2_ASAP7_75t_L g16959 ( 
.A(n_16433),
.B(n_16436),
.Y(n_16959)
);

INVx1_ASAP7_75t_L g16960 ( 
.A(n_16300),
.Y(n_16960)
);

AND2x2_ASAP7_75t_L g16961 ( 
.A(n_16441),
.B(n_9169),
.Y(n_16961)
);

OR2x2_ASAP7_75t_L g16962 ( 
.A(n_16020),
.B(n_9424),
.Y(n_16962)
);

AND2x2_ASAP7_75t_L g16963 ( 
.A(n_16421),
.B(n_16395),
.Y(n_16963)
);

AND2x2_ASAP7_75t_L g16964 ( 
.A(n_16322),
.B(n_9169),
.Y(n_16964)
);

AND2x2_ASAP7_75t_L g16965 ( 
.A(n_16325),
.B(n_9169),
.Y(n_16965)
);

NAND2xp5_ASAP7_75t_L g16966 ( 
.A(n_16345),
.B(n_9449),
.Y(n_16966)
);

HB1xp67_ASAP7_75t_L g16967 ( 
.A(n_16012),
.Y(n_16967)
);

NAND3xp33_ASAP7_75t_L g16968 ( 
.A(n_16078),
.B(n_11551),
.C(n_11545),
.Y(n_16968)
);

AND2x2_ASAP7_75t_L g16969 ( 
.A(n_16328),
.B(n_9251),
.Y(n_16969)
);

AND2x2_ASAP7_75t_L g16970 ( 
.A(n_16329),
.B(n_9251),
.Y(n_16970)
);

INVx2_ASAP7_75t_L g16971 ( 
.A(n_16471),
.Y(n_16971)
);

INVx1_ASAP7_75t_L g16972 ( 
.A(n_16308),
.Y(n_16972)
);

BUFx2_ASAP7_75t_L g16973 ( 
.A(n_16305),
.Y(n_16973)
);

BUFx3_ASAP7_75t_L g16974 ( 
.A(n_16377),
.Y(n_16974)
);

INVx1_ASAP7_75t_L g16975 ( 
.A(n_16366),
.Y(n_16975)
);

HB1xp67_ASAP7_75t_L g16976 ( 
.A(n_16168),
.Y(n_16976)
);

INVx1_ASAP7_75t_SL g16977 ( 
.A(n_16142),
.Y(n_16977)
);

AND2x2_ASAP7_75t_L g16978 ( 
.A(n_16330),
.B(n_9251),
.Y(n_16978)
);

HB1xp67_ASAP7_75t_L g16979 ( 
.A(n_16362),
.Y(n_16979)
);

OR2x2_ASAP7_75t_L g16980 ( 
.A(n_16223),
.B(n_9424),
.Y(n_16980)
);

AND2x2_ASAP7_75t_L g16981 ( 
.A(n_16317),
.B(n_9313),
.Y(n_16981)
);

INVx2_ASAP7_75t_L g16982 ( 
.A(n_16498),
.Y(n_16982)
);

AND2x2_ASAP7_75t_L g16983 ( 
.A(n_16350),
.B(n_9313),
.Y(n_16983)
);

AND2x2_ASAP7_75t_L g16984 ( 
.A(n_16380),
.B(n_9313),
.Y(n_16984)
);

INVx1_ASAP7_75t_L g16985 ( 
.A(n_16143),
.Y(n_16985)
);

AND2x2_ASAP7_75t_L g16986 ( 
.A(n_16408),
.B(n_9350),
.Y(n_16986)
);

AND2x2_ASAP7_75t_L g16987 ( 
.A(n_16424),
.B(n_9350),
.Y(n_16987)
);

AND2x2_ASAP7_75t_L g16988 ( 
.A(n_16171),
.B(n_9350),
.Y(n_16988)
);

HB1xp67_ASAP7_75t_L g16989 ( 
.A(n_16365),
.Y(n_16989)
);

BUFx3_ASAP7_75t_L g16990 ( 
.A(n_16342),
.Y(n_16990)
);

OR2x2_ASAP7_75t_L g16991 ( 
.A(n_16422),
.B(n_9451),
.Y(n_16991)
);

INVx2_ASAP7_75t_L g16992 ( 
.A(n_16458),
.Y(n_16992)
);

NAND2xp5_ASAP7_75t_L g16993 ( 
.A(n_16264),
.B(n_9451),
.Y(n_16993)
);

NAND2xp5_ASAP7_75t_L g16994 ( 
.A(n_16276),
.B(n_16283),
.Y(n_16994)
);

AND2x2_ASAP7_75t_L g16995 ( 
.A(n_16486),
.B(n_9476),
.Y(n_16995)
);

AND2x2_ASAP7_75t_L g16996 ( 
.A(n_16353),
.B(n_9476),
.Y(n_16996)
);

AND2x2_ASAP7_75t_L g16997 ( 
.A(n_16384),
.B(n_9476),
.Y(n_16997)
);

AND2x2_ASAP7_75t_L g16998 ( 
.A(n_16394),
.B(n_9484),
.Y(n_16998)
);

OR2x2_ASAP7_75t_L g16999 ( 
.A(n_16091),
.B(n_9347),
.Y(n_16999)
);

INVx1_ASAP7_75t_L g17000 ( 
.A(n_16154),
.Y(n_17000)
);

HB1xp67_ASAP7_75t_L g17001 ( 
.A(n_16115),
.Y(n_17001)
);

INVx2_ASAP7_75t_L g17002 ( 
.A(n_16460),
.Y(n_17002)
);

NOR2x1_ASAP7_75t_L g17003 ( 
.A(n_16305),
.B(n_11551),
.Y(n_17003)
);

NAND2xp5_ASAP7_75t_L g17004 ( 
.A(n_16295),
.B(n_11554),
.Y(n_17004)
);

AND2x4_ASAP7_75t_L g17005 ( 
.A(n_16348),
.B(n_9484),
.Y(n_17005)
);

HB1xp67_ASAP7_75t_L g17006 ( 
.A(n_16116),
.Y(n_17006)
);

INVx1_ASAP7_75t_L g17007 ( 
.A(n_16169),
.Y(n_17007)
);

INVx2_ASAP7_75t_L g17008 ( 
.A(n_16473),
.Y(n_17008)
);

NAND2xp5_ASAP7_75t_L g17009 ( 
.A(n_16504),
.B(n_11554),
.Y(n_17009)
);

HB1xp67_ASAP7_75t_L g17010 ( 
.A(n_16047),
.Y(n_17010)
);

OR2x2_ASAP7_75t_L g17011 ( 
.A(n_16438),
.B(n_9347),
.Y(n_17011)
);

NAND2xp5_ASAP7_75t_L g17012 ( 
.A(n_16407),
.B(n_11555),
.Y(n_17012)
);

OR2x2_ASAP7_75t_L g17013 ( 
.A(n_16220),
.B(n_9347),
.Y(n_17013)
);

INVx1_ASAP7_75t_L g17014 ( 
.A(n_16386),
.Y(n_17014)
);

INVx1_ASAP7_75t_L g17015 ( 
.A(n_16493),
.Y(n_17015)
);

INVx1_ASAP7_75t_L g17016 ( 
.A(n_16495),
.Y(n_17016)
);

OAI211xp5_ASAP7_75t_L g17017 ( 
.A1(n_16162),
.A2(n_11555),
.B(n_11559),
.C(n_11558),
.Y(n_17017)
);

OR2x2_ASAP7_75t_L g17018 ( 
.A(n_16484),
.B(n_16079),
.Y(n_17018)
);

NOR2xp33_ASAP7_75t_R g17019 ( 
.A(n_16230),
.B(n_7076),
.Y(n_17019)
);

AND2x4_ASAP7_75t_L g17020 ( 
.A(n_16351),
.B(n_9484),
.Y(n_17020)
);

INVxp67_ASAP7_75t_SL g17021 ( 
.A(n_16045),
.Y(n_17021)
);

AOI22xp33_ASAP7_75t_L g17022 ( 
.A1(n_16094),
.A2(n_11565),
.B1(n_11566),
.B2(n_11563),
.Y(n_17022)
);

AND2x2_ASAP7_75t_L g17023 ( 
.A(n_16205),
.B(n_9519),
.Y(n_17023)
);

AND2x2_ASAP7_75t_L g17024 ( 
.A(n_16237),
.B(n_16061),
.Y(n_17024)
);

NAND2xp5_ASAP7_75t_L g17025 ( 
.A(n_16507),
.B(n_11571),
.Y(n_17025)
);

INVx4_ASAP7_75t_L g17026 ( 
.A(n_16520),
.Y(n_17026)
);

INVx1_ASAP7_75t_L g17027 ( 
.A(n_16320),
.Y(n_17027)
);

NAND2xp5_ASAP7_75t_L g17028 ( 
.A(n_16321),
.B(n_11571),
.Y(n_17028)
);

AND2x4_ASAP7_75t_L g17029 ( 
.A(n_16247),
.B(n_9519),
.Y(n_17029)
);

AND2x2_ASAP7_75t_L g17030 ( 
.A(n_16258),
.B(n_9519),
.Y(n_17030)
);

AND2x2_ASAP7_75t_L g17031 ( 
.A(n_16515),
.B(n_11574),
.Y(n_17031)
);

INVx1_ASAP7_75t_L g17032 ( 
.A(n_16289),
.Y(n_17032)
);

AND2x2_ASAP7_75t_L g17033 ( 
.A(n_16215),
.B(n_11574),
.Y(n_17033)
);

AND2x2_ASAP7_75t_L g17034 ( 
.A(n_16217),
.B(n_11575),
.Y(n_17034)
);

INVxp67_ASAP7_75t_L g17035 ( 
.A(n_16070),
.Y(n_17035)
);

INVx4_ASAP7_75t_L g17036 ( 
.A(n_16175),
.Y(n_17036)
);

AND2x2_ASAP7_75t_L g17037 ( 
.A(n_16361),
.B(n_11575),
.Y(n_17037)
);

INVx2_ASAP7_75t_L g17038 ( 
.A(n_16463),
.Y(n_17038)
);

INVx2_ASAP7_75t_L g17039 ( 
.A(n_16496),
.Y(n_17039)
);

INVx1_ASAP7_75t_L g17040 ( 
.A(n_16359),
.Y(n_17040)
);

AND2x4_ASAP7_75t_L g17041 ( 
.A(n_16177),
.B(n_10591),
.Y(n_17041)
);

INVx1_ASAP7_75t_SL g17042 ( 
.A(n_16055),
.Y(n_17042)
);

INVxp67_ASAP7_75t_L g17043 ( 
.A(n_16339),
.Y(n_17043)
);

INVx1_ASAP7_75t_SL g17044 ( 
.A(n_16182),
.Y(n_17044)
);

NAND2xp5_ASAP7_75t_L g17045 ( 
.A(n_16453),
.B(n_11583),
.Y(n_17045)
);

AND2x2_ASAP7_75t_L g17046 ( 
.A(n_16464),
.B(n_11583),
.Y(n_17046)
);

AND2x2_ASAP7_75t_L g17047 ( 
.A(n_16093),
.B(n_11594),
.Y(n_17047)
);

NAND2xp5_ASAP7_75t_L g17048 ( 
.A(n_16454),
.B(n_16457),
.Y(n_17048)
);

INVx1_ASAP7_75t_L g17049 ( 
.A(n_16400),
.Y(n_17049)
);

AND2x2_ASAP7_75t_L g17050 ( 
.A(n_16416),
.B(n_11594),
.Y(n_17050)
);

INVx1_ASAP7_75t_L g17051 ( 
.A(n_16503),
.Y(n_17051)
);

NAND2xp5_ASAP7_75t_L g17052 ( 
.A(n_16461),
.B(n_11610),
.Y(n_17052)
);

INVx1_ASAP7_75t_L g17053 ( 
.A(n_16383),
.Y(n_17053)
);

AND2x2_ASAP7_75t_L g17054 ( 
.A(n_16482),
.B(n_11610),
.Y(n_17054)
);

INVx1_ASAP7_75t_L g17055 ( 
.A(n_16206),
.Y(n_17055)
);

INVx1_ASAP7_75t_L g17056 ( 
.A(n_16203),
.Y(n_17056)
);

INVx2_ASAP7_75t_L g17057 ( 
.A(n_16492),
.Y(n_17057)
);

INVx2_ASAP7_75t_L g17058 ( 
.A(n_16252),
.Y(n_17058)
);

INVx1_ASAP7_75t_L g17059 ( 
.A(n_16302),
.Y(n_17059)
);

AND2x2_ASAP7_75t_L g17060 ( 
.A(n_16508),
.B(n_11616),
.Y(n_17060)
);

OR2x2_ASAP7_75t_L g17061 ( 
.A(n_16428),
.B(n_9367),
.Y(n_17061)
);

INVx1_ASAP7_75t_L g17062 ( 
.A(n_16313),
.Y(n_17062)
);

INVx1_ASAP7_75t_L g17063 ( 
.A(n_16318),
.Y(n_17063)
);

INVx2_ASAP7_75t_L g17064 ( 
.A(n_16279),
.Y(n_17064)
);

HB1xp67_ASAP7_75t_L g17065 ( 
.A(n_16181),
.Y(n_17065)
);

AND2x2_ASAP7_75t_L g17066 ( 
.A(n_16513),
.B(n_11616),
.Y(n_17066)
);

AND2x2_ASAP7_75t_L g17067 ( 
.A(n_16519),
.B(n_11634),
.Y(n_17067)
);

INVx1_ASAP7_75t_L g17068 ( 
.A(n_16331),
.Y(n_17068)
);

INVx2_ASAP7_75t_L g17069 ( 
.A(n_16284),
.Y(n_17069)
);

OR2x2_ASAP7_75t_L g17070 ( 
.A(n_16430),
.B(n_9367),
.Y(n_17070)
);

HB1xp67_ASAP7_75t_L g17071 ( 
.A(n_16194),
.Y(n_17071)
);

OR2x2_ASAP7_75t_L g17072 ( 
.A(n_16432),
.B(n_9367),
.Y(n_17072)
);

HB1xp67_ASAP7_75t_L g17073 ( 
.A(n_16201),
.Y(n_17073)
);

INVx1_ASAP7_75t_L g17074 ( 
.A(n_16344),
.Y(n_17074)
);

NAND2xp5_ASAP7_75t_L g17075 ( 
.A(n_16427),
.B(n_11634),
.Y(n_17075)
);

AND2x2_ASAP7_75t_L g17076 ( 
.A(n_16355),
.B(n_11645),
.Y(n_17076)
);

INVx1_ASAP7_75t_L g17077 ( 
.A(n_16357),
.Y(n_17077)
);

OR2x2_ASAP7_75t_L g17078 ( 
.A(n_16207),
.B(n_16216),
.Y(n_17078)
);

INVx1_ASAP7_75t_L g17079 ( 
.A(n_16323),
.Y(n_17079)
);

AOI22xp33_ASAP7_75t_L g17080 ( 
.A1(n_16500),
.A2(n_11648),
.B1(n_11649),
.B2(n_11645),
.Y(n_17080)
);

INVx1_ASAP7_75t_L g17081 ( 
.A(n_15916),
.Y(n_17081)
);

INVx1_ASAP7_75t_SL g17082 ( 
.A(n_16063),
.Y(n_17082)
);

OR2x6_ASAP7_75t_L g17083 ( 
.A(n_16219),
.B(n_10424),
.Y(n_17083)
);

NAND2x1p5_ASAP7_75t_L g17084 ( 
.A(n_16420),
.B(n_8232),
.Y(n_17084)
);

AND2x2_ASAP7_75t_L g17085 ( 
.A(n_16397),
.B(n_11648),
.Y(n_17085)
);

OR2x6_ASAP7_75t_L g17086 ( 
.A(n_16516),
.B(n_10424),
.Y(n_17086)
);

AND2x2_ASAP7_75t_L g17087 ( 
.A(n_16310),
.B(n_11649),
.Y(n_17087)
);

INVx2_ASAP7_75t_SL g17088 ( 
.A(n_16106),
.Y(n_17088)
);

INVx2_ASAP7_75t_L g17089 ( 
.A(n_16412),
.Y(n_17089)
);

INVx1_ASAP7_75t_L g17090 ( 
.A(n_16297),
.Y(n_17090)
);

INVx2_ASAP7_75t_L g17091 ( 
.A(n_16466),
.Y(n_17091)
);

NOR2x1_ASAP7_75t_L g17092 ( 
.A(n_16447),
.B(n_11650),
.Y(n_17092)
);

OR2x2_ASAP7_75t_L g17093 ( 
.A(n_16411),
.B(n_9369),
.Y(n_17093)
);

HB1xp67_ASAP7_75t_L g17094 ( 
.A(n_16053),
.Y(n_17094)
);

AND2x2_ASAP7_75t_L g17095 ( 
.A(n_16451),
.B(n_11650),
.Y(n_17095)
);

AND2x2_ASAP7_75t_L g17096 ( 
.A(n_16489),
.B(n_11660),
.Y(n_17096)
);

INVx2_ASAP7_75t_L g17097 ( 
.A(n_16466),
.Y(n_17097)
);

INVx2_ASAP7_75t_SL g17098 ( 
.A(n_16231),
.Y(n_17098)
);

AND2x2_ASAP7_75t_L g17099 ( 
.A(n_16499),
.B(n_11660),
.Y(n_17099)
);

OR2x2_ASAP7_75t_L g17100 ( 
.A(n_16232),
.B(n_9369),
.Y(n_17100)
);

INVx2_ASAP7_75t_L g17101 ( 
.A(n_16585),
.Y(n_17101)
);

INVx1_ASAP7_75t_L g17102 ( 
.A(n_16973),
.Y(n_17102)
);

NOR2xp33_ASAP7_75t_L g17103 ( 
.A(n_16723),
.B(n_16437),
.Y(n_17103)
);

NOR3xp33_ASAP7_75t_L g17104 ( 
.A(n_16724),
.B(n_16072),
.C(n_16058),
.Y(n_17104)
);

AND2x2_ASAP7_75t_L g17105 ( 
.A(n_16629),
.B(n_16501),
.Y(n_17105)
);

INVx1_ASAP7_75t_SL g17106 ( 
.A(n_16885),
.Y(n_17106)
);

HB1xp67_ASAP7_75t_L g17107 ( 
.A(n_16973),
.Y(n_17107)
);

NAND2x1p5_ASAP7_75t_L g17108 ( 
.A(n_16673),
.B(n_16440),
.Y(n_17108)
);

OR2x2_ASAP7_75t_L g17109 ( 
.A(n_16575),
.B(n_16135),
.Y(n_17109)
);

NAND2xp5_ASAP7_75t_L g17110 ( 
.A(n_16639),
.B(n_16443),
.Y(n_17110)
);

INVx2_ASAP7_75t_L g17111 ( 
.A(n_16770),
.Y(n_17111)
);

INVx1_ASAP7_75t_L g17112 ( 
.A(n_16853),
.Y(n_17112)
);

INVx1_ASAP7_75t_L g17113 ( 
.A(n_16918),
.Y(n_17113)
);

AND2x2_ASAP7_75t_L g17114 ( 
.A(n_16676),
.B(n_16698),
.Y(n_17114)
);

INVx1_ASAP7_75t_L g17115 ( 
.A(n_16918),
.Y(n_17115)
);

OR2x2_ASAP7_75t_L g17116 ( 
.A(n_16531),
.B(n_16235),
.Y(n_17116)
);

INVx1_ASAP7_75t_L g17117 ( 
.A(n_16810),
.Y(n_17117)
);

INVx1_ASAP7_75t_L g17118 ( 
.A(n_16913),
.Y(n_17118)
);

AOI21xp5_ASAP7_75t_L g17119 ( 
.A1(n_16551),
.A2(n_16193),
.B(n_16510),
.Y(n_17119)
);

NAND2xp5_ASAP7_75t_L g17120 ( 
.A(n_16527),
.B(n_16445),
.Y(n_17120)
);

AND2x4_ASAP7_75t_L g17121 ( 
.A(n_16594),
.B(n_16511),
.Y(n_17121)
);

AND2x2_ASAP7_75t_L g17122 ( 
.A(n_16641),
.B(n_16512),
.Y(n_17122)
);

NAND2x1p5_ASAP7_75t_L g17123 ( 
.A(n_16717),
.B(n_16514),
.Y(n_17123)
);

INVx1_ASAP7_75t_L g17124 ( 
.A(n_16526),
.Y(n_17124)
);

NOR2xp67_ASAP7_75t_L g17125 ( 
.A(n_16544),
.B(n_16112),
.Y(n_17125)
);

AND2x2_ASAP7_75t_L g17126 ( 
.A(n_16701),
.B(n_16517),
.Y(n_17126)
);

AND2x2_ASAP7_75t_L g17127 ( 
.A(n_16943),
.B(n_16521),
.Y(n_17127)
);

NAND2x2_ASAP7_75t_L g17128 ( 
.A(n_16990),
.B(n_16104),
.Y(n_17128)
);

HB1xp67_ASAP7_75t_L g17129 ( 
.A(n_16636),
.Y(n_17129)
);

AND2x4_ASAP7_75t_L g17130 ( 
.A(n_16600),
.B(n_16720),
.Y(n_17130)
);

NAND2xp5_ASAP7_75t_L g17131 ( 
.A(n_16560),
.B(n_16522),
.Y(n_17131)
);

AND2x2_ASAP7_75t_L g17132 ( 
.A(n_16539),
.B(n_16523),
.Y(n_17132)
);

INVx1_ASAP7_75t_SL g17133 ( 
.A(n_16789),
.Y(n_17133)
);

AND2x2_ASAP7_75t_L g17134 ( 
.A(n_16534),
.B(n_16387),
.Y(n_17134)
);

NAND2xp33_ASAP7_75t_SL g17135 ( 
.A(n_16533),
.B(n_16287),
.Y(n_17135)
);

AND2x2_ASAP7_75t_L g17136 ( 
.A(n_16553),
.B(n_16388),
.Y(n_17136)
);

AND2x2_ASAP7_75t_L g17137 ( 
.A(n_16836),
.B(n_16536),
.Y(n_17137)
);

INVx1_ASAP7_75t_L g17138 ( 
.A(n_16574),
.Y(n_17138)
);

INVx2_ASAP7_75t_L g17139 ( 
.A(n_17018),
.Y(n_17139)
);

INVx1_ASAP7_75t_L g17140 ( 
.A(n_17001),
.Y(n_17140)
);

INVx2_ASAP7_75t_L g17141 ( 
.A(n_16636),
.Y(n_17141)
);

AND2x2_ASAP7_75t_L g17142 ( 
.A(n_16909),
.B(n_16393),
.Y(n_17142)
);

AOI221x1_ASAP7_75t_L g17143 ( 
.A1(n_16601),
.A2(n_16077),
.B1(n_16076),
.B2(n_16073),
.C(n_16398),
.Y(n_17143)
);

AND2x2_ASAP7_75t_L g17144 ( 
.A(n_16709),
.B(n_16403),
.Y(n_17144)
);

INVx2_ASAP7_75t_L g17145 ( 
.A(n_16599),
.Y(n_17145)
);

NAND2xp5_ASAP7_75t_L g17146 ( 
.A(n_16977),
.B(n_16405),
.Y(n_17146)
);

INVx4_ASAP7_75t_L g17147 ( 
.A(n_16712),
.Y(n_17147)
);

HB1xp67_ASAP7_75t_L g17148 ( 
.A(n_16734),
.Y(n_17148)
);

AND2x4_ASAP7_75t_L g17149 ( 
.A(n_16530),
.B(n_16410),
.Y(n_17149)
);

INVx2_ASAP7_75t_L g17150 ( 
.A(n_16608),
.Y(n_17150)
);

NOR2x1_ASAP7_75t_SL g17151 ( 
.A(n_16654),
.B(n_16419),
.Y(n_17151)
);

INVx1_ASAP7_75t_L g17152 ( 
.A(n_17006),
.Y(n_17152)
);

INVx1_ASAP7_75t_L g17153 ( 
.A(n_16598),
.Y(n_17153)
);

AND2x4_ASAP7_75t_L g17154 ( 
.A(n_16700),
.B(n_16242),
.Y(n_17154)
);

BUFx2_ASAP7_75t_SL g17155 ( 
.A(n_16543),
.Y(n_17155)
);

AND2x2_ASAP7_75t_L g17156 ( 
.A(n_16623),
.B(n_16103),
.Y(n_17156)
);

NAND2xp5_ASAP7_75t_SL g17157 ( 
.A(n_16566),
.B(n_16234),
.Y(n_17157)
);

INVxp33_ASAP7_75t_L g17158 ( 
.A(n_16646),
.Y(n_17158)
);

HB1xp67_ASAP7_75t_L g17159 ( 
.A(n_16537),
.Y(n_17159)
);

OR2x2_ASAP7_75t_L g17160 ( 
.A(n_16593),
.B(n_16246),
.Y(n_17160)
);

AOI21xp5_ASAP7_75t_L g17161 ( 
.A1(n_16559),
.A2(n_16497),
.B(n_16476),
.Y(n_17161)
);

INVx2_ASAP7_75t_L g17162 ( 
.A(n_16576),
.Y(n_17162)
);

INVx1_ASAP7_75t_L g17163 ( 
.A(n_16682),
.Y(n_17163)
);

AND2x2_ASAP7_75t_L g17164 ( 
.A(n_16622),
.B(n_16266),
.Y(n_17164)
);

INVx3_ASAP7_75t_L g17165 ( 
.A(n_17026),
.Y(n_17165)
);

AND2x2_ASAP7_75t_L g17166 ( 
.A(n_16563),
.B(n_16268),
.Y(n_17166)
);

NOR2x1_ASAP7_75t_L g17167 ( 
.A(n_16525),
.B(n_16110),
.Y(n_17167)
);

AND2x2_ASAP7_75t_L g17168 ( 
.A(n_16768),
.B(n_16277),
.Y(n_17168)
);

INVx1_ASAP7_75t_L g17169 ( 
.A(n_16573),
.Y(n_17169)
);

INVx2_ASAP7_75t_L g17170 ( 
.A(n_16957),
.Y(n_17170)
);

NAND2xp5_ASAP7_75t_L g17171 ( 
.A(n_16569),
.B(n_16583),
.Y(n_17171)
);

AND2x2_ASAP7_75t_L g17172 ( 
.A(n_16572),
.B(n_16286),
.Y(n_17172)
);

INVx1_ASAP7_75t_L g17173 ( 
.A(n_16603),
.Y(n_17173)
);

INVx2_ASAP7_75t_L g17174 ( 
.A(n_16627),
.Y(n_17174)
);

AND2x2_ASAP7_75t_L g17175 ( 
.A(n_16565),
.B(n_16294),
.Y(n_17175)
);

HB1xp67_ASAP7_75t_L g17176 ( 
.A(n_16704),
.Y(n_17176)
);

NAND2xp5_ASAP7_75t_L g17177 ( 
.A(n_16604),
.B(n_16211),
.Y(n_17177)
);

OAI31xp33_ASAP7_75t_SL g17178 ( 
.A1(n_16638),
.A2(n_16138),
.A3(n_16281),
.B(n_11916),
.Y(n_17178)
);

AND2x2_ASAP7_75t_L g17179 ( 
.A(n_16626),
.B(n_16311),
.Y(n_17179)
);

INVx1_ASAP7_75t_L g17180 ( 
.A(n_16678),
.Y(n_17180)
);

AND2x2_ASAP7_75t_L g17181 ( 
.A(n_16835),
.B(n_16354),
.Y(n_17181)
);

HB1xp67_ASAP7_75t_L g17182 ( 
.A(n_16671),
.Y(n_17182)
);

AND2x4_ASAP7_75t_L g17183 ( 
.A(n_16740),
.B(n_16364),
.Y(n_17183)
);

AND2x2_ASAP7_75t_L g17184 ( 
.A(n_16959),
.B(n_16335),
.Y(n_17184)
);

AND2x2_ASAP7_75t_L g17185 ( 
.A(n_16788),
.B(n_16389),
.Y(n_17185)
);

OR2x2_ASAP7_75t_L g17186 ( 
.A(n_16686),
.B(n_16828),
.Y(n_17186)
);

NAND2xp5_ASAP7_75t_L g17187 ( 
.A(n_17021),
.B(n_16449),
.Y(n_17187)
);

NAND2xp5_ASAP7_75t_L g17188 ( 
.A(n_16647),
.B(n_16477),
.Y(n_17188)
);

HB1xp67_ASAP7_75t_L g17189 ( 
.A(n_16689),
.Y(n_17189)
);

NOR3xp33_ASAP7_75t_L g17190 ( 
.A(n_16797),
.B(n_16487),
.C(n_16518),
.Y(n_17190)
);

AND2x2_ASAP7_75t_L g17191 ( 
.A(n_16845),
.B(n_16124),
.Y(n_17191)
);

INVx1_ASAP7_75t_L g17192 ( 
.A(n_16540),
.Y(n_17192)
);

INVx1_ASAP7_75t_L g17193 ( 
.A(n_16542),
.Y(n_17193)
);

AOI22x1_ASAP7_75t_L g17194 ( 
.A1(n_16675),
.A2(n_11824),
.B1(n_11825),
.B2(n_11811),
.Y(n_17194)
);

INVx1_ASAP7_75t_L g17195 ( 
.A(n_16552),
.Y(n_17195)
);

INVx2_ASAP7_75t_L g17196 ( 
.A(n_16591),
.Y(n_17196)
);

NAND2x1_ASAP7_75t_SL g17197 ( 
.A(n_16979),
.B(n_11661),
.Y(n_17197)
);

AND2x2_ASAP7_75t_L g17198 ( 
.A(n_16535),
.B(n_16134),
.Y(n_17198)
);

AND2x2_ASAP7_75t_L g17199 ( 
.A(n_16644),
.B(n_11661),
.Y(n_17199)
);

AND2x4_ASAP7_75t_L g17200 ( 
.A(n_16937),
.B(n_16963),
.Y(n_17200)
);

AND2x2_ASAP7_75t_L g17201 ( 
.A(n_16617),
.B(n_11669),
.Y(n_17201)
);

AND2x4_ASAP7_75t_L g17202 ( 
.A(n_16706),
.B(n_11669),
.Y(n_17202)
);

OR2x2_ASAP7_75t_L g17203 ( 
.A(n_16581),
.B(n_11675),
.Y(n_17203)
);

INVx1_ASAP7_75t_SL g17204 ( 
.A(n_16645),
.Y(n_17204)
);

AND2x2_ASAP7_75t_L g17205 ( 
.A(n_16616),
.B(n_11675),
.Y(n_17205)
);

INVx3_ASAP7_75t_L g17206 ( 
.A(n_16813),
.Y(n_17206)
);

INVx1_ASAP7_75t_L g17207 ( 
.A(n_16783),
.Y(n_17207)
);

INVx2_ASAP7_75t_L g17208 ( 
.A(n_16715),
.Y(n_17208)
);

OR2x2_ASAP7_75t_L g17209 ( 
.A(n_16597),
.B(n_11677),
.Y(n_17209)
);

NAND4xp25_ASAP7_75t_L g17210 ( 
.A(n_16685),
.B(n_11677),
.C(n_11693),
.D(n_11692),
.Y(n_17210)
);

AND2x2_ASAP7_75t_L g17211 ( 
.A(n_16719),
.B(n_11692),
.Y(n_17211)
);

INVx1_ASAP7_75t_SL g17212 ( 
.A(n_17042),
.Y(n_17212)
);

AND2x2_ASAP7_75t_L g17213 ( 
.A(n_16719),
.B(n_11693),
.Y(n_17213)
);

INVx1_ASAP7_75t_L g17214 ( 
.A(n_16783),
.Y(n_17214)
);

INVxp33_ASAP7_75t_L g17215 ( 
.A(n_16596),
.Y(n_17215)
);

INVx1_ASAP7_75t_L g17216 ( 
.A(n_16934),
.Y(n_17216)
);

INVx2_ASAP7_75t_L g17217 ( 
.A(n_16813),
.Y(n_17217)
);

AND2x2_ASAP7_75t_L g17218 ( 
.A(n_16570),
.B(n_11811),
.Y(n_17218)
);

INVx1_ASAP7_75t_L g17219 ( 
.A(n_16735),
.Y(n_17219)
);

NOR2xp33_ASAP7_75t_L g17220 ( 
.A(n_16830),
.B(n_17036),
.Y(n_17220)
);

NOR3xp33_ASAP7_75t_L g17221 ( 
.A(n_16691),
.B(n_11825),
.C(n_11824),
.Y(n_17221)
);

AND2x2_ASAP7_75t_L g17222 ( 
.A(n_16657),
.B(n_16562),
.Y(n_17222)
);

OAI21xp5_ASAP7_75t_L g17223 ( 
.A1(n_16524),
.A2(n_11262),
.B(n_11258),
.Y(n_17223)
);

NAND2xp5_ASAP7_75t_L g17224 ( 
.A(n_16830),
.B(n_11833),
.Y(n_17224)
);

AND2x2_ASAP7_75t_L g17225 ( 
.A(n_16684),
.B(n_11833),
.Y(n_17225)
);

OR2x2_ASAP7_75t_L g17226 ( 
.A(n_16606),
.B(n_11841),
.Y(n_17226)
);

OR2x2_ASAP7_75t_L g17227 ( 
.A(n_16612),
.B(n_11841),
.Y(n_17227)
);

NAND2xp5_ASAP7_75t_L g17228 ( 
.A(n_16830),
.B(n_11846),
.Y(n_17228)
);

OAI21xp33_ASAP7_75t_L g17229 ( 
.A1(n_16642),
.A2(n_11849),
.B(n_11846),
.Y(n_17229)
);

INVx2_ASAP7_75t_L g17230 ( 
.A(n_16869),
.Y(n_17230)
);

OR2x2_ASAP7_75t_L g17231 ( 
.A(n_16726),
.B(n_11849),
.Y(n_17231)
);

AND2x2_ASAP7_75t_L g17232 ( 
.A(n_16613),
.B(n_11851),
.Y(n_17232)
);

INVx1_ASAP7_75t_SL g17233 ( 
.A(n_16628),
.Y(n_17233)
);

INVx1_ASAP7_75t_L g17234 ( 
.A(n_16538),
.Y(n_17234)
);

HB1xp67_ASAP7_75t_L g17235 ( 
.A(n_17003),
.Y(n_17235)
);

INVx1_ASAP7_75t_L g17236 ( 
.A(n_16952),
.Y(n_17236)
);

AND2x2_ASAP7_75t_L g17237 ( 
.A(n_16619),
.B(n_11851),
.Y(n_17237)
);

NAND2xp5_ASAP7_75t_L g17238 ( 
.A(n_17044),
.B(n_11852),
.Y(n_17238)
);

AND2x2_ASAP7_75t_L g17239 ( 
.A(n_16592),
.B(n_11852),
.Y(n_17239)
);

OAI31xp33_ASAP7_75t_L g17240 ( 
.A1(n_17017),
.A2(n_11867),
.A3(n_11871),
.B(n_11854),
.Y(n_17240)
);

AND2x2_ASAP7_75t_L g17241 ( 
.A(n_16660),
.B(n_11854),
.Y(n_17241)
);

HB1xp67_ASAP7_75t_L g17242 ( 
.A(n_16954),
.Y(n_17242)
);

NAND2xp5_ASAP7_75t_L g17243 ( 
.A(n_16656),
.B(n_11867),
.Y(n_17243)
);

AND2x2_ASAP7_75t_L g17244 ( 
.A(n_16743),
.B(n_11871),
.Y(n_17244)
);

INVx1_ASAP7_75t_L g17245 ( 
.A(n_16886),
.Y(n_17245)
);

INVx1_ASAP7_75t_L g17246 ( 
.A(n_16989),
.Y(n_17246)
);

INVx1_ASAP7_75t_L g17247 ( 
.A(n_16854),
.Y(n_17247)
);

AND2x2_ASAP7_75t_L g17248 ( 
.A(n_16936),
.B(n_11874),
.Y(n_17248)
);

AND2x4_ASAP7_75t_L g17249 ( 
.A(n_16974),
.B(n_16567),
.Y(n_17249)
);

INVx1_ASAP7_75t_L g17250 ( 
.A(n_16819),
.Y(n_17250)
);

INVx2_ASAP7_75t_L g17251 ( 
.A(n_17083),
.Y(n_17251)
);

AND2x2_ASAP7_75t_L g17252 ( 
.A(n_16790),
.B(n_11874),
.Y(n_17252)
);

AOI22xp33_ASAP7_75t_L g17253 ( 
.A1(n_16609),
.A2(n_11886),
.B1(n_11909),
.B2(n_11884),
.Y(n_17253)
);

INVx3_ASAP7_75t_L g17254 ( 
.A(n_17083),
.Y(n_17254)
);

INVx1_ASAP7_75t_L g17255 ( 
.A(n_16615),
.Y(n_17255)
);

AND2x2_ASAP7_75t_L g17256 ( 
.A(n_16767),
.B(n_11884),
.Y(n_17256)
);

AND2x2_ASAP7_75t_L g17257 ( 
.A(n_16755),
.B(n_11886),
.Y(n_17257)
);

NAND2x1p5_ASAP7_75t_L g17258 ( 
.A(n_16548),
.B(n_8232),
.Y(n_17258)
);

CKINVDCx6p67_ASAP7_75t_R g17259 ( 
.A(n_16791),
.Y(n_17259)
);

NAND2xp5_ASAP7_75t_L g17260 ( 
.A(n_16651),
.B(n_17089),
.Y(n_17260)
);

OR2x2_ASAP7_75t_L g17261 ( 
.A(n_16632),
.B(n_11909),
.Y(n_17261)
);

INVx1_ASAP7_75t_SL g17262 ( 
.A(n_16554),
.Y(n_17262)
);

AND2x4_ASAP7_75t_L g17263 ( 
.A(n_16874),
.B(n_8494),
.Y(n_17263)
);

AND2x2_ASAP7_75t_L g17264 ( 
.A(n_17041),
.B(n_11920),
.Y(n_17264)
);

OR2x2_ASAP7_75t_L g17265 ( 
.A(n_16633),
.B(n_16637),
.Y(n_17265)
);

NAND2xp5_ASAP7_75t_L g17266 ( 
.A(n_16866),
.B(n_11920),
.Y(n_17266)
);

INVx1_ASAP7_75t_L g17267 ( 
.A(n_16625),
.Y(n_17267)
);

OAI22xp5_ASAP7_75t_L g17268 ( 
.A1(n_16702),
.A2(n_11926),
.B1(n_11936),
.B2(n_11925),
.Y(n_17268)
);

INVx1_ASAP7_75t_L g17269 ( 
.A(n_17065),
.Y(n_17269)
);

INVx1_ASAP7_75t_L g17270 ( 
.A(n_17071),
.Y(n_17270)
);

AND2x2_ASAP7_75t_L g17271 ( 
.A(n_16634),
.B(n_11925),
.Y(n_17271)
);

NOR2xp33_ASAP7_75t_R g17272 ( 
.A(n_16923),
.B(n_7076),
.Y(n_17272)
);

AND2x2_ASAP7_75t_L g17273 ( 
.A(n_16568),
.B(n_16878),
.Y(n_17273)
);

NAND2xp5_ASAP7_75t_L g17274 ( 
.A(n_16661),
.B(n_11926),
.Y(n_17274)
);

AND2x2_ASAP7_75t_L g17275 ( 
.A(n_16669),
.B(n_11936),
.Y(n_17275)
);

AND2x2_ASAP7_75t_L g17276 ( 
.A(n_16561),
.B(n_11937),
.Y(n_17276)
);

AND2x4_ASAP7_75t_L g17277 ( 
.A(n_16580),
.B(n_11937),
.Y(n_17277)
);

NAND2xp5_ASAP7_75t_SL g17278 ( 
.A(n_16586),
.B(n_10539),
.Y(n_17278)
);

OAI21x1_ASAP7_75t_L g17279 ( 
.A1(n_16614),
.A2(n_11952),
.B(n_11939),
.Y(n_17279)
);

INVx1_ASAP7_75t_L g17280 ( 
.A(n_17073),
.Y(n_17280)
);

INVx1_ASAP7_75t_L g17281 ( 
.A(n_17094),
.Y(n_17281)
);

OR2x2_ASAP7_75t_L g17282 ( 
.A(n_16587),
.B(n_16589),
.Y(n_17282)
);

OAI211xp5_ASAP7_75t_SL g17283 ( 
.A1(n_16786),
.A2(n_11952),
.B(n_11959),
.C(n_11939),
.Y(n_17283)
);

AND2x2_ASAP7_75t_L g17284 ( 
.A(n_16831),
.B(n_11959),
.Y(n_17284)
);

OAI21x1_ASAP7_75t_L g17285 ( 
.A1(n_16727),
.A2(n_11916),
.B(n_12078),
.Y(n_17285)
);

INVx1_ASAP7_75t_L g17286 ( 
.A(n_16805),
.Y(n_17286)
);

INVx2_ASAP7_75t_L g17287 ( 
.A(n_17086),
.Y(n_17287)
);

INVx3_ASAP7_75t_L g17288 ( 
.A(n_17086),
.Y(n_17288)
);

AND2x2_ASAP7_75t_L g17289 ( 
.A(n_16590),
.B(n_9434),
.Y(n_17289)
);

NAND3xp33_ASAP7_75t_L g17290 ( 
.A(n_16571),
.B(n_10542),
.C(n_10539),
.Y(n_17290)
);

NAND2xp5_ASAP7_75t_L g17291 ( 
.A(n_16681),
.B(n_9578),
.Y(n_17291)
);

NAND2xp5_ASAP7_75t_L g17292 ( 
.A(n_16683),
.B(n_9578),
.Y(n_17292)
);

OR2x2_ASAP7_75t_L g17293 ( 
.A(n_16595),
.B(n_9369),
.Y(n_17293)
);

OR2x2_ASAP7_75t_L g17294 ( 
.A(n_16618),
.B(n_9321),
.Y(n_17294)
);

INVx1_ASAP7_75t_L g17295 ( 
.A(n_16558),
.Y(n_17295)
);

AND2x2_ASAP7_75t_L g17296 ( 
.A(n_16985),
.B(n_9294),
.Y(n_17296)
);

AND2x2_ASAP7_75t_L g17297 ( 
.A(n_17000),
.B(n_9294),
.Y(n_17297)
);

INVx1_ASAP7_75t_L g17298 ( 
.A(n_16564),
.Y(n_17298)
);

INVx1_ASAP7_75t_L g17299 ( 
.A(n_16908),
.Y(n_17299)
);

NAND2xp5_ASAP7_75t_L g17300 ( 
.A(n_17027),
.B(n_16650),
.Y(n_17300)
);

CKINVDCx5p33_ASAP7_75t_R g17301 ( 
.A(n_17035),
.Y(n_17301)
);

INVx1_ASAP7_75t_L g17302 ( 
.A(n_16631),
.Y(n_17302)
);

INVxp67_ASAP7_75t_L g17303 ( 
.A(n_16872),
.Y(n_17303)
);

INVx1_ASAP7_75t_SL g17304 ( 
.A(n_16547),
.Y(n_17304)
);

INVx2_ASAP7_75t_L g17305 ( 
.A(n_17011),
.Y(n_17305)
);

OR2x2_ASAP7_75t_L g17306 ( 
.A(n_16549),
.B(n_9321),
.Y(n_17306)
);

INVx1_ASAP7_75t_L g17307 ( 
.A(n_16607),
.Y(n_17307)
);

AND2x2_ASAP7_75t_L g17308 ( 
.A(n_17040),
.B(n_9294),
.Y(n_17308)
);

INVx1_ASAP7_75t_L g17309 ( 
.A(n_16577),
.Y(n_17309)
);

AND2x2_ASAP7_75t_L g17310 ( 
.A(n_16588),
.B(n_9294),
.Y(n_17310)
);

INVx1_ASAP7_75t_SL g17311 ( 
.A(n_16610),
.Y(n_17311)
);

AND2x2_ASAP7_75t_L g17312 ( 
.A(n_16605),
.B(n_9294),
.Y(n_17312)
);

HB1xp67_ASAP7_75t_L g17313 ( 
.A(n_16658),
.Y(n_17313)
);

NOR3xp33_ASAP7_75t_SL g17314 ( 
.A(n_16620),
.B(n_9470),
.C(n_9561),
.Y(n_17314)
);

AND2x2_ASAP7_75t_L g17315 ( 
.A(n_16630),
.B(n_16924),
.Y(n_17315)
);

AND2x2_ASAP7_75t_L g17316 ( 
.A(n_16663),
.B(n_9294),
.Y(n_17316)
);

NAND2xp5_ASAP7_75t_L g17317 ( 
.A(n_17082),
.B(n_17015),
.Y(n_17317)
);

AND2x4_ASAP7_75t_L g17318 ( 
.A(n_16889),
.B(n_8494),
.Y(n_17318)
);

OR2x2_ASAP7_75t_L g17319 ( 
.A(n_16611),
.B(n_9321),
.Y(n_17319)
);

OR2x2_ASAP7_75t_L g17320 ( 
.A(n_16693),
.B(n_9328),
.Y(n_17320)
);

INVx1_ASAP7_75t_L g17321 ( 
.A(n_16545),
.Y(n_17321)
);

OR2x6_ASAP7_75t_L g17322 ( 
.A(n_16710),
.B(n_10789),
.Y(n_17322)
);

NAND2xp5_ASAP7_75t_L g17323 ( 
.A(n_17016),
.B(n_9578),
.Y(n_17323)
);

INVx1_ASAP7_75t_L g17324 ( 
.A(n_16546),
.Y(n_17324)
);

INVx1_ASAP7_75t_L g17325 ( 
.A(n_16528),
.Y(n_17325)
);

INVx1_ASAP7_75t_L g17326 ( 
.A(n_16948),
.Y(n_17326)
);

AND2x2_ASAP7_75t_L g17327 ( 
.A(n_17047),
.B(n_9326),
.Y(n_17327)
);

AOI221x1_ASAP7_75t_L g17328 ( 
.A1(n_16541),
.A2(n_10709),
.B1(n_10716),
.B2(n_10700),
.C(n_10668),
.Y(n_17328)
);

OR2x2_ASAP7_75t_L g17329 ( 
.A(n_16832),
.B(n_9328),
.Y(n_17329)
);

INVx2_ASAP7_75t_SL g17330 ( 
.A(n_16863),
.Y(n_17330)
);

AND2x2_ASAP7_75t_L g17331 ( 
.A(n_16729),
.B(n_9326),
.Y(n_17331)
);

INVx2_ASAP7_75t_L g17332 ( 
.A(n_16992),
.Y(n_17332)
);

AND2x2_ASAP7_75t_L g17333 ( 
.A(n_16929),
.B(n_9326),
.Y(n_17333)
);

INVx1_ASAP7_75t_L g17334 ( 
.A(n_16796),
.Y(n_17334)
);

AND2x2_ASAP7_75t_L g17335 ( 
.A(n_16971),
.B(n_9326),
.Y(n_17335)
);

OR2x2_ASAP7_75t_L g17336 ( 
.A(n_16868),
.B(n_9328),
.Y(n_17336)
);

OR2x2_ASAP7_75t_L g17337 ( 
.A(n_16624),
.B(n_8661),
.Y(n_17337)
);

NOR3xp33_ASAP7_75t_L g17338 ( 
.A(n_16578),
.B(n_16579),
.C(n_16946),
.Y(n_17338)
);

NAND2xp5_ASAP7_75t_L g17339 ( 
.A(n_17051),
.B(n_9578),
.Y(n_17339)
);

NAND2xp5_ASAP7_75t_L g17340 ( 
.A(n_16812),
.B(n_9463),
.Y(n_17340)
);

NAND2xp5_ASAP7_75t_L g17341 ( 
.A(n_16859),
.B(n_16950),
.Y(n_17341)
);

INVx1_ASAP7_75t_L g17342 ( 
.A(n_17002),
.Y(n_17342)
);

AND2x2_ASAP7_75t_L g17343 ( 
.A(n_16982),
.B(n_9326),
.Y(n_17343)
);

INVx2_ASAP7_75t_L g17344 ( 
.A(n_17008),
.Y(n_17344)
);

NAND2xp5_ASAP7_75t_SL g17345 ( 
.A(n_16855),
.B(n_10539),
.Y(n_17345)
);

NAND2xp5_ASAP7_75t_L g17346 ( 
.A(n_16758),
.B(n_9463),
.Y(n_17346)
);

AND2x2_ASAP7_75t_L g17347 ( 
.A(n_17057),
.B(n_9326),
.Y(n_17347)
);

AND2x2_ASAP7_75t_L g17348 ( 
.A(n_16659),
.B(n_9382),
.Y(n_17348)
);

NOR2xp33_ASAP7_75t_R g17349 ( 
.A(n_16884),
.B(n_7703),
.Y(n_17349)
);

AND2x2_ASAP7_75t_L g17350 ( 
.A(n_16695),
.B(n_9382),
.Y(n_17350)
);

OR2x2_ASAP7_75t_L g17351 ( 
.A(n_16999),
.B(n_8661),
.Y(n_17351)
);

NAND2xp5_ASAP7_75t_L g17352 ( 
.A(n_17055),
.B(n_10524),
.Y(n_17352)
);

INVx1_ASAP7_75t_L g17353 ( 
.A(n_16705),
.Y(n_17353)
);

AND2x2_ASAP7_75t_L g17354 ( 
.A(n_16699),
.B(n_9382),
.Y(n_17354)
);

AND2x2_ASAP7_75t_L g17355 ( 
.A(n_16668),
.B(n_9382),
.Y(n_17355)
);

NAND2xp5_ASAP7_75t_L g17356 ( 
.A(n_17059),
.B(n_10524),
.Y(n_17356)
);

AND2x2_ASAP7_75t_L g17357 ( 
.A(n_16672),
.B(n_9382),
.Y(n_17357)
);

INVxp67_ASAP7_75t_SL g17358 ( 
.A(n_16584),
.Y(n_17358)
);

INVx1_ASAP7_75t_L g17359 ( 
.A(n_16692),
.Y(n_17359)
);

INVx2_ASAP7_75t_L g17360 ( 
.A(n_17037),
.Y(n_17360)
);

NOR3xp33_ASAP7_75t_L g17361 ( 
.A(n_16764),
.B(n_10700),
.C(n_10668),
.Y(n_17361)
);

HB1xp67_ASAP7_75t_L g17362 ( 
.A(n_16967),
.Y(n_17362)
);

INVx2_ASAP7_75t_L g17363 ( 
.A(n_16602),
.Y(n_17363)
);

INVx2_ASAP7_75t_L g17364 ( 
.A(n_16865),
.Y(n_17364)
);

OR2x2_ASAP7_75t_L g17365 ( 
.A(n_16621),
.B(n_8680),
.Y(n_17365)
);

AND2x4_ASAP7_75t_SL g17366 ( 
.A(n_16858),
.B(n_7703),
.Y(n_17366)
);

INVx1_ASAP7_75t_L g17367 ( 
.A(n_17081),
.Y(n_17367)
);

AND2x2_ASAP7_75t_L g17368 ( 
.A(n_16912),
.B(n_9382),
.Y(n_17368)
);

AND2x2_ASAP7_75t_L g17369 ( 
.A(n_16922),
.B(n_9399),
.Y(n_17369)
);

OR2x2_ASAP7_75t_L g17370 ( 
.A(n_16843),
.B(n_8680),
.Y(n_17370)
);

INVx1_ASAP7_75t_L g17371 ( 
.A(n_16976),
.Y(n_17371)
);

BUFx3_ASAP7_75t_L g17372 ( 
.A(n_16823),
.Y(n_17372)
);

INVx2_ASAP7_75t_L g17373 ( 
.A(n_16792),
.Y(n_17373)
);

INVx1_ASAP7_75t_L g17374 ( 
.A(n_16550),
.Y(n_17374)
);

INVx1_ASAP7_75t_L g17375 ( 
.A(n_16713),
.Y(n_17375)
);

INVx1_ASAP7_75t_L g17376 ( 
.A(n_16747),
.Y(n_17376)
);

AND2x2_ASAP7_75t_L g17377 ( 
.A(n_16762),
.B(n_9399),
.Y(n_17377)
);

AND2x2_ASAP7_75t_L g17378 ( 
.A(n_16763),
.B(n_16806),
.Y(n_17378)
);

AND2x2_ASAP7_75t_L g17379 ( 
.A(n_16757),
.B(n_9399),
.Y(n_17379)
);

NAND2xp5_ASAP7_75t_L g17380 ( 
.A(n_17062),
.B(n_10526),
.Y(n_17380)
);

AOI222xp33_ASAP7_75t_L g17381 ( 
.A1(n_16582),
.A2(n_10771),
.B1(n_10748),
.B2(n_10752),
.C1(n_10745),
.C2(n_10716),
.Y(n_17381)
);

NAND2xp5_ASAP7_75t_L g17382 ( 
.A(n_17063),
.B(n_10528),
.Y(n_17382)
);

NOR2xp33_ASAP7_75t_L g17383 ( 
.A(n_17043),
.B(n_10539),
.Y(n_17383)
);

INVx1_ASAP7_75t_L g17384 ( 
.A(n_17078),
.Y(n_17384)
);

AND2x4_ASAP7_75t_L g17385 ( 
.A(n_16708),
.B(n_8494),
.Y(n_17385)
);

AND2x4_ASAP7_75t_L g17386 ( 
.A(n_16775),
.B(n_8494),
.Y(n_17386)
);

NAND2xp5_ASAP7_75t_L g17387 ( 
.A(n_17068),
.B(n_10528),
.Y(n_17387)
);

AND2x2_ASAP7_75t_L g17388 ( 
.A(n_16902),
.B(n_9399),
.Y(n_17388)
);

AND2x2_ASAP7_75t_SL g17389 ( 
.A(n_16994),
.B(n_10542),
.Y(n_17389)
);

INVx2_ASAP7_75t_L g17390 ( 
.A(n_16787),
.Y(n_17390)
);

INVxp67_ASAP7_75t_SL g17391 ( 
.A(n_16895),
.Y(n_17391)
);

INVx2_ASAP7_75t_L g17392 ( 
.A(n_16802),
.Y(n_17392)
);

INVx1_ASAP7_75t_L g17393 ( 
.A(n_16901),
.Y(n_17393)
);

NOR2xp33_ASAP7_75t_L g17394 ( 
.A(n_16781),
.B(n_10542),
.Y(n_17394)
);

OR2x2_ASAP7_75t_L g17395 ( 
.A(n_16844),
.B(n_8787),
.Y(n_17395)
);

AND2x4_ASAP7_75t_SL g17396 ( 
.A(n_16842),
.B(n_7703),
.Y(n_17396)
);

INVxp67_ASAP7_75t_SL g17397 ( 
.A(n_16850),
.Y(n_17397)
);

AOI221xp5_ASAP7_75t_L g17398 ( 
.A1(n_16532),
.A2(n_10709),
.B1(n_10716),
.B2(n_10700),
.C(n_10668),
.Y(n_17398)
);

NAND2x1_ASAP7_75t_L g17399 ( 
.A(n_16834),
.B(n_10914),
.Y(n_17399)
);

NAND2xp5_ASAP7_75t_L g17400 ( 
.A(n_17074),
.B(n_10534),
.Y(n_17400)
);

INVx1_ASAP7_75t_SL g17401 ( 
.A(n_16677),
.Y(n_17401)
);

AND2x2_ASAP7_75t_L g17402 ( 
.A(n_16904),
.B(n_16680),
.Y(n_17402)
);

AND2x2_ASAP7_75t_L g17403 ( 
.A(n_16679),
.B(n_9399),
.Y(n_17403)
);

NAND3xp33_ASAP7_75t_L g17404 ( 
.A(n_16643),
.B(n_10584),
.C(n_10542),
.Y(n_17404)
);

AND2x2_ASAP7_75t_SL g17405 ( 
.A(n_16652),
.B(n_10542),
.Y(n_17405)
);

AND2x2_ASAP7_75t_L g17406 ( 
.A(n_16742),
.B(n_9399),
.Y(n_17406)
);

AND2x2_ASAP7_75t_L g17407 ( 
.A(n_16759),
.B(n_9446),
.Y(n_17407)
);

INVx2_ASAP7_75t_SL g17408 ( 
.A(n_16804),
.Y(n_17408)
);

INVx1_ASAP7_75t_L g17409 ( 
.A(n_16921),
.Y(n_17409)
);

INVx2_ASAP7_75t_L g17410 ( 
.A(n_16822),
.Y(n_17410)
);

HB1xp67_ASAP7_75t_L g17411 ( 
.A(n_16635),
.Y(n_17411)
);

INVx2_ASAP7_75t_SL g17412 ( 
.A(n_16849),
.Y(n_17412)
);

INVx1_ASAP7_75t_L g17413 ( 
.A(n_16839),
.Y(n_17413)
);

NAND2xp5_ASAP7_75t_L g17414 ( 
.A(n_17077),
.B(n_10534),
.Y(n_17414)
);

OR2x2_ASAP7_75t_L g17415 ( 
.A(n_17014),
.B(n_8787),
.Y(n_17415)
);

AND2x2_ASAP7_75t_L g17416 ( 
.A(n_16848),
.B(n_9446),
.Y(n_17416)
);

INVx1_ASAP7_75t_L g17417 ( 
.A(n_16840),
.Y(n_17417)
);

INVxp67_ASAP7_75t_SL g17418 ( 
.A(n_17049),
.Y(n_17418)
);

AND2x2_ASAP7_75t_L g17419 ( 
.A(n_16667),
.B(n_9446),
.Y(n_17419)
);

AND2x2_ASAP7_75t_L g17420 ( 
.A(n_16877),
.B(n_9446),
.Y(n_17420)
);

INVx1_ASAP7_75t_L g17421 ( 
.A(n_17032),
.Y(n_17421)
);

INVx2_ASAP7_75t_L g17422 ( 
.A(n_16857),
.Y(n_17422)
);

NAND2xp5_ASAP7_75t_SL g17423 ( 
.A(n_16875),
.B(n_10542),
.Y(n_17423)
);

NAND2xp5_ASAP7_75t_L g17424 ( 
.A(n_16861),
.B(n_10541),
.Y(n_17424)
);

INVx1_ASAP7_75t_L g17425 ( 
.A(n_16932),
.Y(n_17425)
);

INVx1_ASAP7_75t_SL g17426 ( 
.A(n_16722),
.Y(n_17426)
);

NAND2xp5_ASAP7_75t_SL g17427 ( 
.A(n_16653),
.B(n_10584),
.Y(n_17427)
);

INVx1_ASAP7_75t_L g17428 ( 
.A(n_16718),
.Y(n_17428)
);

INVx1_ASAP7_75t_L g17429 ( 
.A(n_16928),
.Y(n_17429)
);

INVx2_ASAP7_75t_L g17430 ( 
.A(n_16862),
.Y(n_17430)
);

NAND2xp5_ASAP7_75t_L g17431 ( 
.A(n_16815),
.B(n_10541),
.Y(n_17431)
);

NOR2xp33_ASAP7_75t_L g17432 ( 
.A(n_17088),
.B(n_10584),
.Y(n_17432)
);

NOR3xp33_ASAP7_75t_L g17433 ( 
.A(n_17091),
.B(n_10720),
.C(n_10709),
.Y(n_17433)
);

INVx1_ASAP7_75t_L g17434 ( 
.A(n_16991),
.Y(n_17434)
);

HB1xp67_ASAP7_75t_L g17435 ( 
.A(n_16873),
.Y(n_17435)
);

AND2x2_ASAP7_75t_L g17436 ( 
.A(n_16942),
.B(n_9446),
.Y(n_17436)
);

NOR2xp33_ASAP7_75t_L g17437 ( 
.A(n_17097),
.B(n_10584),
.Y(n_17437)
);

INVx1_ASAP7_75t_L g17438 ( 
.A(n_16816),
.Y(n_17438)
);

NOR2x1_ASAP7_75t_L g17439 ( 
.A(n_16529),
.B(n_8494),
.Y(n_17439)
);

AND2x2_ASAP7_75t_L g17440 ( 
.A(n_16964),
.B(n_9446),
.Y(n_17440)
);

NOR2xp33_ASAP7_75t_L g17441 ( 
.A(n_16664),
.B(n_10584),
.Y(n_17441)
);

INVx1_ASAP7_75t_L g17442 ( 
.A(n_16756),
.Y(n_17442)
);

NAND2xp5_ASAP7_75t_L g17443 ( 
.A(n_16748),
.B(n_10543),
.Y(n_17443)
);

AND2x2_ASAP7_75t_L g17444 ( 
.A(n_16965),
.B(n_16969),
.Y(n_17444)
);

AND2x2_ASAP7_75t_L g17445 ( 
.A(n_16894),
.B(n_9487),
.Y(n_17445)
);

INVx1_ASAP7_75t_L g17446 ( 
.A(n_16800),
.Y(n_17446)
);

AOI21xp5_ASAP7_75t_L g17447 ( 
.A1(n_16655),
.A2(n_12101),
.B(n_12078),
.Y(n_17447)
);

AND2x2_ASAP7_75t_L g17448 ( 
.A(n_16899),
.B(n_16777),
.Y(n_17448)
);

AND2x2_ASAP7_75t_L g17449 ( 
.A(n_16778),
.B(n_9487),
.Y(n_17449)
);

INVx1_ASAP7_75t_L g17450 ( 
.A(n_16935),
.Y(n_17450)
);

AND2x2_ASAP7_75t_L g17451 ( 
.A(n_16714),
.B(n_9487),
.Y(n_17451)
);

NAND2xp5_ASAP7_75t_L g17452 ( 
.A(n_16749),
.B(n_10543),
.Y(n_17452)
);

AND2x2_ASAP7_75t_L g17453 ( 
.A(n_16721),
.B(n_9487),
.Y(n_17453)
);

INVx1_ASAP7_75t_L g17454 ( 
.A(n_17092),
.Y(n_17454)
);

NOR2xp33_ASAP7_75t_L g17455 ( 
.A(n_17098),
.B(n_10584),
.Y(n_17455)
);

AND2x4_ASAP7_75t_L g17456 ( 
.A(n_17058),
.B(n_8514),
.Y(n_17456)
);

NAND2xp5_ASAP7_75t_L g17457 ( 
.A(n_16750),
.B(n_10550),
.Y(n_17457)
);

AND2x2_ASAP7_75t_L g17458 ( 
.A(n_16725),
.B(n_9487),
.Y(n_17458)
);

NAND2xp5_ASAP7_75t_L g17459 ( 
.A(n_16785),
.B(n_10550),
.Y(n_17459)
);

INVx1_ASAP7_75t_L g17460 ( 
.A(n_17010),
.Y(n_17460)
);

INVx1_ASAP7_75t_L g17461 ( 
.A(n_16925),
.Y(n_17461)
);

INVx1_ASAP7_75t_L g17462 ( 
.A(n_16732),
.Y(n_17462)
);

INVx2_ASAP7_75t_L g17463 ( 
.A(n_16926),
.Y(n_17463)
);

AND2x2_ASAP7_75t_L g17464 ( 
.A(n_16738),
.B(n_9487),
.Y(n_17464)
);

NOR2x1_ASAP7_75t_L g17465 ( 
.A(n_16557),
.B(n_8514),
.Y(n_17465)
);

INVx2_ASAP7_75t_L g17466 ( 
.A(n_16940),
.Y(n_17466)
);

AND2x2_ASAP7_75t_L g17467 ( 
.A(n_16741),
.B(n_9495),
.Y(n_17467)
);

INVx1_ASAP7_75t_L g17468 ( 
.A(n_16733),
.Y(n_17468)
);

INVxp67_ASAP7_75t_SL g17469 ( 
.A(n_17048),
.Y(n_17469)
);

INVx1_ASAP7_75t_L g17470 ( 
.A(n_17095),
.Y(n_17470)
);

INVx1_ASAP7_75t_L g17471 ( 
.A(n_17096),
.Y(n_17471)
);

AND2x2_ASAP7_75t_L g17472 ( 
.A(n_16745),
.B(n_9495),
.Y(n_17472)
);

AOI22xp33_ASAP7_75t_L g17473 ( 
.A1(n_17087),
.A2(n_17080),
.B1(n_16906),
.B2(n_16903),
.Y(n_17473)
);

BUFx3_ASAP7_75t_L g17474 ( 
.A(n_16852),
.Y(n_17474)
);

NOR2xp33_ASAP7_75t_L g17475 ( 
.A(n_16780),
.B(n_10659),
.Y(n_17475)
);

AND2x2_ASAP7_75t_L g17476 ( 
.A(n_16730),
.B(n_9495),
.Y(n_17476)
);

AND2x2_ASAP7_75t_L g17477 ( 
.A(n_16736),
.B(n_9495),
.Y(n_17477)
);

AND2x2_ASAP7_75t_L g17478 ( 
.A(n_16737),
.B(n_9495),
.Y(n_17478)
);

AND2x2_ASAP7_75t_L g17479 ( 
.A(n_16744),
.B(n_9495),
.Y(n_17479)
);

INVx1_ASAP7_75t_L g17480 ( 
.A(n_17099),
.Y(n_17480)
);

AOI221xp5_ASAP7_75t_L g17481 ( 
.A1(n_16968),
.A2(n_10726),
.B1(n_10720),
.B2(n_10748),
.C(n_10745),
.Y(n_17481)
);

AND2x2_ASAP7_75t_L g17482 ( 
.A(n_16746),
.B(n_9510),
.Y(n_17482)
);

INVx1_ASAP7_75t_L g17483 ( 
.A(n_17013),
.Y(n_17483)
);

AND2x4_ASAP7_75t_L g17484 ( 
.A(n_17064),
.B(n_8514),
.Y(n_17484)
);

NAND2xp5_ASAP7_75t_L g17485 ( 
.A(n_16949),
.B(n_10552),
.Y(n_17485)
);

AND2x2_ASAP7_75t_L g17486 ( 
.A(n_16779),
.B(n_9510),
.Y(n_17486)
);

INVx1_ASAP7_75t_L g17487 ( 
.A(n_16956),
.Y(n_17487)
);

AND2x4_ASAP7_75t_L g17488 ( 
.A(n_17069),
.B(n_8514),
.Y(n_17488)
);

AND2x2_ASAP7_75t_L g17489 ( 
.A(n_16782),
.B(n_9510),
.Y(n_17489)
);

AND2x2_ASAP7_75t_L g17490 ( 
.A(n_16784),
.B(n_9510),
.Y(n_17490)
);

OAI221xp5_ASAP7_75t_L g17491 ( 
.A1(n_16696),
.A2(n_10726),
.B1(n_10720),
.B2(n_10771),
.C(n_10752),
.Y(n_17491)
);

AND2x2_ASAP7_75t_L g17492 ( 
.A(n_16876),
.B(n_9510),
.Y(n_17492)
);

AND2x2_ASAP7_75t_L g17493 ( 
.A(n_16795),
.B(n_9510),
.Y(n_17493)
);

NOR2x1_ASAP7_75t_L g17494 ( 
.A(n_16648),
.B(n_8514),
.Y(n_17494)
);

INVx2_ASAP7_75t_SL g17495 ( 
.A(n_16793),
.Y(n_17495)
);

AND2x2_ASAP7_75t_L g17496 ( 
.A(n_16927),
.B(n_9531),
.Y(n_17496)
);

AND2x2_ASAP7_75t_L g17497 ( 
.A(n_16987),
.B(n_9531),
.Y(n_17497)
);

NAND2xp5_ASAP7_75t_L g17498 ( 
.A(n_16960),
.B(n_10552),
.Y(n_17498)
);

AND2x2_ASAP7_75t_L g17499 ( 
.A(n_16945),
.B(n_9531),
.Y(n_17499)
);

AND2x2_ASAP7_75t_L g17500 ( 
.A(n_16847),
.B(n_9531),
.Y(n_17500)
);

AND2x2_ASAP7_75t_L g17501 ( 
.A(n_16662),
.B(n_9531),
.Y(n_17501)
);

HB1xp67_ASAP7_75t_L g17502 ( 
.A(n_16807),
.Y(n_17502)
);

BUFx2_ASAP7_75t_L g17503 ( 
.A(n_16817),
.Y(n_17503)
);

AND2x2_ASAP7_75t_L g17504 ( 
.A(n_16947),
.B(n_9531),
.Y(n_17504)
);

INVx1_ASAP7_75t_SL g17505 ( 
.A(n_16666),
.Y(n_17505)
);

AOI211xp5_ASAP7_75t_L g17506 ( 
.A1(n_16649),
.A2(n_8634),
.B(n_9384),
.C(n_12101),
.Y(n_17506)
);

AOI222xp33_ASAP7_75t_L g17507 ( 
.A1(n_16887),
.A2(n_10726),
.B1(n_12119),
.B2(n_10666),
.C1(n_10772),
.C2(n_10682),
.Y(n_17507)
);

INVx1_ASAP7_75t_L g17508 ( 
.A(n_16980),
.Y(n_17508)
);

INVx3_ASAP7_75t_L g17509 ( 
.A(n_17005),
.Y(n_17509)
);

OR2x2_ASAP7_75t_L g17510 ( 
.A(n_16941),
.B(n_8359),
.Y(n_17510)
);

INVx1_ASAP7_75t_L g17511 ( 
.A(n_17012),
.Y(n_17511)
);

AND2x4_ASAP7_75t_L g17512 ( 
.A(n_16880),
.B(n_8542),
.Y(n_17512)
);

AND2x2_ASAP7_75t_L g17513 ( 
.A(n_17024),
.B(n_12149),
.Y(n_17513)
);

OR2x2_ASAP7_75t_L g17514 ( 
.A(n_17093),
.B(n_8386),
.Y(n_17514)
);

OR2x2_ASAP7_75t_L g17515 ( 
.A(n_17100),
.B(n_8438),
.Y(n_17515)
);

NAND5xp2_ASAP7_75t_L g17516 ( 
.A(n_16890),
.B(n_9327),
.C(n_9284),
.D(n_8686),
.E(n_9384),
.Y(n_17516)
);

NAND2xp5_ASAP7_75t_SL g17517 ( 
.A(n_16711),
.B(n_10659),
.Y(n_17517)
);

INVx2_ASAP7_75t_L g17518 ( 
.A(n_16996),
.Y(n_17518)
);

AND2x2_ASAP7_75t_L g17519 ( 
.A(n_16838),
.B(n_12149),
.Y(n_17519)
);

OR2x2_ASAP7_75t_L g17520 ( 
.A(n_16640),
.B(n_8438),
.Y(n_17520)
);

AND2x2_ASAP7_75t_L g17521 ( 
.A(n_16972),
.B(n_12177),
.Y(n_17521)
);

INVx1_ASAP7_75t_L g17522 ( 
.A(n_16687),
.Y(n_17522)
);

INVxp67_ASAP7_75t_L g17523 ( 
.A(n_16555),
.Y(n_17523)
);

AND2x2_ASAP7_75t_L g17524 ( 
.A(n_16975),
.B(n_12177),
.Y(n_17524)
);

INVxp67_ASAP7_75t_L g17525 ( 
.A(n_16556),
.Y(n_17525)
);

OAI33xp33_ASAP7_75t_L g17526 ( 
.A1(n_16825),
.A2(n_10565),
.A3(n_10558),
.B1(n_10571),
.B2(n_10569),
.B3(n_10560),
.Y(n_17526)
);

OR2x2_ASAP7_75t_L g17527 ( 
.A(n_16851),
.B(n_8570),
.Y(n_17527)
);

HB1xp67_ASAP7_75t_L g17528 ( 
.A(n_16881),
.Y(n_17528)
);

INVx2_ASAP7_75t_L g17529 ( 
.A(n_16997),
.Y(n_17529)
);

INVx1_ASAP7_75t_L g17530 ( 
.A(n_16761),
.Y(n_17530)
);

NAND4xp25_ASAP7_75t_L g17531 ( 
.A(n_17022),
.B(n_16690),
.C(n_16751),
.D(n_16688),
.Y(n_17531)
);

INVx1_ASAP7_75t_L g17532 ( 
.A(n_16773),
.Y(n_17532)
);

AND2x2_ASAP7_75t_L g17533 ( 
.A(n_16914),
.B(n_12218),
.Y(n_17533)
);

INVx1_ASAP7_75t_L g17534 ( 
.A(n_16774),
.Y(n_17534)
);

INVx1_ASAP7_75t_SL g17535 ( 
.A(n_16766),
.Y(n_17535)
);

INVx2_ASAP7_75t_L g17536 ( 
.A(n_16998),
.Y(n_17536)
);

OAI33xp33_ASAP7_75t_L g17537 ( 
.A1(n_16665),
.A2(n_10565),
.A3(n_10558),
.B1(n_10571),
.B2(n_10569),
.B3(n_10560),
.Y(n_17537)
);

INVx1_ASAP7_75t_L g17538 ( 
.A(n_16776),
.Y(n_17538)
);

HB1xp67_ASAP7_75t_L g17539 ( 
.A(n_16891),
.Y(n_17539)
);

AND2x2_ASAP7_75t_L g17540 ( 
.A(n_16915),
.B(n_12218),
.Y(n_17540)
);

AND2x2_ASAP7_75t_SL g17541 ( 
.A(n_16769),
.B(n_10659),
.Y(n_17541)
);

BUFx2_ASAP7_75t_L g17542 ( 
.A(n_16670),
.Y(n_17542)
);

INVx1_ASAP7_75t_L g17543 ( 
.A(n_16798),
.Y(n_17543)
);

BUFx2_ASAP7_75t_SL g17544 ( 
.A(n_16818),
.Y(n_17544)
);

AND2x2_ASAP7_75t_L g17545 ( 
.A(n_17030),
.B(n_12251),
.Y(n_17545)
);

OR2x2_ASAP7_75t_L g17546 ( 
.A(n_17061),
.B(n_8570),
.Y(n_17546)
);

INVx1_ASAP7_75t_L g17547 ( 
.A(n_16808),
.Y(n_17547)
);

INVx1_ASAP7_75t_L g17548 ( 
.A(n_16820),
.Y(n_17548)
);

AND2x2_ASAP7_75t_L g17549 ( 
.A(n_17053),
.B(n_12251),
.Y(n_17549)
);

AND2x2_ASAP7_75t_L g17550 ( 
.A(n_16933),
.B(n_8542),
.Y(n_17550)
);

NAND2xp5_ASAP7_75t_L g17551 ( 
.A(n_17085),
.B(n_10575),
.Y(n_17551)
);

AOI22xp33_ASAP7_75t_L g17552 ( 
.A1(n_16882),
.A2(n_8675),
.B1(n_8767),
.B2(n_8498),
.Y(n_17552)
);

OR2x2_ASAP7_75t_L g17553 ( 
.A(n_17070),
.B(n_8612),
.Y(n_17553)
);

AND2x2_ASAP7_75t_L g17554 ( 
.A(n_16905),
.B(n_8542),
.Y(n_17554)
);

OR2x2_ASAP7_75t_L g17555 ( 
.A(n_17072),
.B(n_8612),
.Y(n_17555)
);

INVx1_ASAP7_75t_L g17556 ( 
.A(n_16827),
.Y(n_17556)
);

NAND2xp5_ASAP7_75t_L g17557 ( 
.A(n_17090),
.B(n_10575),
.Y(n_17557)
);

AND2x2_ASAP7_75t_L g17558 ( 
.A(n_16920),
.B(n_17079),
.Y(n_17558)
);

AND2x2_ASAP7_75t_L g17559 ( 
.A(n_16824),
.B(n_8542),
.Y(n_17559)
);

AND2x2_ASAP7_75t_L g17560 ( 
.A(n_16829),
.B(n_8542),
.Y(n_17560)
);

NAND2xp5_ASAP7_75t_L g17561 ( 
.A(n_17007),
.B(n_10576),
.Y(n_17561)
);

INVx4_ASAP7_75t_L g17562 ( 
.A(n_16931),
.Y(n_17562)
);

INVx1_ASAP7_75t_L g17563 ( 
.A(n_16833),
.Y(n_17563)
);

INVx1_ASAP7_75t_L g17564 ( 
.A(n_16993),
.Y(n_17564)
);

AND2x2_ASAP7_75t_L g17565 ( 
.A(n_16870),
.B(n_10659),
.Y(n_17565)
);

INVx1_ASAP7_75t_L g17566 ( 
.A(n_17025),
.Y(n_17566)
);

AND2x2_ASAP7_75t_L g17567 ( 
.A(n_16879),
.B(n_10659),
.Y(n_17567)
);

INVx1_ASAP7_75t_L g17568 ( 
.A(n_17009),
.Y(n_17568)
);

NAND2xp5_ASAP7_75t_L g17569 ( 
.A(n_16898),
.B(n_10576),
.Y(n_17569)
);

OR2x6_ASAP7_75t_L g17570 ( 
.A(n_16897),
.B(n_10789),
.Y(n_17570)
);

INVx1_ASAP7_75t_L g17571 ( 
.A(n_16966),
.Y(n_17571)
);

AND2x2_ASAP7_75t_L g17572 ( 
.A(n_16883),
.B(n_10659),
.Y(n_17572)
);

OR2x2_ASAP7_75t_L g17573 ( 
.A(n_16694),
.B(n_8677),
.Y(n_17573)
);

AND2x2_ASAP7_75t_L g17574 ( 
.A(n_16900),
.B(n_10666),
.Y(n_17574)
);

AND2x2_ASAP7_75t_L g17575 ( 
.A(n_16970),
.B(n_10666),
.Y(n_17575)
);

NAND2xp5_ASAP7_75t_L g17576 ( 
.A(n_17039),
.B(n_10577),
.Y(n_17576)
);

HB1xp67_ASAP7_75t_L g17577 ( 
.A(n_16703),
.Y(n_17577)
);

AND2x2_ASAP7_75t_L g17578 ( 
.A(n_16978),
.B(n_10666),
.Y(n_17578)
);

OAI21xp33_ASAP7_75t_L g17579 ( 
.A1(n_17019),
.A2(n_9055),
.B(n_8871),
.Y(n_17579)
);

OAI211xp5_ASAP7_75t_L g17580 ( 
.A1(n_16938),
.A2(n_8634),
.B(n_12119),
.C(n_10682),
.Y(n_17580)
);

AND2x2_ASAP7_75t_L g17581 ( 
.A(n_16939),
.B(n_10666),
.Y(n_17581)
);

NAND2xp33_ASAP7_75t_R g17582 ( 
.A(n_16739),
.B(n_9252),
.Y(n_17582)
);

AND2x2_ASAP7_75t_L g17583 ( 
.A(n_16953),
.B(n_10666),
.Y(n_17583)
);

INVx2_ASAP7_75t_L g17584 ( 
.A(n_17084),
.Y(n_17584)
);

INVx1_ASAP7_75t_L g17585 ( 
.A(n_17028),
.Y(n_17585)
);

INVx2_ASAP7_75t_L g17586 ( 
.A(n_16962),
.Y(n_17586)
);

OR2x2_ASAP7_75t_L g17587 ( 
.A(n_16864),
.B(n_8677),
.Y(n_17587)
);

INVx1_ASAP7_75t_L g17588 ( 
.A(n_16944),
.Y(n_17588)
);

AND2x2_ASAP7_75t_L g17589 ( 
.A(n_16958),
.B(n_16961),
.Y(n_17589)
);

INVx1_ASAP7_75t_L g17590 ( 
.A(n_16955),
.Y(n_17590)
);

NAND2xp5_ASAP7_75t_L g17591 ( 
.A(n_17029),
.B(n_10577),
.Y(n_17591)
);

AND2x2_ASAP7_75t_L g17592 ( 
.A(n_16907),
.B(n_10682),
.Y(n_17592)
);

AND2x2_ASAP7_75t_L g17593 ( 
.A(n_16910),
.B(n_10682),
.Y(n_17593)
);

INVx1_ASAP7_75t_SL g17594 ( 
.A(n_16856),
.Y(n_17594)
);

OR2x2_ASAP7_75t_L g17595 ( 
.A(n_16826),
.B(n_8738),
.Y(n_17595)
);

HB1xp67_ASAP7_75t_L g17596 ( 
.A(n_16772),
.Y(n_17596)
);

AND2x2_ASAP7_75t_L g17597 ( 
.A(n_16911),
.B(n_10682),
.Y(n_17597)
);

BUFx3_ASAP7_75t_L g17598 ( 
.A(n_16916),
.Y(n_17598)
);

OR2x2_ASAP7_75t_L g17599 ( 
.A(n_16814),
.B(n_8738),
.Y(n_17599)
);

NAND2x1p5_ASAP7_75t_L g17600 ( 
.A(n_16917),
.B(n_8955),
.Y(n_17600)
);

OR2x2_ASAP7_75t_L g17601 ( 
.A(n_16821),
.B(n_8854),
.Y(n_17601)
);

INVx1_ASAP7_75t_L g17602 ( 
.A(n_17045),
.Y(n_17602)
);

INVx2_ASAP7_75t_L g17603 ( 
.A(n_17020),
.Y(n_17603)
);

NAND2xp5_ASAP7_75t_L g17604 ( 
.A(n_17056),
.B(n_10589),
.Y(n_17604)
);

NAND2x1p5_ASAP7_75t_L g17605 ( 
.A(n_16707),
.B(n_8955),
.Y(n_17605)
);

NAND2x1_ASAP7_75t_SL g17606 ( 
.A(n_17038),
.B(n_16809),
.Y(n_17606)
);

AND2x2_ASAP7_75t_L g17607 ( 
.A(n_16984),
.B(n_16765),
.Y(n_17607)
);

AND2x2_ASAP7_75t_L g17608 ( 
.A(n_16986),
.B(n_10682),
.Y(n_17608)
);

INVx1_ASAP7_75t_L g17609 ( 
.A(n_17052),
.Y(n_17609)
);

AND2x2_ASAP7_75t_L g17610 ( 
.A(n_16896),
.B(n_10772),
.Y(n_17610)
);

NAND2xp5_ASAP7_75t_L g17611 ( 
.A(n_17060),
.B(n_10589),
.Y(n_17611)
);

NAND2xp5_ASAP7_75t_L g17612 ( 
.A(n_17066),
.B(n_17067),
.Y(n_17612)
);

INVx1_ASAP7_75t_SL g17613 ( 
.A(n_16760),
.Y(n_17613)
);

AOI33xp33_ASAP7_75t_L g17614 ( 
.A1(n_16811),
.A2(n_7111),
.A3(n_7060),
.B1(n_7127),
.B2(n_7117),
.B3(n_7084),
.Y(n_17614)
);

HB1xp67_ASAP7_75t_L g17615 ( 
.A(n_17004),
.Y(n_17615)
);

INVx1_ASAP7_75t_L g17616 ( 
.A(n_16771),
.Y(n_17616)
);

INVx2_ASAP7_75t_L g17617 ( 
.A(n_16860),
.Y(n_17617)
);

INVx2_ASAP7_75t_L g17618 ( 
.A(n_17046),
.Y(n_17618)
);

INVx2_ASAP7_75t_L g17619 ( 
.A(n_17054),
.Y(n_17619)
);

INVx2_ASAP7_75t_L g17620 ( 
.A(n_17076),
.Y(n_17620)
);

NAND2xp5_ASAP7_75t_L g17621 ( 
.A(n_16837),
.B(n_16799),
.Y(n_17621)
);

AND2x4_ASAP7_75t_L g17622 ( 
.A(n_16951),
.B(n_8871),
.Y(n_17622)
);

AND2x2_ASAP7_75t_L g17623 ( 
.A(n_17023),
.B(n_10772),
.Y(n_17623)
);

AND2x2_ASAP7_75t_L g17624 ( 
.A(n_16930),
.B(n_10772),
.Y(n_17624)
);

INVx3_ASAP7_75t_L g17625 ( 
.A(n_17033),
.Y(n_17625)
);

INVx1_ASAP7_75t_L g17626 ( 
.A(n_16794),
.Y(n_17626)
);

AO21x2_ASAP7_75t_L g17627 ( 
.A1(n_17075),
.A2(n_10588),
.B(n_10502),
.Y(n_17627)
);

INVx1_ASAP7_75t_L g17628 ( 
.A(n_16801),
.Y(n_17628)
);

INVx2_ASAP7_75t_L g17629 ( 
.A(n_17034),
.Y(n_17629)
);

OAI21xp5_ASAP7_75t_L g17630 ( 
.A1(n_16697),
.A2(n_10588),
.B(n_10502),
.Y(n_17630)
);

AND2x2_ASAP7_75t_L g17631 ( 
.A(n_16995),
.B(n_10772),
.Y(n_17631)
);

AND2x4_ASAP7_75t_L g17632 ( 
.A(n_16871),
.B(n_10772),
.Y(n_17632)
);

NAND2xp5_ASAP7_75t_L g17633 ( 
.A(n_16803),
.B(n_10592),
.Y(n_17633)
);

BUFx3_ASAP7_75t_L g17634 ( 
.A(n_16841),
.Y(n_17634)
);

OR2x2_ASAP7_75t_L g17635 ( 
.A(n_16846),
.B(n_8854),
.Y(n_17635)
);

AOI22xp33_ASAP7_75t_L g17636 ( 
.A1(n_16893),
.A2(n_8675),
.B1(n_8767),
.B2(n_8498),
.Y(n_17636)
);

OR2x2_ASAP7_75t_L g17637 ( 
.A(n_16731),
.B(n_8938),
.Y(n_17637)
);

INVx2_ASAP7_75t_L g17638 ( 
.A(n_17031),
.Y(n_17638)
);

NAND2xp5_ASAP7_75t_L g17639 ( 
.A(n_17050),
.B(n_10592),
.Y(n_17639)
);

INVx1_ASAP7_75t_SL g17640 ( 
.A(n_16752),
.Y(n_17640)
);

A2O1A1Ixp33_ASAP7_75t_L g17641 ( 
.A1(n_17178),
.A2(n_16888),
.B(n_16892),
.C(n_16867),
.Y(n_17641)
);

OAI322xp33_ASAP7_75t_L g17642 ( 
.A1(n_17119),
.A2(n_16753),
.A3(n_16716),
.B1(n_16754),
.B2(n_16728),
.C1(n_16674),
.C2(n_16919),
.Y(n_17642)
);

INVx1_ASAP7_75t_L g17643 ( 
.A(n_17107),
.Y(n_17643)
);

AND2x4_ASAP7_75t_L g17644 ( 
.A(n_17130),
.B(n_16981),
.Y(n_17644)
);

HB1xp67_ASAP7_75t_L g17645 ( 
.A(n_17114),
.Y(n_17645)
);

OR2x6_ASAP7_75t_L g17646 ( 
.A(n_17544),
.B(n_16983),
.Y(n_17646)
);

INVx2_ASAP7_75t_SL g17647 ( 
.A(n_17606),
.Y(n_17647)
);

NAND2xp5_ASAP7_75t_L g17648 ( 
.A(n_17106),
.B(n_16988),
.Y(n_17648)
);

INVx1_ASAP7_75t_L g17649 ( 
.A(n_17137),
.Y(n_17649)
);

INVx1_ASAP7_75t_L g17650 ( 
.A(n_17411),
.Y(n_17650)
);

OR2x2_ASAP7_75t_L g17651 ( 
.A(n_17212),
.B(n_8938),
.Y(n_17651)
);

HB1xp67_ASAP7_75t_L g17652 ( 
.A(n_17129),
.Y(n_17652)
);

NOR2x1_ASAP7_75t_L g17653 ( 
.A(n_17147),
.B(n_10799),
.Y(n_17653)
);

AND2x4_ASAP7_75t_SL g17654 ( 
.A(n_17200),
.B(n_7703),
.Y(n_17654)
);

OR2x2_ASAP7_75t_L g17655 ( 
.A(n_17304),
.B(n_9044),
.Y(n_17655)
);

NAND2xp5_ASAP7_75t_L g17656 ( 
.A(n_17378),
.B(n_10597),
.Y(n_17656)
);

AOI22xp5_ASAP7_75t_L g17657 ( 
.A1(n_17204),
.A2(n_10732),
.B1(n_10664),
.B2(n_10799),
.Y(n_17657)
);

NAND2xp5_ASAP7_75t_L g17658 ( 
.A(n_17311),
.B(n_10597),
.Y(n_17658)
);

INVx1_ASAP7_75t_L g17659 ( 
.A(n_17313),
.Y(n_17659)
);

AOI22xp5_ASAP7_75t_L g17660 ( 
.A1(n_17301),
.A2(n_10732),
.B1(n_10664),
.B2(n_10799),
.Y(n_17660)
);

INVx1_ASAP7_75t_L g17661 ( 
.A(n_17126),
.Y(n_17661)
);

INVx2_ASAP7_75t_SL g17662 ( 
.A(n_17273),
.Y(n_17662)
);

INVx2_ASAP7_75t_L g17663 ( 
.A(n_17197),
.Y(n_17663)
);

AOI33xp33_ASAP7_75t_L g17664 ( 
.A1(n_17253),
.A2(n_17133),
.A3(n_17262),
.B1(n_17233),
.B2(n_17118),
.B3(n_17473),
.Y(n_17664)
);

OAI21xp33_ASAP7_75t_L g17665 ( 
.A1(n_17158),
.A2(n_9055),
.B(n_8871),
.Y(n_17665)
);

BUFx2_ASAP7_75t_L g17666 ( 
.A(n_17108),
.Y(n_17666)
);

INVx1_ASAP7_75t_L g17667 ( 
.A(n_17171),
.Y(n_17667)
);

AOI22xp33_ASAP7_75t_L g17668 ( 
.A1(n_17190),
.A2(n_8498),
.B1(n_8767),
.B2(n_8675),
.Y(n_17668)
);

OAI21xp5_ASAP7_75t_SL g17669 ( 
.A1(n_17216),
.A2(n_8687),
.B(n_8686),
.Y(n_17669)
);

AOI32xp33_ASAP7_75t_L g17670 ( 
.A1(n_17167),
.A2(n_10594),
.A3(n_10721),
.B1(n_10683),
.B2(n_10678),
.Y(n_17670)
);

INVx1_ASAP7_75t_L g17671 ( 
.A(n_17528),
.Y(n_17671)
);

INVx1_ASAP7_75t_SL g17672 ( 
.A(n_17259),
.Y(n_17672)
);

OA222x2_ASAP7_75t_L g17673 ( 
.A1(n_17454),
.A2(n_9230),
.B1(n_9055),
.B2(n_9298),
.C1(n_9186),
.C2(n_8871),
.Y(n_17673)
);

AOI22xp5_ASAP7_75t_L g17674 ( 
.A1(n_17582),
.A2(n_10732),
.B1(n_10664),
.B2(n_10799),
.Y(n_17674)
);

OAI33xp33_ASAP7_75t_L g17675 ( 
.A1(n_17157),
.A2(n_17102),
.A3(n_17214),
.B1(n_17207),
.B2(n_17138),
.B3(n_17299),
.Y(n_17675)
);

INVx1_ASAP7_75t_L g17676 ( 
.A(n_17539),
.Y(n_17676)
);

AND2x4_ASAP7_75t_L g17677 ( 
.A(n_17141),
.B(n_10799),
.Y(n_17677)
);

INVx1_ASAP7_75t_L g17678 ( 
.A(n_17503),
.Y(n_17678)
);

AOI32xp33_ASAP7_75t_L g17679 ( 
.A1(n_17103),
.A2(n_10594),
.A3(n_10721),
.B1(n_10683),
.B2(n_10678),
.Y(n_17679)
);

INVx2_ASAP7_75t_L g17680 ( 
.A(n_17151),
.Y(n_17680)
);

INVx2_ASAP7_75t_L g17681 ( 
.A(n_17123),
.Y(n_17681)
);

INVx1_ASAP7_75t_L g17682 ( 
.A(n_17503),
.Y(n_17682)
);

INVx1_ASAP7_75t_L g17683 ( 
.A(n_17542),
.Y(n_17683)
);

OA222x2_ASAP7_75t_L g17684 ( 
.A1(n_17372),
.A2(n_17110),
.B1(n_17474),
.B2(n_17598),
.C1(n_17250),
.C2(n_17219),
.Y(n_17684)
);

NAND2xp5_ASAP7_75t_L g17685 ( 
.A(n_17166),
.B(n_10598),
.Y(n_17685)
);

HB1xp67_ASAP7_75t_L g17686 ( 
.A(n_17235),
.Y(n_17686)
);

INVx2_ASAP7_75t_L g17687 ( 
.A(n_17322),
.Y(n_17687)
);

INVx1_ASAP7_75t_L g17688 ( 
.A(n_17542),
.Y(n_17688)
);

INVx2_ASAP7_75t_SL g17689 ( 
.A(n_17315),
.Y(n_17689)
);

AND2x2_ASAP7_75t_L g17690 ( 
.A(n_17155),
.B(n_10799),
.Y(n_17690)
);

AND2x2_ASAP7_75t_L g17691 ( 
.A(n_17127),
.B(n_10864),
.Y(n_17691)
);

INVx1_ASAP7_75t_L g17692 ( 
.A(n_17144),
.Y(n_17692)
);

NAND4xp75_ASAP7_75t_L g17693 ( 
.A(n_17125),
.B(n_9489),
.C(n_9194),
.D(n_9215),
.Y(n_17693)
);

OR2x2_ASAP7_75t_L g17694 ( 
.A(n_17535),
.B(n_9044),
.Y(n_17694)
);

AOI22xp5_ASAP7_75t_L g17695 ( 
.A1(n_17188),
.A2(n_10732),
.B1(n_10664),
.B2(n_10864),
.Y(n_17695)
);

AND2x4_ASAP7_75t_SL g17696 ( 
.A(n_17111),
.B(n_9143),
.Y(n_17696)
);

NAND2xp5_ASAP7_75t_L g17697 ( 
.A(n_17164),
.B(n_10598),
.Y(n_17697)
);

INVx1_ASAP7_75t_L g17698 ( 
.A(n_17132),
.Y(n_17698)
);

OA222x2_ASAP7_75t_L g17699 ( 
.A1(n_17170),
.A2(n_9298),
.B1(n_9186),
.B2(n_9325),
.C1(n_9230),
.C2(n_9055),
.Y(n_17699)
);

NOR2xp67_ASAP7_75t_L g17700 ( 
.A(n_17165),
.B(n_9143),
.Y(n_17700)
);

INVx1_ASAP7_75t_L g17701 ( 
.A(n_17134),
.Y(n_17701)
);

INVx2_ASAP7_75t_SL g17702 ( 
.A(n_17154),
.Y(n_17702)
);

AND2x2_ASAP7_75t_L g17703 ( 
.A(n_17105),
.B(n_17122),
.Y(n_17703)
);

INVx1_ASAP7_75t_L g17704 ( 
.A(n_17136),
.Y(n_17704)
);

AOI32xp33_ASAP7_75t_L g17705 ( 
.A1(n_17215),
.A2(n_10594),
.A3(n_10721),
.B1(n_10683),
.B2(n_10678),
.Y(n_17705)
);

INVx1_ASAP7_75t_L g17706 ( 
.A(n_17148),
.Y(n_17706)
);

INVx2_ASAP7_75t_L g17707 ( 
.A(n_17322),
.Y(n_17707)
);

OR2x2_ASAP7_75t_L g17708 ( 
.A(n_17139),
.B(n_9160),
.Y(n_17708)
);

AOI322xp5_ASAP7_75t_L g17709 ( 
.A1(n_17435),
.A2(n_9273),
.A3(n_9127),
.B1(n_9340),
.B2(n_9293),
.C1(n_8993),
.C2(n_7041),
.Y(n_17709)
);

NOR2xp33_ASAP7_75t_L g17710 ( 
.A(n_17562),
.B(n_10864),
.Y(n_17710)
);

INVx2_ASAP7_75t_L g17711 ( 
.A(n_17184),
.Y(n_17711)
);

INVx1_ASAP7_75t_L g17712 ( 
.A(n_17159),
.Y(n_17712)
);

AND2x2_ASAP7_75t_L g17713 ( 
.A(n_17222),
.B(n_10864),
.Y(n_17713)
);

AOI22xp33_ASAP7_75t_L g17714 ( 
.A1(n_17640),
.A2(n_8498),
.B1(n_8767),
.B2(n_8675),
.Y(n_17714)
);

HB1xp67_ASAP7_75t_L g17715 ( 
.A(n_17189),
.Y(n_17715)
);

INVx1_ASAP7_75t_L g17716 ( 
.A(n_17260),
.Y(n_17716)
);

INVx1_ASAP7_75t_L g17717 ( 
.A(n_17242),
.Y(n_17717)
);

OR2x2_ASAP7_75t_L g17718 ( 
.A(n_17145),
.B(n_9160),
.Y(n_17718)
);

INVx1_ASAP7_75t_L g17719 ( 
.A(n_17109),
.Y(n_17719)
);

INVxp67_ASAP7_75t_SL g17720 ( 
.A(n_17220),
.Y(n_17720)
);

OAI211xp5_ASAP7_75t_L g17721 ( 
.A1(n_17143),
.A2(n_17418),
.B(n_17397),
.C(n_17391),
.Y(n_17721)
);

INVx2_ASAP7_75t_SL g17722 ( 
.A(n_17249),
.Y(n_17722)
);

INVx1_ASAP7_75t_L g17723 ( 
.A(n_17176),
.Y(n_17723)
);

OR2x2_ASAP7_75t_L g17724 ( 
.A(n_17426),
.B(n_9173),
.Y(n_17724)
);

OAI31xp33_ASAP7_75t_L g17725 ( 
.A1(n_17182),
.A2(n_9525),
.A3(n_9132),
.B(n_9210),
.Y(n_17725)
);

AND2x2_ASAP7_75t_L g17726 ( 
.A(n_17181),
.B(n_10864),
.Y(n_17726)
);

AND2x2_ASAP7_75t_L g17727 ( 
.A(n_17175),
.B(n_17185),
.Y(n_17727)
);

OAI22xp5_ASAP7_75t_L g17728 ( 
.A1(n_17163),
.A2(n_10879),
.B1(n_10926),
.B2(n_10864),
.Y(n_17728)
);

INVx1_ASAP7_75t_L g17729 ( 
.A(n_17120),
.Y(n_17729)
);

INVx2_ASAP7_75t_SL g17730 ( 
.A(n_17249),
.Y(n_17730)
);

HB1xp67_ASAP7_75t_L g17731 ( 
.A(n_17208),
.Y(n_17731)
);

AOI22xp5_ASAP7_75t_L g17732 ( 
.A1(n_17191),
.A2(n_10926),
.B1(n_10932),
.B2(n_10879),
.Y(n_17732)
);

OAI22xp33_ASAP7_75t_L g17733 ( 
.A1(n_17401),
.A2(n_10926),
.B1(n_10932),
.B2(n_10879),
.Y(n_17733)
);

NAND2xp5_ASAP7_75t_L g17734 ( 
.A(n_17183),
.B(n_10600),
.Y(n_17734)
);

OAI332xp33_ASAP7_75t_L g17735 ( 
.A1(n_17505),
.A2(n_17113),
.A3(n_17115),
.B1(n_17594),
.B2(n_17358),
.B3(n_17131),
.C1(n_17613),
.C2(n_17317),
.Y(n_17735)
);

INVx1_ASAP7_75t_L g17736 ( 
.A(n_17502),
.Y(n_17736)
);

INVxp67_ASAP7_75t_SL g17737 ( 
.A(n_17577),
.Y(n_17737)
);

INVx1_ASAP7_75t_L g17738 ( 
.A(n_17247),
.Y(n_17738)
);

INVx2_ASAP7_75t_L g17739 ( 
.A(n_17282),
.Y(n_17739)
);

NAND2xp5_ASAP7_75t_L g17740 ( 
.A(n_17172),
.B(n_10600),
.Y(n_17740)
);

INVxp67_ASAP7_75t_L g17741 ( 
.A(n_17135),
.Y(n_17741)
);

AO221x1_ASAP7_75t_L g17742 ( 
.A1(n_17254),
.A2(n_10914),
.B1(n_10926),
.B2(n_10932),
.C(n_10879),
.Y(n_17742)
);

HB1xp67_ASAP7_75t_L g17743 ( 
.A(n_17192),
.Y(n_17743)
);

AND2x2_ASAP7_75t_L g17744 ( 
.A(n_17150),
.B(n_10879),
.Y(n_17744)
);

INVx1_ASAP7_75t_L g17745 ( 
.A(n_17265),
.Y(n_17745)
);

AND2x2_ASAP7_75t_L g17746 ( 
.A(n_17174),
.B(n_10879),
.Y(n_17746)
);

NAND2x1_ASAP7_75t_L g17747 ( 
.A(n_17149),
.B(n_17206),
.Y(n_17747)
);

INVx1_ASAP7_75t_L g17748 ( 
.A(n_17193),
.Y(n_17748)
);

OAI22xp5_ASAP7_75t_L g17749 ( 
.A1(n_17128),
.A2(n_10932),
.B1(n_10936),
.B2(n_10926),
.Y(n_17749)
);

AOI22xp5_ASAP7_75t_L g17750 ( 
.A1(n_17198),
.A2(n_10932),
.B1(n_10936),
.B2(n_10926),
.Y(n_17750)
);

NOR2x1_ASAP7_75t_L g17751 ( 
.A(n_17245),
.B(n_10932),
.Y(n_17751)
);

INVx1_ASAP7_75t_L g17752 ( 
.A(n_17168),
.Y(n_17752)
);

OR2x2_ASAP7_75t_L g17753 ( 
.A(n_17408),
.B(n_9173),
.Y(n_17753)
);

OAI21xp33_ASAP7_75t_L g17754 ( 
.A1(n_17516),
.A2(n_9230),
.B(n_9186),
.Y(n_17754)
);

INVxp33_ASAP7_75t_L g17755 ( 
.A(n_17338),
.Y(n_17755)
);

INVx2_ASAP7_75t_SL g17756 ( 
.A(n_17121),
.Y(n_17756)
);

A2O1A1Ixp33_ASAP7_75t_L g17757 ( 
.A1(n_17223),
.A2(n_10803),
.B(n_10855),
.C(n_9655),
.Y(n_17757)
);

INVxp67_ASAP7_75t_L g17758 ( 
.A(n_17596),
.Y(n_17758)
);

INVx2_ASAP7_75t_L g17759 ( 
.A(n_17363),
.Y(n_17759)
);

AOI211xp5_ASAP7_75t_L g17760 ( 
.A1(n_17531),
.A2(n_10936),
.B(n_10997),
.C(n_10985),
.Y(n_17760)
);

OR2x2_ASAP7_75t_L g17761 ( 
.A(n_17412),
.B(n_9247),
.Y(n_17761)
);

OAI32xp33_ASAP7_75t_L g17762 ( 
.A1(n_17104),
.A2(n_8623),
.A3(n_8698),
.B1(n_8688),
.B2(n_8618),
.Y(n_17762)
);

INVxp67_ASAP7_75t_SL g17763 ( 
.A(n_17177),
.Y(n_17763)
);

AOI22xp5_ASAP7_75t_L g17764 ( 
.A1(n_17187),
.A2(n_10936),
.B1(n_10997),
.B2(n_10985),
.Y(n_17764)
);

INVx2_ASAP7_75t_L g17765 ( 
.A(n_17196),
.Y(n_17765)
);

AOI33xp33_ASAP7_75t_L g17766 ( 
.A1(n_17153),
.A2(n_7117),
.A3(n_7060),
.B1(n_7183),
.B2(n_7127),
.B3(n_7111),
.Y(n_17766)
);

INVx1_ASAP7_75t_L g17767 ( 
.A(n_17124),
.Y(n_17767)
);

INVx2_ASAP7_75t_SL g17768 ( 
.A(n_17101),
.Y(n_17768)
);

HB1xp67_ASAP7_75t_L g17769 ( 
.A(n_17162),
.Y(n_17769)
);

AOI32xp33_ASAP7_75t_L g17770 ( 
.A1(n_17244),
.A2(n_10803),
.A3(n_10855),
.B1(n_8252),
.B2(n_8250),
.Y(n_17770)
);

INVx1_ASAP7_75t_L g17771 ( 
.A(n_17428),
.Y(n_17771)
);

NAND2xp5_ASAP7_75t_L g17772 ( 
.A(n_17469),
.B(n_10601),
.Y(n_17772)
);

INVx1_ASAP7_75t_L g17773 ( 
.A(n_17462),
.Y(n_17773)
);

HB1xp67_ASAP7_75t_L g17774 ( 
.A(n_17332),
.Y(n_17774)
);

INVx1_ASAP7_75t_L g17775 ( 
.A(n_17468),
.Y(n_17775)
);

INVx1_ASAP7_75t_L g17776 ( 
.A(n_17326),
.Y(n_17776)
);

OAI22xp5_ASAP7_75t_L g17777 ( 
.A1(n_17112),
.A2(n_10985),
.B1(n_10997),
.B2(n_10936),
.Y(n_17777)
);

AOI32xp33_ASAP7_75t_L g17778 ( 
.A1(n_17513),
.A2(n_10803),
.A3(n_10855),
.B1(n_8252),
.B2(n_8250),
.Y(n_17778)
);

AND2x2_ASAP7_75t_L g17779 ( 
.A(n_17310),
.B(n_17312),
.Y(n_17779)
);

INVx1_ASAP7_75t_L g17780 ( 
.A(n_17186),
.Y(n_17780)
);

NAND2xp5_ASAP7_75t_L g17781 ( 
.A(n_17169),
.B(n_10601),
.Y(n_17781)
);

INVx1_ASAP7_75t_L g17782 ( 
.A(n_17353),
.Y(n_17782)
);

INVx1_ASAP7_75t_L g17783 ( 
.A(n_17344),
.Y(n_17783)
);

NOR2xp67_ASAP7_75t_L g17784 ( 
.A(n_17210),
.B(n_9247),
.Y(n_17784)
);

INVx1_ASAP7_75t_L g17785 ( 
.A(n_17179),
.Y(n_17785)
);

AND2x2_ASAP7_75t_L g17786 ( 
.A(n_17156),
.B(n_10936),
.Y(n_17786)
);

INVx2_ASAP7_75t_L g17787 ( 
.A(n_17634),
.Y(n_17787)
);

INVxp33_ASAP7_75t_L g17788 ( 
.A(n_17612),
.Y(n_17788)
);

NAND2xp5_ASAP7_75t_L g17789 ( 
.A(n_17173),
.B(n_10614),
.Y(n_17789)
);

NOR2xp67_ASAP7_75t_SL g17790 ( 
.A(n_17117),
.B(n_17180),
.Y(n_17790)
);

NAND2xp5_ASAP7_75t_L g17791 ( 
.A(n_17409),
.B(n_10614),
.Y(n_17791)
);

INVx2_ASAP7_75t_L g17792 ( 
.A(n_17570),
.Y(n_17792)
);

A2O1A1Ixp33_ASAP7_75t_L g17793 ( 
.A1(n_17161),
.A2(n_9655),
.B(n_10044),
.C(n_8274),
.Y(n_17793)
);

INVx1_ASAP7_75t_L g17794 ( 
.A(n_17142),
.Y(n_17794)
);

HB1xp67_ASAP7_75t_L g17795 ( 
.A(n_17305),
.Y(n_17795)
);

XNOR2xp5_ASAP7_75t_L g17796 ( 
.A(n_17589),
.B(n_17607),
.Y(n_17796)
);

INVx1_ASAP7_75t_L g17797 ( 
.A(n_17341),
.Y(n_17797)
);

INVx1_ASAP7_75t_L g17798 ( 
.A(n_17205),
.Y(n_17798)
);

INVx2_ASAP7_75t_L g17799 ( 
.A(n_17570),
.Y(n_17799)
);

HB1xp67_ASAP7_75t_L g17800 ( 
.A(n_17364),
.Y(n_17800)
);

INVx3_ASAP7_75t_L g17801 ( 
.A(n_17625),
.Y(n_17801)
);

INVx1_ASAP7_75t_L g17802 ( 
.A(n_17116),
.Y(n_17802)
);

AOI22xp5_ASAP7_75t_L g17803 ( 
.A1(n_17342),
.A2(n_10997),
.B1(n_10985),
.B2(n_10949),
.Y(n_17803)
);

OR2x2_ASAP7_75t_L g17804 ( 
.A(n_17373),
.B(n_9296),
.Y(n_17804)
);

AND2x2_ASAP7_75t_L g17805 ( 
.A(n_17448),
.B(n_10985),
.Y(n_17805)
);

NAND2xp5_ASAP7_75t_L g17806 ( 
.A(n_17393),
.B(n_10635),
.Y(n_17806)
);

NAND4xp75_ASAP7_75t_SL g17807 ( 
.A(n_17437),
.B(n_8967),
.C(n_8179),
.D(n_10929),
.Y(n_17807)
);

OR2x2_ASAP7_75t_L g17808 ( 
.A(n_17390),
.B(n_9296),
.Y(n_17808)
);

OR2x2_ASAP7_75t_L g17809 ( 
.A(n_17392),
.B(n_9300),
.Y(n_17809)
);

AND2x2_ASAP7_75t_L g17810 ( 
.A(n_17355),
.B(n_10985),
.Y(n_17810)
);

NAND2xp5_ASAP7_75t_L g17811 ( 
.A(n_17232),
.B(n_10635),
.Y(n_17811)
);

NAND2x1_ASAP7_75t_SL g17812 ( 
.A(n_17362),
.B(n_9300),
.Y(n_17812)
);

NAND2xp5_ASAP7_75t_L g17813 ( 
.A(n_17237),
.B(n_10644),
.Y(n_17813)
);

OAI22xp5_ASAP7_75t_L g17814 ( 
.A1(n_17337),
.A2(n_10997),
.B1(n_10648),
.B2(n_10649),
.Y(n_17814)
);

INVx1_ASAP7_75t_L g17815 ( 
.A(n_17442),
.Y(n_17815)
);

NAND4xp75_ASAP7_75t_L g17816 ( 
.A(n_17446),
.B(n_9489),
.C(n_9194),
.D(n_9215),
.Y(n_17816)
);

BUFx2_ASAP7_75t_L g17817 ( 
.A(n_17410),
.Y(n_17817)
);

INVx1_ASAP7_75t_L g17818 ( 
.A(n_17300),
.Y(n_17818)
);

NAND2xp5_ASAP7_75t_L g17819 ( 
.A(n_17276),
.B(n_10644),
.Y(n_17819)
);

AO221x1_ASAP7_75t_L g17820 ( 
.A1(n_17288),
.A2(n_10997),
.B1(n_8623),
.B2(n_8698),
.C(n_8688),
.Y(n_17820)
);

HB1xp67_ASAP7_75t_L g17821 ( 
.A(n_17422),
.Y(n_17821)
);

OAI33xp33_ASAP7_75t_L g17822 ( 
.A1(n_17321),
.A2(n_10656),
.A3(n_10648),
.B1(n_10660),
.B2(n_10657),
.B3(n_10649),
.Y(n_17822)
);

NAND2xp5_ASAP7_75t_L g17823 ( 
.A(n_17461),
.B(n_10656),
.Y(n_17823)
);

NAND2xp5_ASAP7_75t_L g17824 ( 
.A(n_17384),
.B(n_10657),
.Y(n_17824)
);

AOI22xp33_ASAP7_75t_L g17825 ( 
.A1(n_17433),
.A2(n_8498),
.B1(n_8767),
.B2(n_8675),
.Y(n_17825)
);

AND2x2_ASAP7_75t_L g17826 ( 
.A(n_17357),
.B(n_8573),
.Y(n_17826)
);

NOR3xp33_ASAP7_75t_L g17827 ( 
.A(n_17146),
.B(n_9273),
.C(n_9041),
.Y(n_17827)
);

INVx1_ASAP7_75t_L g17828 ( 
.A(n_17615),
.Y(n_17828)
);

HB1xp67_ASAP7_75t_L g17829 ( 
.A(n_17430),
.Y(n_17829)
);

INVx1_ASAP7_75t_L g17830 ( 
.A(n_17375),
.Y(n_17830)
);

NAND2xp5_ASAP7_75t_SL g17831 ( 
.A(n_17460),
.B(n_8955),
.Y(n_17831)
);

AOI32xp33_ASAP7_75t_L g17832 ( 
.A1(n_17487),
.A2(n_8252),
.A3(n_8250),
.B1(n_10044),
.B2(n_9639),
.Y(n_17832)
);

NAND2xp5_ASAP7_75t_L g17833 ( 
.A(n_17413),
.B(n_10660),
.Y(n_17833)
);

NAND2xp5_ASAP7_75t_L g17834 ( 
.A(n_17417),
.B(n_10667),
.Y(n_17834)
);

OAI32xp33_ASAP7_75t_L g17835 ( 
.A1(n_17365),
.A2(n_17246),
.A3(n_17280),
.B1(n_17270),
.B2(n_17269),
.Y(n_17835)
);

OR2x2_ASAP7_75t_L g17836 ( 
.A(n_17618),
.B(n_9317),
.Y(n_17836)
);

AND2x2_ASAP7_75t_L g17837 ( 
.A(n_17619),
.B(n_17444),
.Y(n_17837)
);

AND2x2_ASAP7_75t_L g17838 ( 
.A(n_17558),
.B(n_17416),
.Y(n_17838)
);

NOR2xp33_ASAP7_75t_L g17839 ( 
.A(n_17303),
.B(n_17523),
.Y(n_17839)
);

AND2x2_ASAP7_75t_L g17840 ( 
.A(n_17406),
.B(n_8573),
.Y(n_17840)
);

NAND2xp5_ASAP7_75t_L g17841 ( 
.A(n_17376),
.B(n_10667),
.Y(n_17841)
);

NAND2xp5_ASAP7_75t_L g17842 ( 
.A(n_17470),
.B(n_10673),
.Y(n_17842)
);

INVx1_ASAP7_75t_L g17843 ( 
.A(n_17360),
.Y(n_17843)
);

AND2x4_ASAP7_75t_L g17844 ( 
.A(n_17438),
.B(n_17359),
.Y(n_17844)
);

AOI32xp33_ASAP7_75t_L g17845 ( 
.A1(n_17483),
.A2(n_10044),
.A3(n_9639),
.B1(n_9630),
.B2(n_10115),
.Y(n_17845)
);

INVx1_ASAP7_75t_L g17846 ( 
.A(n_17319),
.Y(n_17846)
);

OR2x2_ASAP7_75t_L g17847 ( 
.A(n_17351),
.B(n_9317),
.Y(n_17847)
);

INVx1_ASAP7_75t_L g17848 ( 
.A(n_17231),
.Y(n_17848)
);

OR2x2_ASAP7_75t_L g17849 ( 
.A(n_17370),
.B(n_9364),
.Y(n_17849)
);

OAI21xp5_ASAP7_75t_L g17850 ( 
.A1(n_17394),
.A2(n_9639),
.B(n_9630),
.Y(n_17850)
);

NAND4xp75_ASAP7_75t_L g17851 ( 
.A(n_17140),
.B(n_9284),
.C(n_9327),
.D(n_9570),
.Y(n_17851)
);

OR2x2_ASAP7_75t_L g17852 ( 
.A(n_17395),
.B(n_9364),
.Y(n_17852)
);

AND2x2_ASAP7_75t_L g17853 ( 
.A(n_17449),
.B(n_8573),
.Y(n_17853)
);

INVxp67_ASAP7_75t_SL g17854 ( 
.A(n_17522),
.Y(n_17854)
);

AOI22xp5_ASAP7_75t_L g17855 ( 
.A1(n_17330),
.A2(n_10949),
.B1(n_10929),
.B2(n_10610),
.Y(n_17855)
);

NOR2x1p5_ASAP7_75t_SL g17856 ( 
.A(n_17160),
.B(n_10673),
.Y(n_17856)
);

INVx1_ASAP7_75t_SL g17857 ( 
.A(n_17241),
.Y(n_17857)
);

AND2x2_ASAP7_75t_L g17858 ( 
.A(n_17451),
.B(n_8581),
.Y(n_17858)
);

NAND2xp5_ASAP7_75t_L g17859 ( 
.A(n_17471),
.B(n_10676),
.Y(n_17859)
);

OAI322xp33_ASAP7_75t_L g17860 ( 
.A1(n_17325),
.A2(n_8623),
.A3(n_8698),
.B1(n_8688),
.B2(n_8868),
.C1(n_8819),
.C2(n_8618),
.Y(n_17860)
);

OR2x2_ASAP7_75t_L g17861 ( 
.A(n_17415),
.B(n_9393),
.Y(n_17861)
);

AOI22xp5_ASAP7_75t_L g17862 ( 
.A1(n_17255),
.A2(n_10949),
.B1(n_10929),
.B2(n_10610),
.Y(n_17862)
);

INVxp67_ASAP7_75t_L g17863 ( 
.A(n_17480),
.Y(n_17863)
);

INVx1_ASAP7_75t_L g17864 ( 
.A(n_17152),
.Y(n_17864)
);

INVx1_ASAP7_75t_L g17865 ( 
.A(n_17530),
.Y(n_17865)
);

AOI22xp33_ASAP7_75t_L g17866 ( 
.A1(n_17361),
.A2(n_8498),
.B1(n_8835),
.B2(n_8767),
.Y(n_17866)
);

INVx2_ASAP7_75t_L g17867 ( 
.A(n_17500),
.Y(n_17867)
);

NOR2x1p5_ASAP7_75t_SL g17868 ( 
.A(n_17251),
.B(n_10676),
.Y(n_17868)
);

AOI211xp5_ASAP7_75t_L g17869 ( 
.A1(n_17281),
.A2(n_9426),
.B(n_8767),
.C(n_8837),
.Y(n_17869)
);

INVx1_ASAP7_75t_L g17870 ( 
.A(n_17532),
.Y(n_17870)
);

AOI22xp5_ASAP7_75t_L g17871 ( 
.A1(n_17267),
.A2(n_10949),
.B1(n_10929),
.B2(n_10610),
.Y(n_17871)
);

INVx2_ASAP7_75t_L g17872 ( 
.A(n_17389),
.Y(n_17872)
);

INVx1_ASAP7_75t_L g17873 ( 
.A(n_17534),
.Y(n_17873)
);

OR2x2_ASAP7_75t_L g17874 ( 
.A(n_17538),
.B(n_9393),
.Y(n_17874)
);

INVxp67_ASAP7_75t_SL g17875 ( 
.A(n_17543),
.Y(n_17875)
);

OAI31xp33_ASAP7_75t_L g17876 ( 
.A1(n_17339),
.A2(n_9525),
.A3(n_9132),
.B(n_9210),
.Y(n_17876)
);

INVx1_ASAP7_75t_L g17877 ( 
.A(n_17547),
.Y(n_17877)
);

AND2x2_ASAP7_75t_L g17878 ( 
.A(n_17453),
.B(n_8581),
.Y(n_17878)
);

INVx1_ASAP7_75t_L g17879 ( 
.A(n_17548),
.Y(n_17879)
);

AOI211xp5_ASAP7_75t_L g17880 ( 
.A1(n_17371),
.A2(n_9426),
.B(n_8835),
.C(n_8943),
.Y(n_17880)
);

INVx1_ASAP7_75t_L g17881 ( 
.A(n_17556),
.Y(n_17881)
);

AND2x2_ASAP7_75t_L g17882 ( 
.A(n_17458),
.B(n_8581),
.Y(n_17882)
);

NAND2xp5_ASAP7_75t_L g17883 ( 
.A(n_17425),
.B(n_10684),
.Y(n_17883)
);

INVx1_ASAP7_75t_L g17884 ( 
.A(n_17563),
.Y(n_17884)
);

NOR2xp33_ASAP7_75t_L g17885 ( 
.A(n_17525),
.B(n_10684),
.Y(n_17885)
);

AND2x2_ASAP7_75t_L g17886 ( 
.A(n_17464),
.B(n_8581),
.Y(n_17886)
);

HB1xp67_ASAP7_75t_L g17887 ( 
.A(n_17218),
.Y(n_17887)
);

AND2x2_ASAP7_75t_L g17888 ( 
.A(n_17467),
.B(n_8581),
.Y(n_17888)
);

INVx2_ASAP7_75t_SL g17889 ( 
.A(n_17275),
.Y(n_17889)
);

AOI21x1_ASAP7_75t_L g17890 ( 
.A1(n_17374),
.A2(n_9522),
.B(n_9462),
.Y(n_17890)
);

INVx1_ASAP7_75t_L g17891 ( 
.A(n_17225),
.Y(n_17891)
);

AOI32xp33_ASAP7_75t_L g17892 ( 
.A1(n_17309),
.A2(n_9630),
.A3(n_10115),
.B1(n_10103),
.B2(n_8509),
.Y(n_17892)
);

INVx1_ASAP7_75t_SL g17893 ( 
.A(n_17199),
.Y(n_17893)
);

A2O1A1Ixp33_ASAP7_75t_L g17894 ( 
.A1(n_17447),
.A2(n_8270),
.B(n_8274),
.C(n_10115),
.Y(n_17894)
);

INVx2_ASAP7_75t_L g17895 ( 
.A(n_17403),
.Y(n_17895)
);

INVx2_ASAP7_75t_L g17896 ( 
.A(n_17350),
.Y(n_17896)
);

INVx2_ASAP7_75t_SL g17897 ( 
.A(n_17271),
.Y(n_17897)
);

INVxp67_ASAP7_75t_L g17898 ( 
.A(n_17224),
.Y(n_17898)
);

NOR2xp33_ASAP7_75t_L g17899 ( 
.A(n_17307),
.B(n_10686),
.Y(n_17899)
);

AOI22xp33_ASAP7_75t_L g17900 ( 
.A1(n_17586),
.A2(n_17324),
.B1(n_17292),
.B2(n_17291),
.Y(n_17900)
);

OAI22xp5_ASAP7_75t_L g17901 ( 
.A1(n_17234),
.A2(n_10687),
.B1(n_10688),
.B2(n_10686),
.Y(n_17901)
);

HB1xp67_ASAP7_75t_L g17902 ( 
.A(n_17279),
.Y(n_17902)
);

AND2x2_ASAP7_75t_L g17903 ( 
.A(n_17472),
.B(n_17493),
.Y(n_17903)
);

INVxp67_ASAP7_75t_L g17904 ( 
.A(n_17228),
.Y(n_17904)
);

INVx2_ASAP7_75t_L g17905 ( 
.A(n_17354),
.Y(n_17905)
);

INVxp33_ASAP7_75t_L g17906 ( 
.A(n_17432),
.Y(n_17906)
);

NOR2xp67_ASAP7_75t_SL g17907 ( 
.A(n_17421),
.B(n_9090),
.Y(n_17907)
);

BUFx2_ASAP7_75t_L g17908 ( 
.A(n_17263),
.Y(n_17908)
);

NOR2xp33_ASAP7_75t_L g17909 ( 
.A(n_17334),
.B(n_10687),
.Y(n_17909)
);

INVx1_ASAP7_75t_L g17910 ( 
.A(n_17508),
.Y(n_17910)
);

INVx2_ASAP7_75t_L g17911 ( 
.A(n_17377),
.Y(n_17911)
);

INVx1_ASAP7_75t_L g17912 ( 
.A(n_17434),
.Y(n_17912)
);

NAND4xp75_ASAP7_75t_L g17913 ( 
.A(n_17236),
.B(n_17450),
.C(n_17195),
.D(n_17367),
.Y(n_17913)
);

INVx1_ASAP7_75t_L g17914 ( 
.A(n_17329),
.Y(n_17914)
);

INVx1_ASAP7_75t_L g17915 ( 
.A(n_17336),
.Y(n_17915)
);

XNOR2xp5_ASAP7_75t_L g17916 ( 
.A(n_17286),
.B(n_17302),
.Y(n_17916)
);

NAND4xp25_ASAP7_75t_L g17917 ( 
.A(n_17383),
.B(n_9230),
.C(n_9298),
.D(n_9186),
.Y(n_17917)
);

OAI33xp33_ASAP7_75t_L g17918 ( 
.A1(n_17295),
.A2(n_10701),
.A3(n_10688),
.B1(n_10719),
.B2(n_10712),
.B3(n_10692),
.Y(n_17918)
);

INVx1_ASAP7_75t_L g17919 ( 
.A(n_17621),
.Y(n_17919)
);

AND2x4_ASAP7_75t_L g17920 ( 
.A(n_17638),
.B(n_17495),
.Y(n_17920)
);

AND2x2_ASAP7_75t_L g17921 ( 
.A(n_17501),
.B(n_8581),
.Y(n_17921)
);

INVx2_ASAP7_75t_L g17922 ( 
.A(n_17476),
.Y(n_17922)
);

OAI22xp33_ASAP7_75t_L g17923 ( 
.A1(n_17323),
.A2(n_8837),
.B1(n_8943),
.B2(n_8835),
.Y(n_17923)
);

NOR2xp33_ASAP7_75t_L g17924 ( 
.A(n_17293),
.B(n_17463),
.Y(n_17924)
);

INVx1_ASAP7_75t_L g17925 ( 
.A(n_17294),
.Y(n_17925)
);

NAND2xp5_ASAP7_75t_L g17926 ( 
.A(n_17504),
.B(n_10692),
.Y(n_17926)
);

INVx3_ASAP7_75t_L g17927 ( 
.A(n_17202),
.Y(n_17927)
);

OR2x2_ASAP7_75t_L g17928 ( 
.A(n_17320),
.B(n_9462),
.Y(n_17928)
);

OAI32xp33_ASAP7_75t_L g17929 ( 
.A1(n_17238),
.A2(n_8623),
.A3(n_8698),
.B1(n_8688),
.B2(n_8618),
.Y(n_17929)
);

INVx1_ASAP7_75t_L g17930 ( 
.A(n_17261),
.Y(n_17930)
);

INVxp67_ASAP7_75t_SL g17931 ( 
.A(n_17620),
.Y(n_17931)
);

OR2x2_ASAP7_75t_L g17932 ( 
.A(n_17629),
.B(n_9522),
.Y(n_17932)
);

AOI22xp5_ASAP7_75t_L g17933 ( 
.A1(n_17327),
.A2(n_10610),
.B1(n_10814),
.B2(n_10591),
.Y(n_17933)
);

AO221x1_ASAP7_75t_L g17934 ( 
.A1(n_17509),
.A2(n_8688),
.B1(n_8698),
.B2(n_8623),
.C(n_8618),
.Y(n_17934)
);

INVx1_ASAP7_75t_L g17935 ( 
.A(n_17306),
.Y(n_17935)
);

INVx2_ASAP7_75t_L g17936 ( 
.A(n_17477),
.Y(n_17936)
);

INVx1_ASAP7_75t_L g17937 ( 
.A(n_17257),
.Y(n_17937)
);

NOR2xp33_ASAP7_75t_L g17938 ( 
.A(n_17466),
.B(n_10701),
.Y(n_17938)
);

INVx1_ASAP7_75t_L g17939 ( 
.A(n_17284),
.Y(n_17939)
);

NAND2xp5_ASAP7_75t_L g17940 ( 
.A(n_17541),
.B(n_10712),
.Y(n_17940)
);

NAND2xp5_ASAP7_75t_L g17941 ( 
.A(n_17496),
.B(n_10719),
.Y(n_17941)
);

O2A1O1Ixp33_ASAP7_75t_SL g17942 ( 
.A1(n_17399),
.A2(n_9555),
.B(n_10736),
.C(n_10734),
.Y(n_17942)
);

OAI32xp33_ASAP7_75t_L g17943 ( 
.A1(n_17221),
.A2(n_8819),
.A3(n_8870),
.B1(n_8868),
.B2(n_8618),
.Y(n_17943)
);

OR2x2_ASAP7_75t_L g17944 ( 
.A(n_17429),
.B(n_9555),
.Y(n_17944)
);

AND2x2_ASAP7_75t_L g17945 ( 
.A(n_17289),
.B(n_8695),
.Y(n_17945)
);

INVx1_ASAP7_75t_L g17946 ( 
.A(n_17201),
.Y(n_17946)
);

AOI22xp5_ASAP7_75t_L g17947 ( 
.A1(n_17521),
.A2(n_10814),
.B1(n_10959),
.B2(n_10591),
.Y(n_17947)
);

NAND2xp5_ASAP7_75t_L g17948 ( 
.A(n_17333),
.B(n_10734),
.Y(n_17948)
);

NOR2xp33_ASAP7_75t_L g17949 ( 
.A(n_17518),
.B(n_10736),
.Y(n_17949)
);

INVx1_ASAP7_75t_L g17950 ( 
.A(n_17256),
.Y(n_17950)
);

OR2x2_ASAP7_75t_L g17951 ( 
.A(n_17510),
.B(n_10741),
.Y(n_17951)
);

AOI22xp5_ASAP7_75t_L g17952 ( 
.A1(n_17524),
.A2(n_10814),
.B1(n_10959),
.B2(n_10591),
.Y(n_17952)
);

INVx1_ASAP7_75t_L g17953 ( 
.A(n_17203),
.Y(n_17953)
);

INVx2_ASAP7_75t_L g17954 ( 
.A(n_17478),
.Y(n_17954)
);

OR2x2_ASAP7_75t_L g17955 ( 
.A(n_17546),
.B(n_17553),
.Y(n_17955)
);

AND2x2_ASAP7_75t_SL g17956 ( 
.A(n_17217),
.B(n_10814),
.Y(n_17956)
);

NAND2xp5_ASAP7_75t_L g17957 ( 
.A(n_17335),
.B(n_10741),
.Y(n_17957)
);

NAND2xp5_ASAP7_75t_L g17958 ( 
.A(n_17343),
.B(n_10762),
.Y(n_17958)
);

INVx2_ASAP7_75t_L g17959 ( 
.A(n_17479),
.Y(n_17959)
);

INVx1_ASAP7_75t_L g17960 ( 
.A(n_17209),
.Y(n_17960)
);

INVx3_ASAP7_75t_L g17961 ( 
.A(n_17277),
.Y(n_17961)
);

INVx2_ASAP7_75t_L g17962 ( 
.A(n_17482),
.Y(n_17962)
);

AO221x1_ASAP7_75t_L g17963 ( 
.A1(n_17298),
.A2(n_8870),
.B1(n_8983),
.B2(n_8868),
.C(n_8819),
.Y(n_17963)
);

NAND2x2_ASAP7_75t_L g17964 ( 
.A(n_17226),
.B(n_9298),
.Y(n_17964)
);

NAND2xp5_ASAP7_75t_L g17965 ( 
.A(n_17347),
.B(n_10762),
.Y(n_17965)
);

OAI22xp33_ASAP7_75t_L g17966 ( 
.A1(n_17568),
.A2(n_8837),
.B1(n_8943),
.B2(n_8835),
.Y(n_17966)
);

INVx1_ASAP7_75t_SL g17967 ( 
.A(n_17402),
.Y(n_17967)
);

OAI32xp33_ASAP7_75t_L g17968 ( 
.A1(n_17340),
.A2(n_8868),
.A3(n_8983),
.B1(n_8870),
.B2(n_8819),
.Y(n_17968)
);

NAND4xp75_ASAP7_75t_L g17969 ( 
.A(n_17566),
.B(n_9570),
.C(n_9355),
.D(n_9405),
.Y(n_17969)
);

NOR2x1p5_ASAP7_75t_SL g17970 ( 
.A(n_17287),
.B(n_10766),
.Y(n_17970)
);

INVx1_ASAP7_75t_L g17971 ( 
.A(n_17227),
.Y(n_17971)
);

OAI322xp33_ASAP7_75t_L g17972 ( 
.A1(n_17637),
.A2(n_8868),
.A3(n_8819),
.B1(n_8999),
.B2(n_9009),
.C1(n_8983),
.C2(n_8870),
.Y(n_17972)
);

NAND4xp75_ASAP7_75t_SL g17973 ( 
.A(n_17455),
.B(n_8967),
.C(n_8179),
.D(n_8105),
.Y(n_17973)
);

NAND2xp5_ASAP7_75t_L g17974 ( 
.A(n_17296),
.B(n_10766),
.Y(n_17974)
);

OAI21xp5_ASAP7_75t_L g17975 ( 
.A1(n_17290),
.A2(n_10103),
.B(n_9851),
.Y(n_17975)
);

NOR2xp33_ASAP7_75t_L g17976 ( 
.A(n_17529),
.B(n_10767),
.Y(n_17976)
);

O2A1O1Ixp33_ASAP7_75t_L g17977 ( 
.A1(n_17616),
.A2(n_8870),
.B(n_8999),
.C(n_8983),
.Y(n_17977)
);

OAI32xp33_ASAP7_75t_L g17978 ( 
.A1(n_17346),
.A2(n_9009),
.A3(n_9011),
.B1(n_8999),
.B2(n_8983),
.Y(n_17978)
);

INVxp33_ASAP7_75t_L g17979 ( 
.A(n_17441),
.Y(n_17979)
);

NAND2xp5_ASAP7_75t_L g17980 ( 
.A(n_17297),
.B(n_10767),
.Y(n_17980)
);

INVx2_ASAP7_75t_L g17981 ( 
.A(n_17486),
.Y(n_17981)
);

AND2x2_ASAP7_75t_L g17982 ( 
.A(n_17308),
.B(n_8695),
.Y(n_17982)
);

AOI32xp33_ASAP7_75t_L g17983 ( 
.A1(n_17239),
.A2(n_10103),
.A3(n_8509),
.B1(n_8523),
.B2(n_8519),
.Y(n_17983)
);

INVx1_ASAP7_75t_L g17984 ( 
.A(n_17443),
.Y(n_17984)
);

NAND2xp5_ASAP7_75t_L g17985 ( 
.A(n_17211),
.B(n_10779),
.Y(n_17985)
);

NAND2xp5_ASAP7_75t_L g17986 ( 
.A(n_17213),
.B(n_10779),
.Y(n_17986)
);

OAI22xp33_ASAP7_75t_L g17987 ( 
.A1(n_17243),
.A2(n_8835),
.B1(n_8943),
.B2(n_8837),
.Y(n_17987)
);

INVx1_ASAP7_75t_L g17988 ( 
.A(n_17452),
.Y(n_17988)
);

INVx1_ASAP7_75t_L g17989 ( 
.A(n_17457),
.Y(n_17989)
);

INVx1_ASAP7_75t_L g17990 ( 
.A(n_17459),
.Y(n_17990)
);

NOR3xp33_ASAP7_75t_L g17991 ( 
.A(n_17602),
.B(n_9041),
.C(n_8964),
.Y(n_17991)
);

AND2x2_ASAP7_75t_L g17992 ( 
.A(n_17536),
.B(n_8695),
.Y(n_17992)
);

OAI322xp33_ASAP7_75t_L g17993 ( 
.A1(n_17587),
.A2(n_9065),
.A3(n_9009),
.B1(n_9207),
.B2(n_9214),
.C1(n_9011),
.C2(n_8999),
.Y(n_17993)
);

AND2x2_ASAP7_75t_L g17994 ( 
.A(n_17314),
.B(n_8695),
.Y(n_17994)
);

INVxp67_ASAP7_75t_L g17995 ( 
.A(n_17475),
.Y(n_17995)
);

INVx1_ASAP7_75t_L g17996 ( 
.A(n_17248),
.Y(n_17996)
);

AND2x2_ASAP7_75t_L g17997 ( 
.A(n_17366),
.B(n_8695),
.Y(n_17997)
);

INVx1_ASAP7_75t_L g17998 ( 
.A(n_17252),
.Y(n_17998)
);

HB1xp67_ASAP7_75t_L g17999 ( 
.A(n_17494),
.Y(n_17999)
);

OAI32xp33_ASAP7_75t_L g18000 ( 
.A1(n_17266),
.A2(n_8999),
.A3(n_9065),
.B1(n_9011),
.B2(n_9009),
.Y(n_18000)
);

NAND2xp5_ASAP7_75t_L g18001 ( 
.A(n_17581),
.B(n_17592),
.Y(n_18001)
);

NAND2xp5_ASAP7_75t_L g18002 ( 
.A(n_17593),
.B(n_10785),
.Y(n_18002)
);

INVx2_ASAP7_75t_SL g18003 ( 
.A(n_17396),
.Y(n_18003)
);

OR3x2_ASAP7_75t_L g18004 ( 
.A(n_17628),
.B(n_8179),
.C(n_8967),
.Y(n_18004)
);

AND2x2_ASAP7_75t_L g18005 ( 
.A(n_17622),
.B(n_8695),
.Y(n_18005)
);

INVx2_ASAP7_75t_SL g18006 ( 
.A(n_17385),
.Y(n_18006)
);

AOI22xp33_ASAP7_75t_L g18007 ( 
.A1(n_17571),
.A2(n_8837),
.B1(n_8943),
.B2(n_8835),
.Y(n_18007)
);

INVx1_ASAP7_75t_L g18008 ( 
.A(n_17520),
.Y(n_18008)
);

AND2x2_ASAP7_75t_L g18009 ( 
.A(n_17603),
.B(n_8742),
.Y(n_18009)
);

INVx2_ASAP7_75t_L g18010 ( 
.A(n_17489),
.Y(n_18010)
);

INVx2_ASAP7_75t_L g18011 ( 
.A(n_17490),
.Y(n_18011)
);

INVx1_ASAP7_75t_L g18012 ( 
.A(n_17573),
.Y(n_18012)
);

INVx1_ASAP7_75t_L g18013 ( 
.A(n_17431),
.Y(n_18013)
);

INVx1_ASAP7_75t_L g18014 ( 
.A(n_17277),
.Y(n_18014)
);

O2A1O1Ixp5_ASAP7_75t_R g18015 ( 
.A1(n_17274),
.A2(n_9564),
.B(n_9574),
.C(n_9467),
.Y(n_18015)
);

INVx2_ASAP7_75t_L g18016 ( 
.A(n_17316),
.Y(n_18016)
);

NOR2xp33_ASAP7_75t_L g18017 ( 
.A(n_17230),
.B(n_17588),
.Y(n_18017)
);

OAI22xp5_ASAP7_75t_SL g18018 ( 
.A1(n_17626),
.A2(n_9163),
.B1(n_9439),
.B2(n_8955),
.Y(n_18018)
);

OR2x2_ASAP7_75t_L g18019 ( 
.A(n_17555),
.B(n_10785),
.Y(n_18019)
);

INVx1_ASAP7_75t_L g18020 ( 
.A(n_17590),
.Y(n_18020)
);

OA222x2_ASAP7_75t_L g18021 ( 
.A1(n_17609),
.A2(n_9496),
.B1(n_9344),
.B2(n_9498),
.C1(n_9460),
.C2(n_9325),
.Y(n_18021)
);

INVx1_ASAP7_75t_L g18022 ( 
.A(n_17564),
.Y(n_18022)
);

NAND2xp5_ASAP7_75t_L g18023 ( 
.A(n_17597),
.B(n_10790),
.Y(n_18023)
);

AND2x4_ASAP7_75t_L g18024 ( 
.A(n_17511),
.B(n_9325),
.Y(n_18024)
);

INVx2_ASAP7_75t_L g18025 ( 
.A(n_17348),
.Y(n_18025)
);

AND2x2_ASAP7_75t_L g18026 ( 
.A(n_17386),
.B(n_8742),
.Y(n_18026)
);

INVx1_ASAP7_75t_L g18027 ( 
.A(n_17585),
.Y(n_18027)
);

INVx2_ASAP7_75t_L g18028 ( 
.A(n_17605),
.Y(n_18028)
);

INVx1_ASAP7_75t_L g18029 ( 
.A(n_17611),
.Y(n_18029)
);

OAI322xp33_ASAP7_75t_L g18030 ( 
.A1(n_17527),
.A2(n_9207),
.A3(n_9011),
.B1(n_9214),
.B2(n_9223),
.C1(n_9065),
.C2(n_9009),
.Y(n_18030)
);

INVx1_ASAP7_75t_L g18031 ( 
.A(n_17551),
.Y(n_18031)
);

INVx1_ASAP7_75t_L g18032 ( 
.A(n_17639),
.Y(n_18032)
);

AND2x2_ASAP7_75t_L g18033 ( 
.A(n_17379),
.B(n_17610),
.Y(n_18033)
);

INVx1_ASAP7_75t_L g18034 ( 
.A(n_17633),
.Y(n_18034)
);

AND2x2_ASAP7_75t_L g18035 ( 
.A(n_17492),
.B(n_8742),
.Y(n_18035)
);

NAND2xp5_ASAP7_75t_L g18036 ( 
.A(n_17264),
.B(n_10790),
.Y(n_18036)
);

AND2x2_ASAP7_75t_L g18037 ( 
.A(n_17368),
.B(n_8742),
.Y(n_18037)
);

XNOR2x1_ASAP7_75t_L g18038 ( 
.A(n_17549),
.B(n_10789),
.Y(n_18038)
);

NAND5xp2_ASAP7_75t_L g18039 ( 
.A(n_17240),
.B(n_9527),
.C(n_9429),
.D(n_9411),
.E(n_9375),
.Y(n_18039)
);

OR2x2_ASAP7_75t_L g18040 ( 
.A(n_17514),
.B(n_10794),
.Y(n_18040)
);

INVx1_ASAP7_75t_L g18041 ( 
.A(n_17485),
.Y(n_18041)
);

AOI22xp33_ASAP7_75t_L g18042 ( 
.A1(n_17545),
.A2(n_8837),
.B1(n_8943),
.B2(n_8835),
.Y(n_18042)
);

OA222x2_ASAP7_75t_L g18043 ( 
.A1(n_17617),
.A2(n_17584),
.B1(n_17424),
.B2(n_17595),
.C1(n_17601),
.C2(n_17599),
.Y(n_18043)
);

AOI22xp33_ASAP7_75t_L g18044 ( 
.A1(n_17533),
.A2(n_8837),
.B1(n_8943),
.B2(n_8835),
.Y(n_18044)
);

INVx1_ASAP7_75t_L g18045 ( 
.A(n_17498),
.Y(n_18045)
);

OR2x2_ASAP7_75t_L g18046 ( 
.A(n_17515),
.B(n_10794),
.Y(n_18046)
);

INVx1_ASAP7_75t_L g18047 ( 
.A(n_17635),
.Y(n_18047)
);

INVx1_ASAP7_75t_L g18048 ( 
.A(n_17352),
.Y(n_18048)
);

AOI22xp5_ASAP7_75t_L g18049 ( 
.A1(n_17540),
.A2(n_10959),
.B1(n_9244),
.B2(n_9253),
.Y(n_18049)
);

AOI211xp5_ASAP7_75t_L g18050 ( 
.A1(n_17278),
.A2(n_8837),
.B(n_8951),
.C(n_8943),
.Y(n_18050)
);

OAI322xp33_ASAP7_75t_L g18051 ( 
.A1(n_17427),
.A2(n_9011),
.A3(n_9207),
.B1(n_9223),
.B2(n_9237),
.C1(n_9214),
.C2(n_9065),
.Y(n_18051)
);

INVx1_ASAP7_75t_L g18052 ( 
.A(n_17356),
.Y(n_18052)
);

NAND2xp5_ASAP7_75t_L g18053 ( 
.A(n_17512),
.B(n_10798),
.Y(n_18053)
);

AND2x4_ASAP7_75t_L g18054 ( 
.A(n_17559),
.B(n_9325),
.Y(n_18054)
);

OR2x2_ASAP7_75t_L g18055 ( 
.A(n_17569),
.B(n_10798),
.Y(n_18055)
);

AOI22xp5_ASAP7_75t_L g18056 ( 
.A1(n_17229),
.A2(n_10959),
.B1(n_9244),
.B2(n_9253),
.Y(n_18056)
);

INVx1_ASAP7_75t_L g18057 ( 
.A(n_17380),
.Y(n_18057)
);

INVx1_ASAP7_75t_L g18058 ( 
.A(n_17382),
.Y(n_18058)
);

O2A1O1Ixp5_ASAP7_75t_SL g18059 ( 
.A1(n_17423),
.A2(n_10804),
.B(n_10806),
.C(n_10802),
.Y(n_18059)
);

INVx1_ASAP7_75t_L g18060 ( 
.A(n_17387),
.Y(n_18060)
);

INVx1_ASAP7_75t_L g18061 ( 
.A(n_17400),
.Y(n_18061)
);

OAI31xp67_ASAP7_75t_L g18062 ( 
.A1(n_17272),
.A2(n_9377),
.A3(n_9851),
.B(n_9716),
.Y(n_18062)
);

OR2x2_ASAP7_75t_L g18063 ( 
.A(n_17576),
.B(n_10802),
.Y(n_18063)
);

INVx2_ASAP7_75t_L g18064 ( 
.A(n_17258),
.Y(n_18064)
);

INVx2_ASAP7_75t_L g18065 ( 
.A(n_17600),
.Y(n_18065)
);

OR2x2_ASAP7_75t_L g18066 ( 
.A(n_17414),
.B(n_10804),
.Y(n_18066)
);

AOI22xp5_ASAP7_75t_L g18067 ( 
.A1(n_17519),
.A2(n_9244),
.B1(n_9253),
.B2(n_9222),
.Y(n_18067)
);

INVx2_ASAP7_75t_L g18068 ( 
.A(n_17194),
.Y(n_18068)
);

INVx1_ASAP7_75t_L g18069 ( 
.A(n_17561),
.Y(n_18069)
);

OAI21xp33_ASAP7_75t_L g18070 ( 
.A1(n_17349),
.A2(n_9460),
.B(n_9344),
.Y(n_18070)
);

AOI211xp5_ASAP7_75t_L g18071 ( 
.A1(n_17283),
.A2(n_8951),
.B(n_9031),
.C(n_8969),
.Y(n_18071)
);

NAND2xp5_ASAP7_75t_L g18072 ( 
.A(n_17560),
.B(n_10806),
.Y(n_18072)
);

INVx2_ASAP7_75t_SL g18073 ( 
.A(n_17318),
.Y(n_18073)
);

NAND2x1p5_ASAP7_75t_L g18074 ( 
.A(n_17439),
.B(n_8955),
.Y(n_18074)
);

BUFx2_ASAP7_75t_L g18075 ( 
.A(n_17456),
.Y(n_18075)
);

INVx1_ASAP7_75t_L g18076 ( 
.A(n_17557),
.Y(n_18076)
);

NAND2xp5_ASAP7_75t_L g18077 ( 
.A(n_17484),
.B(n_10809),
.Y(n_18077)
);

AND2x2_ASAP7_75t_L g18078 ( 
.A(n_17445),
.B(n_8742),
.Y(n_18078)
);

AOI22xp5_ASAP7_75t_L g18079 ( 
.A1(n_17405),
.A2(n_17507),
.B1(n_17632),
.B2(n_17583),
.Y(n_18079)
);

NAND2xp33_ASAP7_75t_L g18080 ( 
.A(n_17465),
.B(n_8951),
.Y(n_18080)
);

INVx2_ASAP7_75t_SL g18081 ( 
.A(n_17488),
.Y(n_18081)
);

INVx2_ASAP7_75t_L g18082 ( 
.A(n_17440),
.Y(n_18082)
);

HB1xp67_ASAP7_75t_L g18083 ( 
.A(n_17645),
.Y(n_18083)
);

INVx1_ASAP7_75t_L g18084 ( 
.A(n_17795),
.Y(n_18084)
);

INVx2_ASAP7_75t_L g18085 ( 
.A(n_17727),
.Y(n_18085)
);

INVxp67_ASAP7_75t_L g18086 ( 
.A(n_17703),
.Y(n_18086)
);

INVxp67_ASAP7_75t_L g18087 ( 
.A(n_17769),
.Y(n_18087)
);

AOI21xp5_ASAP7_75t_L g18088 ( 
.A1(n_17721),
.A2(n_17604),
.B(n_17345),
.Y(n_18088)
);

OR2x2_ASAP7_75t_L g18089 ( 
.A(n_17722),
.B(n_17591),
.Y(n_18089)
);

NAND2xp5_ASAP7_75t_SL g18090 ( 
.A(n_17647),
.B(n_17632),
.Y(n_18090)
);

INVx3_ASAP7_75t_SL g18091 ( 
.A(n_17730),
.Y(n_18091)
);

NAND2xp5_ASAP7_75t_L g18092 ( 
.A(n_17796),
.B(n_17497),
.Y(n_18092)
);

INVx2_ASAP7_75t_L g18093 ( 
.A(n_17739),
.Y(n_18093)
);

NAND2xp5_ASAP7_75t_L g18094 ( 
.A(n_17756),
.B(n_17499),
.Y(n_18094)
);

AND2x2_ASAP7_75t_L g18095 ( 
.A(n_17684),
.B(n_17369),
.Y(n_18095)
);

AND2x2_ASAP7_75t_L g18096 ( 
.A(n_18043),
.B(n_17331),
.Y(n_18096)
);

NAND2xp33_ASAP7_75t_SL g18097 ( 
.A(n_17747),
.B(n_17623),
.Y(n_18097)
);

NAND2xp5_ASAP7_75t_SL g18098 ( 
.A(n_17666),
.B(n_17404),
.Y(n_18098)
);

AOI22xp33_ASAP7_75t_L g18099 ( 
.A1(n_17900),
.A2(n_17491),
.B1(n_17398),
.B2(n_17481),
.Y(n_18099)
);

NAND2xp5_ASAP7_75t_L g18100 ( 
.A(n_17737),
.B(n_17388),
.Y(n_18100)
);

AND2x2_ASAP7_75t_L g18101 ( 
.A(n_17837),
.B(n_17419),
.Y(n_18101)
);

OR2x6_ASAP7_75t_L g18102 ( 
.A(n_17671),
.B(n_17285),
.Y(n_18102)
);

NAND2x1_ASAP7_75t_L g18103 ( 
.A(n_17961),
.B(n_17565),
.Y(n_18103)
);

NOR2xp33_ASAP7_75t_L g18104 ( 
.A(n_17788),
.B(n_17526),
.Y(n_18104)
);

INVx4_ASAP7_75t_L g18105 ( 
.A(n_17801),
.Y(n_18105)
);

AOI21xp33_ASAP7_75t_L g18106 ( 
.A1(n_17755),
.A2(n_17268),
.B(n_17580),
.Y(n_18106)
);

AND2x2_ASAP7_75t_L g18107 ( 
.A(n_17817),
.B(n_17420),
.Y(n_18107)
);

HB1xp67_ASAP7_75t_L g18108 ( 
.A(n_17887),
.Y(n_18108)
);

NOR3xp33_ASAP7_75t_L g18109 ( 
.A(n_17735),
.B(n_17676),
.C(n_17854),
.Y(n_18109)
);

AND2x2_ASAP7_75t_L g18110 ( 
.A(n_17838),
.B(n_17436),
.Y(n_18110)
);

OAI31xp33_ASAP7_75t_L g18111 ( 
.A1(n_17715),
.A2(n_17608),
.A3(n_17567),
.B(n_17574),
.Y(n_18111)
);

NAND3xp33_ASAP7_75t_SL g18112 ( 
.A(n_17664),
.B(n_17506),
.C(n_17614),
.Y(n_18112)
);

AND2x2_ASAP7_75t_L g18113 ( 
.A(n_17689),
.B(n_17407),
.Y(n_18113)
);

NAND2xp33_ASAP7_75t_SL g18114 ( 
.A(n_17812),
.B(n_17624),
.Y(n_18114)
);

NAND2xp33_ASAP7_75t_L g18115 ( 
.A(n_17652),
.B(n_17631),
.Y(n_18115)
);

INVx1_ASAP7_75t_L g18116 ( 
.A(n_17774),
.Y(n_18116)
);

NAND2xp5_ASAP7_75t_L g18117 ( 
.A(n_17662),
.B(n_17967),
.Y(n_18117)
);

NAND2xp5_ASAP7_75t_L g18118 ( 
.A(n_17763),
.B(n_17572),
.Y(n_18118)
);

NOR4xp25_ASAP7_75t_SL g18119 ( 
.A(n_17678),
.B(n_17517),
.C(n_17579),
.D(n_17537),
.Y(n_18119)
);

BUFx3_ASAP7_75t_L g18120 ( 
.A(n_17920),
.Y(n_18120)
);

AOI21xp5_ASAP7_75t_L g18121 ( 
.A1(n_17875),
.A2(n_17578),
.B(n_17575),
.Y(n_18121)
);

INVx5_ASAP7_75t_L g18122 ( 
.A(n_17768),
.Y(n_18122)
);

NOR2xp33_ASAP7_75t_L g18123 ( 
.A(n_17893),
.B(n_17554),
.Y(n_18123)
);

INVx1_ASAP7_75t_L g18124 ( 
.A(n_17731),
.Y(n_18124)
);

OR2x2_ASAP7_75t_L g18125 ( 
.A(n_17649),
.B(n_17550),
.Y(n_18125)
);

OR2x2_ASAP7_75t_L g18126 ( 
.A(n_17759),
.B(n_17630),
.Y(n_18126)
);

AND2x2_ASAP7_75t_L g18127 ( 
.A(n_17800),
.B(n_17627),
.Y(n_18127)
);

INVx1_ASAP7_75t_L g18128 ( 
.A(n_17821),
.Y(n_18128)
);

NAND2xp5_ASAP7_75t_L g18129 ( 
.A(n_17711),
.B(n_17636),
.Y(n_18129)
);

AND2x2_ASAP7_75t_SL g18130 ( 
.A(n_17920),
.B(n_17552),
.Y(n_18130)
);

NOR3xp33_ASAP7_75t_L g18131 ( 
.A(n_17650),
.B(n_17328),
.C(n_17381),
.Y(n_18131)
);

AND2x4_ASAP7_75t_L g18132 ( 
.A(n_17644),
.B(n_9344),
.Y(n_18132)
);

AOI221xp5_ASAP7_75t_SL g18133 ( 
.A1(n_17741),
.A2(n_10812),
.B1(n_10813),
.B2(n_10810),
.C(n_10809),
.Y(n_18133)
);

INVx2_ASAP7_75t_L g18134 ( 
.A(n_17691),
.Y(n_18134)
);

OR2x2_ASAP7_75t_L g18135 ( 
.A(n_17745),
.B(n_10810),
.Y(n_18135)
);

HB1xp67_ASAP7_75t_L g18136 ( 
.A(n_17829),
.Y(n_18136)
);

INVx1_ASAP7_75t_L g18137 ( 
.A(n_17856),
.Y(n_18137)
);

NOR3xp33_ASAP7_75t_L g18138 ( 
.A(n_17686),
.B(n_10789),
.C(n_8509),
.Y(n_18138)
);

NAND2xp5_ASAP7_75t_L g18139 ( 
.A(n_17682),
.B(n_10812),
.Y(n_18139)
);

NAND2xp5_ASAP7_75t_L g18140 ( 
.A(n_17683),
.B(n_10813),
.Y(n_18140)
);

AND2x2_ASAP7_75t_L g18141 ( 
.A(n_17994),
.B(n_8742),
.Y(n_18141)
);

INVx1_ASAP7_75t_L g18142 ( 
.A(n_17743),
.Y(n_18142)
);

INVx1_ASAP7_75t_L g18143 ( 
.A(n_17688),
.Y(n_18143)
);

AND2x2_ASAP7_75t_L g18144 ( 
.A(n_17765),
.B(n_8783),
.Y(n_18144)
);

AOI22xp5_ASAP7_75t_L g18145 ( 
.A1(n_17857),
.A2(n_8969),
.B1(n_9031),
.B2(n_8951),
.Y(n_18145)
);

INVx1_ASAP7_75t_SL g18146 ( 
.A(n_17672),
.Y(n_18146)
);

INVx2_ASAP7_75t_SL g18147 ( 
.A(n_17644),
.Y(n_18147)
);

NOR2x1p5_ASAP7_75t_L g18148 ( 
.A(n_17931),
.B(n_9344),
.Y(n_18148)
);

AND2x2_ASAP7_75t_L g18149 ( 
.A(n_17661),
.B(n_8783),
.Y(n_18149)
);

AND2x2_ASAP7_75t_L g18150 ( 
.A(n_17681),
.B(n_8783),
.Y(n_18150)
);

NAND2xp5_ASAP7_75t_L g18151 ( 
.A(n_17785),
.B(n_17889),
.Y(n_18151)
);

OR2x2_ASAP7_75t_L g18152 ( 
.A(n_17702),
.B(n_10815),
.Y(n_18152)
);

NAND2xp5_ASAP7_75t_L g18153 ( 
.A(n_17802),
.B(n_10815),
.Y(n_18153)
);

NOR3xp33_ASAP7_75t_L g18154 ( 
.A(n_17712),
.B(n_9121),
.C(n_9065),
.Y(n_18154)
);

AND2x4_ASAP7_75t_L g18155 ( 
.A(n_17844),
.B(n_9460),
.Y(n_18155)
);

INVx2_ASAP7_75t_L g18156 ( 
.A(n_18074),
.Y(n_18156)
);

INVx1_ASAP7_75t_L g18157 ( 
.A(n_17902),
.Y(n_18157)
);

INVx1_ASAP7_75t_L g18158 ( 
.A(n_17868),
.Y(n_18158)
);

INVx2_ASAP7_75t_L g18159 ( 
.A(n_18038),
.Y(n_18159)
);

INVx1_ASAP7_75t_L g18160 ( 
.A(n_17970),
.Y(n_18160)
);

INVx2_ASAP7_75t_L g18161 ( 
.A(n_17786),
.Y(n_18161)
);

INVx1_ASAP7_75t_L g18162 ( 
.A(n_17780),
.Y(n_18162)
);

INVxp67_ASAP7_75t_L g18163 ( 
.A(n_17839),
.Y(n_18163)
);

BUFx2_ASAP7_75t_L g18164 ( 
.A(n_17646),
.Y(n_18164)
);

CKINVDCx5p33_ASAP7_75t_R g18165 ( 
.A(n_17916),
.Y(n_18165)
);

AND2x2_ASAP7_75t_SL g18166 ( 
.A(n_17844),
.B(n_8951),
.Y(n_18166)
);

INVx2_ASAP7_75t_L g18167 ( 
.A(n_17726),
.Y(n_18167)
);

AO21x1_ASAP7_75t_L g18168 ( 
.A1(n_17924),
.A2(n_18014),
.B(n_18017),
.Y(n_18168)
);

BUFx3_ASAP7_75t_L g18169 ( 
.A(n_17783),
.Y(n_18169)
);

INVx2_ASAP7_75t_L g18170 ( 
.A(n_17805),
.Y(n_18170)
);

HB1xp67_ASAP7_75t_L g18171 ( 
.A(n_17700),
.Y(n_18171)
);

INVx2_ASAP7_75t_L g18172 ( 
.A(n_17945),
.Y(n_18172)
);

NOR2xp33_ASAP7_75t_L g18173 ( 
.A(n_17719),
.B(n_10819),
.Y(n_18173)
);

AND2x2_ASAP7_75t_L g18174 ( 
.A(n_17692),
.B(n_8783),
.Y(n_18174)
);

NAND2xp33_ASAP7_75t_SL g18175 ( 
.A(n_17790),
.B(n_17680),
.Y(n_18175)
);

AND2x2_ASAP7_75t_L g18176 ( 
.A(n_17698),
.B(n_8783),
.Y(n_18176)
);

NAND2xp5_ASAP7_75t_L g18177 ( 
.A(n_17927),
.B(n_10819),
.Y(n_18177)
);

AND2x2_ASAP7_75t_L g18178 ( 
.A(n_17701),
.B(n_8783),
.Y(n_18178)
);

NOR2xp33_ASAP7_75t_L g18179 ( 
.A(n_17794),
.B(n_10823),
.Y(n_18179)
);

NAND3xp33_ASAP7_75t_L g18180 ( 
.A(n_17758),
.B(n_8969),
.C(n_8951),
.Y(n_18180)
);

NAND2xp5_ASAP7_75t_L g18181 ( 
.A(n_17704),
.B(n_17752),
.Y(n_18181)
);

OAI22xp5_ASAP7_75t_L g18182 ( 
.A1(n_17717),
.A2(n_10828),
.B1(n_10830),
.B2(n_10823),
.Y(n_18182)
);

AOI21xp5_ASAP7_75t_L g18183 ( 
.A1(n_17675),
.A2(n_17648),
.B(n_17835),
.Y(n_18183)
);

AND2x2_ASAP7_75t_L g18184 ( 
.A(n_17787),
.B(n_8884),
.Y(n_18184)
);

INVx2_ASAP7_75t_SL g18185 ( 
.A(n_17646),
.Y(n_18185)
);

INVxp67_ASAP7_75t_L g18186 ( 
.A(n_17653),
.Y(n_18186)
);

NOR2xp33_ASAP7_75t_L g18187 ( 
.A(n_17723),
.B(n_17736),
.Y(n_18187)
);

OAI221xp5_ASAP7_75t_L g18188 ( 
.A1(n_17641),
.A2(n_9223),
.B1(n_9237),
.B2(n_9214),
.C(n_9207),
.Y(n_18188)
);

AOI211xp5_ASAP7_75t_L g18189 ( 
.A1(n_17706),
.A2(n_17642),
.B(n_17659),
.C(n_17979),
.Y(n_18189)
);

OR2x2_ASAP7_75t_L g18190 ( 
.A(n_17798),
.B(n_10828),
.Y(n_18190)
);

OAI31xp33_ASAP7_75t_L g18191 ( 
.A1(n_17663),
.A2(n_9299),
.A3(n_9518),
.B(n_9281),
.Y(n_18191)
);

NAND2xp5_ASAP7_75t_L g18192 ( 
.A(n_17903),
.B(n_10830),
.Y(n_18192)
);

OR2x2_ASAP7_75t_L g18193 ( 
.A(n_17914),
.B(n_10833),
.Y(n_18193)
);

INVx1_ASAP7_75t_L g18194 ( 
.A(n_17915),
.Y(n_18194)
);

AND2x2_ASAP7_75t_L g18195 ( 
.A(n_17992),
.B(n_8884),
.Y(n_18195)
);

NAND2xp5_ASAP7_75t_L g18196 ( 
.A(n_17713),
.B(n_10833),
.Y(n_18196)
);

INVx1_ASAP7_75t_SL g18197 ( 
.A(n_17690),
.Y(n_18197)
);

AND2x2_ASAP7_75t_L g18198 ( 
.A(n_17846),
.B(n_8884),
.Y(n_18198)
);

INVx1_ASAP7_75t_L g18199 ( 
.A(n_17643),
.Y(n_18199)
);

AOI22xp5_ASAP7_75t_L g18200 ( 
.A1(n_17895),
.A2(n_8969),
.B1(n_9031),
.B2(n_8951),
.Y(n_18200)
);

INVx4_ASAP7_75t_L g18201 ( 
.A(n_17828),
.Y(n_18201)
);

INVx2_ASAP7_75t_L g18202 ( 
.A(n_17955),
.Y(n_18202)
);

AND2x2_ASAP7_75t_L g18203 ( 
.A(n_18009),
.B(n_8884),
.Y(n_18203)
);

NOR2xp33_ASAP7_75t_L g18204 ( 
.A(n_17754),
.B(n_10841),
.Y(n_18204)
);

NOR2xp33_ASAP7_75t_L g18205 ( 
.A(n_17797),
.B(n_10841),
.Y(n_18205)
);

CKINVDCx20_ASAP7_75t_R g18206 ( 
.A(n_17667),
.Y(n_18206)
);

OR2x2_ASAP7_75t_L g18207 ( 
.A(n_17891),
.B(n_17897),
.Y(n_18207)
);

AND2x4_ASAP7_75t_L g18208 ( 
.A(n_17930),
.B(n_9460),
.Y(n_18208)
);

AND2x2_ASAP7_75t_L g18209 ( 
.A(n_17843),
.B(n_8884),
.Y(n_18209)
);

NAND2xp5_ASAP7_75t_L g18210 ( 
.A(n_17919),
.B(n_10851),
.Y(n_18210)
);

AND2x2_ASAP7_75t_L g18211 ( 
.A(n_17935),
.B(n_8884),
.Y(n_18211)
);

NAND2xp5_ASAP7_75t_L g18212 ( 
.A(n_17925),
.B(n_10851),
.Y(n_18212)
);

AO21x1_ASAP7_75t_L g18213 ( 
.A1(n_17720),
.A2(n_10854),
.B(n_10853),
.Y(n_18213)
);

INVx1_ASAP7_75t_L g18214 ( 
.A(n_17939),
.Y(n_18214)
);

NOR2x1p5_ASAP7_75t_L g18215 ( 
.A(n_17913),
.B(n_9496),
.Y(n_18215)
);

NAND2xp5_ASAP7_75t_L g18216 ( 
.A(n_17946),
.B(n_10853),
.Y(n_18216)
);

AND2x2_ASAP7_75t_L g18217 ( 
.A(n_18033),
.B(n_8897),
.Y(n_18217)
);

OR2x2_ASAP7_75t_L g18218 ( 
.A(n_17953),
.B(n_10854),
.Y(n_18218)
);

AND2x2_ASAP7_75t_L g18219 ( 
.A(n_17779),
.B(n_8897),
.Y(n_18219)
);

INVx2_ASAP7_75t_L g18220 ( 
.A(n_17956),
.Y(n_18220)
);

NAND2xp5_ASAP7_75t_L g18221 ( 
.A(n_17960),
.B(n_10857),
.Y(n_18221)
);

NOR2xp33_ASAP7_75t_L g18222 ( 
.A(n_17716),
.B(n_10857),
.Y(n_18222)
);

AND2x2_ASAP7_75t_L g18223 ( 
.A(n_17818),
.B(n_8897),
.Y(n_18223)
);

AND2x2_ASAP7_75t_L g18224 ( 
.A(n_18082),
.B(n_8897),
.Y(n_18224)
);

AND2x2_ASAP7_75t_L g18225 ( 
.A(n_17910),
.B(n_8897),
.Y(n_18225)
);

NAND2xp5_ASAP7_75t_L g18226 ( 
.A(n_17971),
.B(n_10859),
.Y(n_18226)
);

OAI21xp5_ASAP7_75t_L g18227 ( 
.A1(n_17863),
.A2(n_9716),
.B(n_10844),
.Y(n_18227)
);

AND2x2_ASAP7_75t_L g18228 ( 
.A(n_17912),
.B(n_8897),
.Y(n_18228)
);

OR2x2_ASAP7_75t_L g18229 ( 
.A(n_17848),
.B(n_10859),
.Y(n_18229)
);

INVx1_ASAP7_75t_L g18230 ( 
.A(n_17937),
.Y(n_18230)
);

OAI32xp33_ASAP7_75t_L g18231 ( 
.A1(n_17964),
.A2(n_9214),
.A3(n_9237),
.B1(n_9223),
.B2(n_9207),
.Y(n_18231)
);

INVx1_ASAP7_75t_L g18232 ( 
.A(n_17890),
.Y(n_18232)
);

NOR3xp33_ASAP7_75t_L g18233 ( 
.A(n_17898),
.B(n_9237),
.C(n_9223),
.Y(n_18233)
);

INVx2_ASAP7_75t_SL g18234 ( 
.A(n_17696),
.Y(n_18234)
);

NAND2xp33_ASAP7_75t_R g18235 ( 
.A(n_18075),
.B(n_9237),
.Y(n_18235)
);

INVx1_ASAP7_75t_L g18236 ( 
.A(n_17651),
.Y(n_18236)
);

NOR2xp33_ASAP7_75t_L g18237 ( 
.A(n_17906),
.B(n_10868),
.Y(n_18237)
);

HB1xp67_ASAP7_75t_L g18238 ( 
.A(n_17999),
.Y(n_18238)
);

OR2x2_ASAP7_75t_L g18239 ( 
.A(n_17708),
.B(n_10868),
.Y(n_18239)
);

NAND2xp5_ASAP7_75t_L g18240 ( 
.A(n_17908),
.B(n_10874),
.Y(n_18240)
);

OR2x2_ASAP7_75t_L g18241 ( 
.A(n_17655),
.B(n_10874),
.Y(n_18241)
);

INVx1_ASAP7_75t_L g18242 ( 
.A(n_17782),
.Y(n_18242)
);

NAND2xp5_ASAP7_75t_L g18243 ( 
.A(n_18020),
.B(n_10875),
.Y(n_18243)
);

OR2x2_ASAP7_75t_L g18244 ( 
.A(n_17849),
.B(n_10875),
.Y(n_18244)
);

NAND2xp5_ASAP7_75t_L g18245 ( 
.A(n_17922),
.B(n_10878),
.Y(n_18245)
);

INVx2_ASAP7_75t_L g18246 ( 
.A(n_17677),
.Y(n_18246)
);

HB1xp67_ASAP7_75t_L g18247 ( 
.A(n_17751),
.Y(n_18247)
);

OAI211xp5_ASAP7_75t_L g18248 ( 
.A1(n_17776),
.A2(n_9163),
.B(n_9439),
.C(n_8955),
.Y(n_18248)
);

OAI31xp33_ASAP7_75t_L g18249 ( 
.A1(n_17904),
.A2(n_9281),
.A3(n_9518),
.B(n_9299),
.Y(n_18249)
);

BUFx2_ASAP7_75t_L g18250 ( 
.A(n_17896),
.Y(n_18250)
);

OR2x2_ASAP7_75t_L g18251 ( 
.A(n_17852),
.B(n_10878),
.Y(n_18251)
);

AND2x2_ASAP7_75t_L g18252 ( 
.A(n_17729),
.B(n_8921),
.Y(n_18252)
);

OR2x2_ASAP7_75t_L g18253 ( 
.A(n_17861),
.B(n_10891),
.Y(n_18253)
);

INVx2_ASAP7_75t_L g18254 ( 
.A(n_17677),
.Y(n_18254)
);

AND2x2_ASAP7_75t_L g18255 ( 
.A(n_17748),
.B(n_8921),
.Y(n_18255)
);

NOR4xp25_ASAP7_75t_SL g18256 ( 
.A(n_17771),
.B(n_10891),
.C(n_10896),
.D(n_10894),
.Y(n_18256)
);

NAND2xp5_ASAP7_75t_L g18257 ( 
.A(n_17936),
.B(n_10894),
.Y(n_18257)
);

NOR2xp33_ASAP7_75t_L g18258 ( 
.A(n_17996),
.B(n_10896),
.Y(n_18258)
);

NOR2xp33_ASAP7_75t_R g18259 ( 
.A(n_17767),
.B(n_7049),
.Y(n_18259)
);

NAND2xp5_ASAP7_75t_L g18260 ( 
.A(n_17954),
.B(n_10898),
.Y(n_18260)
);

NAND2xp5_ASAP7_75t_L g18261 ( 
.A(n_17959),
.B(n_10898),
.Y(n_18261)
);

AND2x4_ASAP7_75t_L g18262 ( 
.A(n_17905),
.B(n_9496),
.Y(n_18262)
);

INVx1_ASAP7_75t_L g18263 ( 
.A(n_17998),
.Y(n_18263)
);

AND2x2_ASAP7_75t_L g18264 ( 
.A(n_17654),
.B(n_8921),
.Y(n_18264)
);

AND2x4_ASAP7_75t_L g18265 ( 
.A(n_17911),
.B(n_9496),
.Y(n_18265)
);

INVxp67_ASAP7_75t_SL g18266 ( 
.A(n_17950),
.Y(n_18266)
);

NOR2xp33_ASAP7_75t_L g18267 ( 
.A(n_17773),
.B(n_10902),
.Y(n_18267)
);

AND2x2_ASAP7_75t_L g18268 ( 
.A(n_17792),
.B(n_8921),
.Y(n_18268)
);

AND2x2_ASAP7_75t_L g18269 ( 
.A(n_17799),
.B(n_8921),
.Y(n_18269)
);

OR2x2_ASAP7_75t_L g18270 ( 
.A(n_18016),
.B(n_10902),
.Y(n_18270)
);

NAND2xp5_ASAP7_75t_L g18271 ( 
.A(n_17962),
.B(n_10905),
.Y(n_18271)
);

NAND2xp5_ASAP7_75t_L g18272 ( 
.A(n_17981),
.B(n_10905),
.Y(n_18272)
);

AND2x2_ASAP7_75t_L g18273 ( 
.A(n_17865),
.B(n_8921),
.Y(n_18273)
);

INVx1_ASAP7_75t_L g18274 ( 
.A(n_17847),
.Y(n_18274)
);

OAI221xp5_ASAP7_75t_L g18275 ( 
.A1(n_18079),
.A2(n_9444),
.B1(n_9445),
.B2(n_9286),
.C(n_9280),
.Y(n_18275)
);

OAI33xp33_ASAP7_75t_L g18276 ( 
.A1(n_17738),
.A2(n_10915),
.A3(n_10907),
.B1(n_10919),
.B2(n_10917),
.B3(n_10908),
.Y(n_18276)
);

INVx2_ASAP7_75t_L g18277 ( 
.A(n_17810),
.Y(n_18277)
);

INVx1_ASAP7_75t_SL g18278 ( 
.A(n_17718),
.Y(n_18278)
);

AND2x2_ASAP7_75t_L g18279 ( 
.A(n_17870),
.B(n_17873),
.Y(n_18279)
);

NOR4xp25_ASAP7_75t_SL g18280 ( 
.A(n_17775),
.B(n_10907),
.C(n_10915),
.D(n_10908),
.Y(n_18280)
);

NOR2xp33_ASAP7_75t_L g18281 ( 
.A(n_17815),
.B(n_10917),
.Y(n_18281)
);

AND2x2_ASAP7_75t_L g18282 ( 
.A(n_17877),
.B(n_8922),
.Y(n_18282)
);

INVx1_ASAP7_75t_L g18283 ( 
.A(n_17879),
.Y(n_18283)
);

OR2x2_ASAP7_75t_L g18284 ( 
.A(n_18025),
.B(n_10919),
.Y(n_18284)
);

BUFx2_ASAP7_75t_L g18285 ( 
.A(n_18010),
.Y(n_18285)
);

NOR2x1_ASAP7_75t_L g18286 ( 
.A(n_17881),
.B(n_10922),
.Y(n_18286)
);

HB1xp67_ASAP7_75t_L g18287 ( 
.A(n_18011),
.Y(n_18287)
);

AND2x2_ASAP7_75t_L g18288 ( 
.A(n_17884),
.B(n_8922),
.Y(n_18288)
);

INVx1_ASAP7_75t_L g18289 ( 
.A(n_17740),
.Y(n_18289)
);

INVxp67_ASAP7_75t_L g18290 ( 
.A(n_17710),
.Y(n_18290)
);

A2O1A1Ixp33_ASAP7_75t_L g18291 ( 
.A1(n_17784),
.A2(n_17674),
.B(n_17867),
.C(n_17707),
.Y(n_18291)
);

AND2x4_ASAP7_75t_L g18292 ( 
.A(n_18006),
.B(n_9498),
.Y(n_18292)
);

AND2x2_ASAP7_75t_L g18293 ( 
.A(n_17744),
.B(n_8922),
.Y(n_18293)
);

AND2x2_ASAP7_75t_L g18294 ( 
.A(n_17746),
.B(n_17830),
.Y(n_18294)
);

AND2x2_ASAP7_75t_L g18295 ( 
.A(n_17864),
.B(n_8922),
.Y(n_18295)
);

HB1xp67_ASAP7_75t_L g18296 ( 
.A(n_17687),
.Y(n_18296)
);

INVx2_ASAP7_75t_L g18297 ( 
.A(n_17826),
.Y(n_18297)
);

AND2x2_ASAP7_75t_L g18298 ( 
.A(n_17853),
.B(n_8922),
.Y(n_18298)
);

AOI21xp5_ASAP7_75t_L g18299 ( 
.A1(n_17942),
.A2(n_10928),
.B(n_10922),
.Y(n_18299)
);

INVx2_ASAP7_75t_L g18300 ( 
.A(n_17742),
.Y(n_18300)
);

AOI22xp33_ASAP7_75t_L g18301 ( 
.A1(n_18004),
.A2(n_8969),
.B1(n_9031),
.B2(n_8951),
.Y(n_18301)
);

INVx1_ASAP7_75t_L g18302 ( 
.A(n_17694),
.Y(n_18302)
);

INVx1_ASAP7_75t_L g18303 ( 
.A(n_17724),
.Y(n_18303)
);

INVx1_ASAP7_75t_L g18304 ( 
.A(n_17685),
.Y(n_18304)
);

INVx1_ASAP7_75t_L g18305 ( 
.A(n_17697),
.Y(n_18305)
);

AND2x2_ASAP7_75t_L g18306 ( 
.A(n_17858),
.B(n_8922),
.Y(n_18306)
);

NAND2xp5_ASAP7_75t_L g18307 ( 
.A(n_18024),
.B(n_10928),
.Y(n_18307)
);

BUFx2_ASAP7_75t_L g18308 ( 
.A(n_18024),
.Y(n_18308)
);

INVx2_ASAP7_75t_L g18309 ( 
.A(n_18054),
.Y(n_18309)
);

NOR2xp33_ASAP7_75t_L g18310 ( 
.A(n_18008),
.B(n_10931),
.Y(n_18310)
);

HB1xp67_ASAP7_75t_L g18311 ( 
.A(n_18068),
.Y(n_18311)
);

HB1xp67_ASAP7_75t_L g18312 ( 
.A(n_18012),
.Y(n_18312)
);

AND2x2_ASAP7_75t_L g18313 ( 
.A(n_17878),
.B(n_8975),
.Y(n_18313)
);

AND2x2_ASAP7_75t_L g18314 ( 
.A(n_17882),
.B(n_8975),
.Y(n_18314)
);

HB1xp67_ASAP7_75t_L g18315 ( 
.A(n_17753),
.Y(n_18315)
);

INVx1_ASAP7_75t_L g18316 ( 
.A(n_17761),
.Y(n_18316)
);

NAND2xp5_ASAP7_75t_L g18317 ( 
.A(n_18022),
.B(n_10931),
.Y(n_18317)
);

OR2x2_ASAP7_75t_L g18318 ( 
.A(n_17804),
.B(n_17808),
.Y(n_18318)
);

INVx1_ASAP7_75t_L g18319 ( 
.A(n_17809),
.Y(n_18319)
);

NAND3xp33_ASAP7_75t_SL g18320 ( 
.A(n_18047),
.B(n_9229),
.C(n_9250),
.Y(n_18320)
);

INVxp67_ASAP7_75t_L g18321 ( 
.A(n_18001),
.Y(n_18321)
);

NAND2xp5_ASAP7_75t_L g18322 ( 
.A(n_18081),
.B(n_10937),
.Y(n_18322)
);

NAND2xp5_ASAP7_75t_L g18323 ( 
.A(n_18027),
.B(n_10937),
.Y(n_18323)
);

INVx2_ASAP7_75t_SL g18324 ( 
.A(n_17836),
.Y(n_18324)
);

AND2x2_ASAP7_75t_L g18325 ( 
.A(n_17886),
.B(n_8975),
.Y(n_18325)
);

NOR3xp33_ASAP7_75t_L g18326 ( 
.A(n_18041),
.B(n_9286),
.C(n_9280),
.Y(n_18326)
);

INVx2_ASAP7_75t_L g18327 ( 
.A(n_18054),
.Y(n_18327)
);

INVx2_ASAP7_75t_L g18328 ( 
.A(n_17888),
.Y(n_18328)
);

INVx1_ASAP7_75t_L g18329 ( 
.A(n_17874),
.Y(n_18329)
);

NAND3x1_ASAP7_75t_SL g18330 ( 
.A(n_18015),
.B(n_9405),
.C(n_9377),
.Y(n_18330)
);

INVx1_ASAP7_75t_L g18331 ( 
.A(n_17656),
.Y(n_18331)
);

AND2x2_ASAP7_75t_L g18332 ( 
.A(n_17921),
.B(n_8975),
.Y(n_18332)
);

OR2x2_ASAP7_75t_L g18333 ( 
.A(n_17928),
.B(n_10938),
.Y(n_18333)
);

NOR2xp33_ASAP7_75t_L g18334 ( 
.A(n_17907),
.B(n_10938),
.Y(n_18334)
);

NAND2xp5_ASAP7_75t_L g18335 ( 
.A(n_18073),
.B(n_10941),
.Y(n_18335)
);

INVx1_ASAP7_75t_L g18336 ( 
.A(n_17932),
.Y(n_18336)
);

OR2x2_ASAP7_75t_L g18337 ( 
.A(n_17944),
.B(n_10941),
.Y(n_18337)
);

NAND2xp5_ASAP7_75t_L g18338 ( 
.A(n_17872),
.B(n_10944),
.Y(n_18338)
);

NAND2xp33_ASAP7_75t_R g18339 ( 
.A(n_18048),
.B(n_9280),
.Y(n_18339)
);

NAND2xp5_ASAP7_75t_L g18340 ( 
.A(n_18034),
.B(n_10944),
.Y(n_18340)
);

NOR2x1_ASAP7_75t_L g18341 ( 
.A(n_18045),
.B(n_10945),
.Y(n_18341)
);

INVx2_ASAP7_75t_L g18342 ( 
.A(n_17840),
.Y(n_18342)
);

OAI322xp33_ASAP7_75t_L g18343 ( 
.A1(n_17995),
.A2(n_9445),
.A3(n_9286),
.B1(n_9444),
.B2(n_9280),
.C1(n_9196),
.C2(n_9054),
.Y(n_18343)
);

HB1xp67_ASAP7_75t_L g18344 ( 
.A(n_17658),
.Y(n_18344)
);

OR2x2_ASAP7_75t_L g18345 ( 
.A(n_18052),
.B(n_10945),
.Y(n_18345)
);

OR2x2_ASAP7_75t_L g18346 ( 
.A(n_18057),
.B(n_18058),
.Y(n_18346)
);

NAND2xp5_ASAP7_75t_L g18347 ( 
.A(n_18069),
.B(n_10950),
.Y(n_18347)
);

INVx1_ASAP7_75t_L g18348 ( 
.A(n_17811),
.Y(n_18348)
);

NAND2xp5_ASAP7_75t_L g18349 ( 
.A(n_18076),
.B(n_10950),
.Y(n_18349)
);

AND2x2_ASAP7_75t_L g18350 ( 
.A(n_17982),
.B(n_8975),
.Y(n_18350)
);

INVx1_ASAP7_75t_SL g18351 ( 
.A(n_17984),
.Y(n_18351)
);

INVx1_ASAP7_75t_L g18352 ( 
.A(n_17813),
.Y(n_18352)
);

NAND2xp5_ASAP7_75t_L g18353 ( 
.A(n_18060),
.B(n_18061),
.Y(n_18353)
);

INVx2_ASAP7_75t_L g18354 ( 
.A(n_18026),
.Y(n_18354)
);

OR2x2_ASAP7_75t_L g18355 ( 
.A(n_17883),
.B(n_10951),
.Y(n_18355)
);

OR2x2_ASAP7_75t_L g18356 ( 
.A(n_17926),
.B(n_10951),
.Y(n_18356)
);

AND2x2_ASAP7_75t_L g18357 ( 
.A(n_18003),
.B(n_8975),
.Y(n_18357)
);

INVx2_ASAP7_75t_SL g18358 ( 
.A(n_18064),
.Y(n_18358)
);

NAND2xp5_ASAP7_75t_L g18359 ( 
.A(n_17988),
.B(n_10953),
.Y(n_18359)
);

AND2x4_ASAP7_75t_L g18360 ( 
.A(n_18031),
.B(n_9498),
.Y(n_18360)
);

INVx1_ASAP7_75t_L g18361 ( 
.A(n_17819),
.Y(n_18361)
);

AND2x2_ASAP7_75t_L g18362 ( 
.A(n_17997),
.B(n_8977),
.Y(n_18362)
);

AND2x2_ASAP7_75t_L g18363 ( 
.A(n_18035),
.B(n_8977),
.Y(n_18363)
);

INVx2_ASAP7_75t_L g18364 ( 
.A(n_17693),
.Y(n_18364)
);

NAND2xp5_ASAP7_75t_L g18365 ( 
.A(n_17989),
.B(n_10953),
.Y(n_18365)
);

AND2x4_ASAP7_75t_L g18366 ( 
.A(n_17990),
.B(n_18013),
.Y(n_18366)
);

NAND2xp5_ASAP7_75t_L g18367 ( 
.A(n_18032),
.B(n_10955),
.Y(n_18367)
);

CKINVDCx8_ASAP7_75t_R g18368 ( 
.A(n_17885),
.Y(n_18368)
);

NOR2xp33_ASAP7_75t_L g18369 ( 
.A(n_17822),
.B(n_10955),
.Y(n_18369)
);

NAND2x1p5_ASAP7_75t_L g18370 ( 
.A(n_18029),
.B(n_9163),
.Y(n_18370)
);

NAND2xp5_ASAP7_75t_SL g18371 ( 
.A(n_17733),
.B(n_17760),
.Y(n_18371)
);

NAND2xp5_ASAP7_75t_L g18372 ( 
.A(n_17938),
.B(n_10968),
.Y(n_18372)
);

NOR2xp33_ASAP7_75t_L g18373 ( 
.A(n_17918),
.B(n_10968),
.Y(n_18373)
);

INVx1_ASAP7_75t_L g18374 ( 
.A(n_17772),
.Y(n_18374)
);

NAND2xp5_ASAP7_75t_L g18375 ( 
.A(n_17949),
.B(n_17976),
.Y(n_18375)
);

INVx1_ASAP7_75t_L g18376 ( 
.A(n_17734),
.Y(n_18376)
);

INVx1_ASAP7_75t_L g18377 ( 
.A(n_17941),
.Y(n_18377)
);

AND2x2_ASAP7_75t_L g18378 ( 
.A(n_18078),
.B(n_8977),
.Y(n_18378)
);

OR2x2_ASAP7_75t_L g18379 ( 
.A(n_17974),
.B(n_10975),
.Y(n_18379)
);

INVx1_ASAP7_75t_L g18380 ( 
.A(n_18019),
.Y(n_18380)
);

NAND2xp5_ASAP7_75t_L g18381 ( 
.A(n_17899),
.B(n_10975),
.Y(n_18381)
);

NAND2xp5_ASAP7_75t_L g18382 ( 
.A(n_17909),
.B(n_10977),
.Y(n_18382)
);

NAND4xp25_ASAP7_75t_L g18383 ( 
.A(n_18039),
.B(n_17669),
.C(n_17665),
.D(n_18028),
.Y(n_18383)
);

NAND2xp5_ASAP7_75t_L g18384 ( 
.A(n_18065),
.B(n_10977),
.Y(n_18384)
);

AND2x2_ASAP7_75t_L g18385 ( 
.A(n_18037),
.B(n_18005),
.Y(n_18385)
);

AND2x2_ASAP7_75t_L g18386 ( 
.A(n_17851),
.B(n_8977),
.Y(n_18386)
);

NAND2xp5_ASAP7_75t_L g18387 ( 
.A(n_17814),
.B(n_10979),
.Y(n_18387)
);

INVx1_ASAP7_75t_L g18388 ( 
.A(n_18040),
.Y(n_18388)
);

NAND2xp5_ASAP7_75t_L g18389 ( 
.A(n_17980),
.B(n_10979),
.Y(n_18389)
);

AND2x2_ASAP7_75t_L g18390 ( 
.A(n_17673),
.B(n_8977),
.Y(n_18390)
);

INVx1_ASAP7_75t_L g18391 ( 
.A(n_18046),
.Y(n_18391)
);

OAI321xp33_ASAP7_75t_L g18392 ( 
.A1(n_17679),
.A2(n_17670),
.A3(n_17705),
.B1(n_17806),
.B2(n_17823),
.C(n_17791),
.Y(n_18392)
);

NOR2xp33_ASAP7_75t_R g18393 ( 
.A(n_17824),
.B(n_7049),
.Y(n_18393)
);

NAND2xp5_ASAP7_75t_L g18394 ( 
.A(n_17948),
.B(n_10982),
.Y(n_18394)
);

INVx1_ASAP7_75t_SL g18395 ( 
.A(n_17781),
.Y(n_18395)
);

NOR2xp67_ASAP7_75t_SL g18396 ( 
.A(n_17969),
.B(n_9163),
.Y(n_18396)
);

INVx1_ASAP7_75t_L g18397 ( 
.A(n_18066),
.Y(n_18397)
);

NOR3xp33_ASAP7_75t_SL g18398 ( 
.A(n_17749),
.B(n_17789),
.C(n_17833),
.Y(n_18398)
);

INVx1_ASAP7_75t_L g18399 ( 
.A(n_17957),
.Y(n_18399)
);

NAND2xp5_ASAP7_75t_L g18400 ( 
.A(n_17958),
.B(n_10982),
.Y(n_18400)
);

INVx2_ASAP7_75t_L g18401 ( 
.A(n_17816),
.Y(n_18401)
);

INVx1_ASAP7_75t_L g18402 ( 
.A(n_17965),
.Y(n_18402)
);

NOR2xp33_ASAP7_75t_L g18403 ( 
.A(n_18036),
.B(n_10983),
.Y(n_18403)
);

HB1xp67_ASAP7_75t_L g18404 ( 
.A(n_17834),
.Y(n_18404)
);

NOR2x1p5_ASAP7_75t_L g18405 ( 
.A(n_17841),
.B(n_9498),
.Y(n_18405)
);

BUFx2_ASAP7_75t_L g18406 ( 
.A(n_17842),
.Y(n_18406)
);

AND2x2_ASAP7_75t_L g18407 ( 
.A(n_17947),
.B(n_8977),
.Y(n_18407)
);

INVx2_ASAP7_75t_L g18408 ( 
.A(n_18055),
.Y(n_18408)
);

INVx1_ASAP7_75t_SL g18409 ( 
.A(n_17859),
.Y(n_18409)
);

INVx1_ASAP7_75t_L g18410 ( 
.A(n_18063),
.Y(n_18410)
);

INVxp67_ASAP7_75t_SL g18411 ( 
.A(n_17985),
.Y(n_18411)
);

INVx1_ASAP7_75t_L g18412 ( 
.A(n_17951),
.Y(n_18412)
);

NAND5xp2_ASAP7_75t_SL g18413 ( 
.A(n_17827),
.B(n_9375),
.C(n_9415),
.D(n_9397),
.E(n_9355),
.Y(n_18413)
);

AOI211xp5_ASAP7_75t_L g18414 ( 
.A1(n_17728),
.A2(n_8969),
.B(n_9054),
.C(n_9031),
.Y(n_18414)
);

INVx1_ASAP7_75t_L g18415 ( 
.A(n_17986),
.Y(n_18415)
);

INVx1_ASAP7_75t_L g18416 ( 
.A(n_18002),
.Y(n_18416)
);

AND2x2_ASAP7_75t_L g18417 ( 
.A(n_17952),
.B(n_17933),
.Y(n_18417)
);

NAND2xp5_ASAP7_75t_L g18418 ( 
.A(n_18023),
.B(n_10983),
.Y(n_18418)
);

NAND2xp5_ASAP7_75t_L g18419 ( 
.A(n_18072),
.B(n_10984),
.Y(n_18419)
);

HB1xp67_ASAP7_75t_L g18420 ( 
.A(n_17940),
.Y(n_18420)
);

INVx1_ASAP7_75t_SL g18421 ( 
.A(n_18053),
.Y(n_18421)
);

INVx1_ASAP7_75t_SL g18422 ( 
.A(n_18077),
.Y(n_18422)
);

AND2x2_ASAP7_75t_L g18423 ( 
.A(n_17991),
.B(n_9089),
.Y(n_18423)
);

AOI22xp5_ASAP7_75t_L g18424 ( 
.A1(n_17657),
.A2(n_9031),
.B1(n_9054),
.B2(n_8969),
.Y(n_18424)
);

AND2x2_ASAP7_75t_L g18425 ( 
.A(n_18021),
.B(n_9089),
.Y(n_18425)
);

AND2x2_ASAP7_75t_L g18426 ( 
.A(n_17699),
.B(n_9089),
.Y(n_18426)
);

CKINVDCx5p33_ASAP7_75t_R g18427 ( 
.A(n_17777),
.Y(n_18427)
);

AND2x2_ASAP7_75t_L g18428 ( 
.A(n_17766),
.B(n_9089),
.Y(n_18428)
);

AND2x2_ASAP7_75t_L g18429 ( 
.A(n_17750),
.B(n_9089),
.Y(n_18429)
);

OR2x2_ASAP7_75t_L g18430 ( 
.A(n_17917),
.B(n_10984),
.Y(n_18430)
);

OR2x2_ASAP7_75t_L g18431 ( 
.A(n_17901),
.B(n_10987),
.Y(n_18431)
);

AND2x2_ASAP7_75t_L g18432 ( 
.A(n_18071),
.B(n_9089),
.Y(n_18432)
);

AND2x4_ASAP7_75t_L g18433 ( 
.A(n_17831),
.B(n_9517),
.Y(n_18433)
);

NAND2xp5_ASAP7_75t_SL g18434 ( 
.A(n_17764),
.B(n_9163),
.Y(n_18434)
);

INVxp33_ASAP7_75t_L g18435 ( 
.A(n_17732),
.Y(n_18435)
);

OR2x2_ASAP7_75t_L g18436 ( 
.A(n_17862),
.B(n_10987),
.Y(n_18436)
);

AND2x2_ASAP7_75t_L g18437 ( 
.A(n_18070),
.B(n_9377),
.Y(n_18437)
);

INVx1_ASAP7_75t_L g18438 ( 
.A(n_18056),
.Y(n_18438)
);

NAND2xp5_ASAP7_75t_L g18439 ( 
.A(n_18059),
.B(n_10993),
.Y(n_18439)
);

OR2x2_ASAP7_75t_L g18440 ( 
.A(n_17871),
.B(n_10993),
.Y(n_18440)
);

INVx1_ASAP7_75t_L g18441 ( 
.A(n_18049),
.Y(n_18441)
);

AND2x2_ASAP7_75t_L g18442 ( 
.A(n_17820),
.B(n_9377),
.Y(n_18442)
);

OR2x2_ASAP7_75t_L g18443 ( 
.A(n_17668),
.B(n_10996),
.Y(n_18443)
);

AND2x2_ASAP7_75t_L g18444 ( 
.A(n_17880),
.B(n_9377),
.Y(n_18444)
);

INVx1_ASAP7_75t_L g18445 ( 
.A(n_17803),
.Y(n_18445)
);

NOR2xp33_ASAP7_75t_L g18446 ( 
.A(n_17793),
.B(n_10996),
.Y(n_18446)
);

OR2x2_ASAP7_75t_L g18447 ( 
.A(n_17855),
.B(n_11006),
.Y(n_18447)
);

OR2x2_ASAP7_75t_L g18448 ( 
.A(n_17757),
.B(n_17894),
.Y(n_18448)
);

BUFx2_ASAP7_75t_L g18449 ( 
.A(n_17850),
.Y(n_18449)
);

AND2x2_ASAP7_75t_L g18450 ( 
.A(n_17869),
.B(n_9377),
.Y(n_18450)
);

AND2x4_ASAP7_75t_L g18451 ( 
.A(n_18007),
.B(n_9517),
.Y(n_18451)
);

AND2x2_ASAP7_75t_L g18452 ( 
.A(n_17963),
.B(n_9377),
.Y(n_18452)
);

INVx1_ASAP7_75t_L g18453 ( 
.A(n_17695),
.Y(n_18453)
);

INVx4_ASAP7_75t_L g18454 ( 
.A(n_18062),
.Y(n_18454)
);

AND2x2_ASAP7_75t_L g18455 ( 
.A(n_17934),
.B(n_11006),
.Y(n_18455)
);

INVx1_ASAP7_75t_L g18456 ( 
.A(n_17660),
.Y(n_18456)
);

AND2x2_ASAP7_75t_L g18457 ( 
.A(n_18050),
.B(n_11007),
.Y(n_18457)
);

NAND3xp33_ASAP7_75t_SL g18458 ( 
.A(n_17725),
.B(n_9229),
.C(n_9250),
.Y(n_18458)
);

AND2x2_ASAP7_75t_L g18459 ( 
.A(n_17714),
.B(n_11007),
.Y(n_18459)
);

NAND2xp5_ASAP7_75t_L g18460 ( 
.A(n_17845),
.B(n_11008),
.Y(n_18460)
);

INVx1_ASAP7_75t_L g18461 ( 
.A(n_18080),
.Y(n_18461)
);

INVx1_ASAP7_75t_L g18462 ( 
.A(n_18067),
.Y(n_18462)
);

AND4x1_ASAP7_75t_L g18463 ( 
.A(n_17876),
.B(n_9411),
.C(n_9527),
.D(n_9429),
.Y(n_18463)
);

AOI22xp5_ASAP7_75t_SL g18464 ( 
.A1(n_17973),
.A2(n_9517),
.B1(n_9286),
.B2(n_9444),
.Y(n_18464)
);

INVx1_ASAP7_75t_L g18465 ( 
.A(n_17977),
.Y(n_18465)
);

INVx1_ASAP7_75t_L g18466 ( 
.A(n_17966),
.Y(n_18466)
);

INVx1_ASAP7_75t_L g18467 ( 
.A(n_17807),
.Y(n_18467)
);

AND2x2_ASAP7_75t_L g18468 ( 
.A(n_17709),
.B(n_11008),
.Y(n_18468)
);

NAND2xp5_ASAP7_75t_L g18469 ( 
.A(n_17892),
.B(n_11010),
.Y(n_18469)
);

NAND2xp5_ASAP7_75t_L g18470 ( 
.A(n_17778),
.B(n_11010),
.Y(n_18470)
);

INVx2_ASAP7_75t_L g18471 ( 
.A(n_18018),
.Y(n_18471)
);

AND2x2_ASAP7_75t_L g18472 ( 
.A(n_18042),
.B(n_11011),
.Y(n_18472)
);

INVx1_ASAP7_75t_L g18473 ( 
.A(n_17972),
.Y(n_18473)
);

INVx2_ASAP7_75t_L g18474 ( 
.A(n_17975),
.Y(n_18474)
);

NAND2xp5_ASAP7_75t_L g18475 ( 
.A(n_17770),
.B(n_11011),
.Y(n_18475)
);

OR2x2_ASAP7_75t_L g18476 ( 
.A(n_17866),
.B(n_11012),
.Y(n_18476)
);

AOI211xp5_ASAP7_75t_L g18477 ( 
.A1(n_17923),
.A2(n_8969),
.B(n_9054),
.C(n_9031),
.Y(n_18477)
);

INVx1_ASAP7_75t_L g18478 ( 
.A(n_17762),
.Y(n_18478)
);

AND2x2_ASAP7_75t_L g18479 ( 
.A(n_18044),
.B(n_11012),
.Y(n_18479)
);

NAND2xp5_ASAP7_75t_L g18480 ( 
.A(n_17832),
.B(n_11016),
.Y(n_18480)
);

OR2x2_ASAP7_75t_L g18481 ( 
.A(n_17825),
.B(n_11016),
.Y(n_18481)
);

NOR2xp33_ASAP7_75t_R g18482 ( 
.A(n_17943),
.B(n_7049),
.Y(n_18482)
);

NAND2xp5_ASAP7_75t_L g18483 ( 
.A(n_17983),
.B(n_11022),
.Y(n_18483)
);

INVx1_ASAP7_75t_L g18484 ( 
.A(n_17993),
.Y(n_18484)
);

OAI211xp5_ASAP7_75t_L g18485 ( 
.A1(n_17978),
.A2(n_9439),
.B(n_9163),
.C(n_9286),
.Y(n_18485)
);

INVx1_ASAP7_75t_L g18486 ( 
.A(n_17860),
.Y(n_18486)
);

INVx1_ASAP7_75t_L g18487 ( 
.A(n_18030),
.Y(n_18487)
);

AND2x2_ASAP7_75t_L g18488 ( 
.A(n_17929),
.B(n_11022),
.Y(n_18488)
);

NAND2xp33_ASAP7_75t_R g18489 ( 
.A(n_17968),
.B(n_9280),
.Y(n_18489)
);

NAND2xp33_ASAP7_75t_R g18490 ( 
.A(n_18000),
.B(n_9444),
.Y(n_18490)
);

NOR2xp33_ASAP7_75t_R g18491 ( 
.A(n_17987),
.B(n_7049),
.Y(n_18491)
);

CKINVDCx16_ASAP7_75t_R g18492 ( 
.A(n_18051),
.Y(n_18492)
);

AND2x2_ASAP7_75t_L g18493 ( 
.A(n_17703),
.B(n_9517),
.Y(n_18493)
);

OAI221xp5_ASAP7_75t_L g18494 ( 
.A1(n_17721),
.A2(n_9445),
.B1(n_9444),
.B2(n_9031),
.C(n_9197),
.Y(n_18494)
);

OR2x2_ASAP7_75t_L g18495 ( 
.A(n_17645),
.B(n_9467),
.Y(n_18495)
);

INVxp67_ASAP7_75t_L g18496 ( 
.A(n_17645),
.Y(n_18496)
);

INVx1_ASAP7_75t_L g18497 ( 
.A(n_17645),
.Y(n_18497)
);

AND2x2_ASAP7_75t_L g18498 ( 
.A(n_17703),
.B(n_10844),
.Y(n_18498)
);

INVx1_ASAP7_75t_L g18499 ( 
.A(n_17645),
.Y(n_18499)
);

INVx1_ASAP7_75t_L g18500 ( 
.A(n_18120),
.Y(n_18500)
);

NAND2xp5_ASAP7_75t_L g18501 ( 
.A(n_18122),
.B(n_9222),
.Y(n_18501)
);

HB1xp67_ASAP7_75t_L g18502 ( 
.A(n_18136),
.Y(n_18502)
);

INVx1_ASAP7_75t_SL g18503 ( 
.A(n_18091),
.Y(n_18503)
);

NAND2xp33_ASAP7_75t_SL g18504 ( 
.A(n_18206),
.B(n_7049),
.Y(n_18504)
);

NAND2xp5_ASAP7_75t_L g18505 ( 
.A(n_18122),
.B(n_9222),
.Y(n_18505)
);

OR2x2_ASAP7_75t_L g18506 ( 
.A(n_18147),
.B(n_9564),
.Y(n_18506)
);

OR2x2_ASAP7_75t_L g18507 ( 
.A(n_18083),
.B(n_9574),
.Y(n_18507)
);

INVx1_ASAP7_75t_L g18508 ( 
.A(n_18108),
.Y(n_18508)
);

INVx1_ASAP7_75t_L g18509 ( 
.A(n_18168),
.Y(n_18509)
);

INVxp67_ASAP7_75t_SL g18510 ( 
.A(n_18287),
.Y(n_18510)
);

NAND2xp5_ASAP7_75t_L g18511 ( 
.A(n_18122),
.B(n_18096),
.Y(n_18511)
);

AOI22xp33_ASAP7_75t_L g18512 ( 
.A1(n_18131),
.A2(n_9196),
.B1(n_9197),
.B2(n_9054),
.Y(n_18512)
);

INVx1_ASAP7_75t_SL g18513 ( 
.A(n_18097),
.Y(n_18513)
);

INVx1_ASAP7_75t_L g18514 ( 
.A(n_18250),
.Y(n_18514)
);

INVx1_ASAP7_75t_L g18515 ( 
.A(n_18285),
.Y(n_18515)
);

INVx1_ASAP7_75t_L g18516 ( 
.A(n_18312),
.Y(n_18516)
);

OR2x2_ASAP7_75t_L g18517 ( 
.A(n_18085),
.B(n_9577),
.Y(n_18517)
);

NAND2xp5_ASAP7_75t_L g18518 ( 
.A(n_18165),
.B(n_9222),
.Y(n_18518)
);

NAND2xp5_ASAP7_75t_L g18519 ( 
.A(n_18095),
.B(n_9222),
.Y(n_18519)
);

INVx1_ASAP7_75t_SL g18520 ( 
.A(n_18107),
.Y(n_18520)
);

OR2x2_ASAP7_75t_L g18521 ( 
.A(n_18202),
.B(n_9577),
.Y(n_18521)
);

AND2x2_ASAP7_75t_L g18522 ( 
.A(n_18110),
.B(n_10900),
.Y(n_18522)
);

AND2x2_ASAP7_75t_L g18523 ( 
.A(n_18164),
.B(n_10900),
.Y(n_18523)
);

INVxp67_ASAP7_75t_L g18524 ( 
.A(n_18238),
.Y(n_18524)
);

INVx1_ASAP7_75t_SL g18525 ( 
.A(n_18146),
.Y(n_18525)
);

AND2x2_ASAP7_75t_L g18526 ( 
.A(n_18101),
.B(n_10981),
.Y(n_18526)
);

INVx1_ASAP7_75t_L g18527 ( 
.A(n_18117),
.Y(n_18527)
);

INVxp67_ASAP7_75t_L g18528 ( 
.A(n_18296),
.Y(n_18528)
);

NAND2xp5_ASAP7_75t_L g18529 ( 
.A(n_18084),
.B(n_9244),
.Y(n_18529)
);

AOI22xp33_ASAP7_75t_L g18530 ( 
.A1(n_18157),
.A2(n_9196),
.B1(n_9197),
.B2(n_9054),
.Y(n_18530)
);

NOR2xp33_ASAP7_75t_L g18531 ( 
.A(n_18087),
.B(n_9244),
.Y(n_18531)
);

INVx1_ASAP7_75t_L g18532 ( 
.A(n_18093),
.Y(n_18532)
);

INVx1_ASAP7_75t_L g18533 ( 
.A(n_18124),
.Y(n_18533)
);

AOI222xp33_ASAP7_75t_L g18534 ( 
.A1(n_18127),
.A2(n_9218),
.B1(n_9196),
.B2(n_9315),
.C1(n_9197),
.C2(n_9054),
.Y(n_18534)
);

OR2x6_ASAP7_75t_L g18535 ( 
.A(n_18358),
.B(n_8544),
.Y(n_18535)
);

AND2x4_ASAP7_75t_L g18536 ( 
.A(n_18185),
.B(n_9163),
.Y(n_18536)
);

INVx2_ASAP7_75t_L g18537 ( 
.A(n_18390),
.Y(n_18537)
);

INVxp67_ASAP7_75t_SL g18538 ( 
.A(n_18496),
.Y(n_18538)
);

AND2x2_ASAP7_75t_L g18539 ( 
.A(n_18086),
.B(n_10981),
.Y(n_18539)
);

AND2x2_ASAP7_75t_L g18540 ( 
.A(n_18128),
.B(n_9390),
.Y(n_18540)
);

AND2x2_ASAP7_75t_L g18541 ( 
.A(n_18217),
.B(n_9390),
.Y(n_18541)
);

AOI22xp33_ASAP7_75t_L g18542 ( 
.A1(n_18453),
.A2(n_9196),
.B1(n_9197),
.B2(n_9054),
.Y(n_18542)
);

INVx1_ASAP7_75t_SL g18543 ( 
.A(n_18175),
.Y(n_18543)
);

INVx1_ASAP7_75t_L g18544 ( 
.A(n_18171),
.Y(n_18544)
);

INVxp67_ASAP7_75t_L g18545 ( 
.A(n_18308),
.Y(n_18545)
);

AND3x1_ASAP7_75t_L g18546 ( 
.A(n_18119),
.B(n_9445),
.C(n_7258),
.Y(n_18546)
);

INVx1_ASAP7_75t_L g18547 ( 
.A(n_18497),
.Y(n_18547)
);

INVx1_ASAP7_75t_SL g18548 ( 
.A(n_18130),
.Y(n_18548)
);

NAND2xp5_ASAP7_75t_L g18549 ( 
.A(n_18499),
.B(n_9253),
.Y(n_18549)
);

AND2x2_ASAP7_75t_L g18550 ( 
.A(n_18219),
.B(n_9390),
.Y(n_18550)
);

NAND2xp5_ASAP7_75t_L g18551 ( 
.A(n_18116),
.B(n_9253),
.Y(n_18551)
);

HB1xp67_ASAP7_75t_L g18552 ( 
.A(n_18103),
.Y(n_18552)
);

INVxp67_ASAP7_75t_L g18553 ( 
.A(n_18092),
.Y(n_18553)
);

NOR2xp33_ASAP7_75t_L g18554 ( 
.A(n_18142),
.B(n_9260),
.Y(n_18554)
);

OAI22xp5_ASAP7_75t_L g18555 ( 
.A1(n_18266),
.A2(n_9445),
.B1(n_9196),
.B2(n_9218),
.Y(n_18555)
);

AND2x2_ASAP7_75t_L g18556 ( 
.A(n_18113),
.B(n_9390),
.Y(n_18556)
);

AND2x2_ASAP7_75t_L g18557 ( 
.A(n_18198),
.B(n_9390),
.Y(n_18557)
);

INVx3_ASAP7_75t_L g18558 ( 
.A(n_18155),
.Y(n_18558)
);

INVx1_ASAP7_75t_L g18559 ( 
.A(n_18137),
.Y(n_18559)
);

AOI22xp33_ASAP7_75t_L g18560 ( 
.A1(n_18456),
.A2(n_9197),
.B1(n_9218),
.B2(n_9196),
.Y(n_18560)
);

AND2x2_ASAP7_75t_L g18561 ( 
.A(n_18211),
.B(n_18493),
.Y(n_18561)
);

AND2x2_ASAP7_75t_L g18562 ( 
.A(n_18105),
.B(n_18209),
.Y(n_18562)
);

AND2x2_ASAP7_75t_L g18563 ( 
.A(n_18169),
.B(n_9390),
.Y(n_18563)
);

INVx4_ASAP7_75t_L g18564 ( 
.A(n_18201),
.Y(n_18564)
);

AOI22xp5_ASAP7_75t_L g18565 ( 
.A1(n_18104),
.A2(n_9196),
.B1(n_9218),
.B2(n_9197),
.Y(n_18565)
);

BUFx2_ASAP7_75t_L g18566 ( 
.A(n_18155),
.Y(n_18566)
);

NOR2x1p5_ASAP7_75t_L g18567 ( 
.A(n_18100),
.B(n_9197),
.Y(n_18567)
);

AOI22xp5_ASAP7_75t_L g18568 ( 
.A1(n_18474),
.A2(n_9218),
.B1(n_9335),
.B2(n_9315),
.Y(n_18568)
);

INVx1_ASAP7_75t_L g18569 ( 
.A(n_18279),
.Y(n_18569)
);

INVx1_ASAP7_75t_L g18570 ( 
.A(n_18158),
.Y(n_18570)
);

INVx3_ASAP7_75t_SL g18571 ( 
.A(n_18366),
.Y(n_18571)
);

INVx1_ASAP7_75t_L g18572 ( 
.A(n_18160),
.Y(n_18572)
);

AOI21xp5_ASAP7_75t_L g18573 ( 
.A1(n_18183),
.A2(n_9372),
.B(n_9371),
.Y(n_18573)
);

HB1xp67_ASAP7_75t_L g18574 ( 
.A(n_18247),
.Y(n_18574)
);

INVx1_ASAP7_75t_L g18575 ( 
.A(n_18315),
.Y(n_18575)
);

AND2x2_ASAP7_75t_L g18576 ( 
.A(n_18144),
.B(n_9390),
.Y(n_18576)
);

INVx2_ASAP7_75t_SL g18577 ( 
.A(n_18148),
.Y(n_18577)
);

INVx1_ASAP7_75t_L g18578 ( 
.A(n_18207),
.Y(n_18578)
);

NAND2xp5_ASAP7_75t_SL g18579 ( 
.A(n_18109),
.B(n_9163),
.Y(n_18579)
);

NAND2xp5_ASAP7_75t_L g18580 ( 
.A(n_18351),
.B(n_9260),
.Y(n_18580)
);

NAND2xp5_ASAP7_75t_L g18581 ( 
.A(n_18321),
.B(n_9260),
.Y(n_18581)
);

OR2x2_ASAP7_75t_L g18582 ( 
.A(n_18094),
.B(n_9371),
.Y(n_18582)
);

INVx1_ASAP7_75t_SL g18583 ( 
.A(n_18114),
.Y(n_18583)
);

INVx1_ASAP7_75t_SL g18584 ( 
.A(n_18089),
.Y(n_18584)
);

INVx1_ASAP7_75t_L g18585 ( 
.A(n_18194),
.Y(n_18585)
);

INVx2_ASAP7_75t_L g18586 ( 
.A(n_18425),
.Y(n_18586)
);

NAND2xp5_ASAP7_75t_SL g18587 ( 
.A(n_18492),
.B(n_9163),
.Y(n_18587)
);

AOI22xp33_ASAP7_75t_L g18588 ( 
.A1(n_18438),
.A2(n_9315),
.B1(n_9335),
.B2(n_9218),
.Y(n_18588)
);

BUFx3_ASAP7_75t_L g18589 ( 
.A(n_18162),
.Y(n_18589)
);

NOR2xp33_ASAP7_75t_L g18590 ( 
.A(n_18278),
.B(n_9260),
.Y(n_18590)
);

NAND2x1_ASAP7_75t_L g18591 ( 
.A(n_18102),
.B(n_8995),
.Y(n_18591)
);

BUFx4f_ASAP7_75t_L g18592 ( 
.A(n_18199),
.Y(n_18592)
);

INVx1_ASAP7_75t_SL g18593 ( 
.A(n_18294),
.Y(n_18593)
);

AOI221xp5_ASAP7_75t_L g18594 ( 
.A1(n_18392),
.A2(n_8993),
.B1(n_9335),
.B2(n_9315),
.C(n_9218),
.Y(n_18594)
);

AND2x2_ASAP7_75t_L g18595 ( 
.A(n_18255),
.B(n_9390),
.Y(n_18595)
);

INVx2_ASAP7_75t_L g18596 ( 
.A(n_18346),
.Y(n_18596)
);

NAND2x1p5_ASAP7_75t_L g18597 ( 
.A(n_18090),
.B(n_9439),
.Y(n_18597)
);

NAND2xp5_ASAP7_75t_L g18598 ( 
.A(n_18395),
.B(n_9260),
.Y(n_18598)
);

INVx2_ASAP7_75t_SL g18599 ( 
.A(n_18215),
.Y(n_18599)
);

INVx1_ASAP7_75t_L g18600 ( 
.A(n_18213),
.Y(n_18600)
);

OR2x2_ASAP7_75t_L g18601 ( 
.A(n_18118),
.B(n_9372),
.Y(n_18601)
);

OR2x2_ASAP7_75t_L g18602 ( 
.A(n_18151),
.B(n_9374),
.Y(n_18602)
);

INVx1_ASAP7_75t_SL g18603 ( 
.A(n_18318),
.Y(n_18603)
);

INVx1_ASAP7_75t_SL g18604 ( 
.A(n_18125),
.Y(n_18604)
);

AND2x2_ASAP7_75t_L g18605 ( 
.A(n_18225),
.B(n_9423),
.Y(n_18605)
);

AND2x2_ASAP7_75t_L g18606 ( 
.A(n_18228),
.B(n_9423),
.Y(n_18606)
);

INVxp33_ASAP7_75t_L g18607 ( 
.A(n_18123),
.Y(n_18607)
);

NAND2xp5_ASAP7_75t_L g18608 ( 
.A(n_18409),
.B(n_9319),
.Y(n_18608)
);

NAND2xp5_ASAP7_75t_L g18609 ( 
.A(n_18406),
.B(n_9319),
.Y(n_18609)
);

INVx1_ASAP7_75t_L g18610 ( 
.A(n_18115),
.Y(n_18610)
);

AND2x2_ASAP7_75t_L g18611 ( 
.A(n_18273),
.B(n_9423),
.Y(n_18611)
);

INVx1_ASAP7_75t_SL g18612 ( 
.A(n_18197),
.Y(n_18612)
);

AND2x2_ASAP7_75t_L g18613 ( 
.A(n_18282),
.B(n_9423),
.Y(n_18613)
);

AO21x2_ASAP7_75t_L g18614 ( 
.A1(n_18181),
.A2(n_10998),
.B(n_10990),
.Y(n_18614)
);

NOR2x1_ASAP7_75t_L g18615 ( 
.A(n_18232),
.B(n_9561),
.Y(n_18615)
);

INVx2_ASAP7_75t_L g18616 ( 
.A(n_18166),
.Y(n_18616)
);

AND2x2_ASAP7_75t_L g18617 ( 
.A(n_18288),
.B(n_9423),
.Y(n_18617)
);

INVx1_ASAP7_75t_L g18618 ( 
.A(n_18404),
.Y(n_18618)
);

OR2x2_ASAP7_75t_L g18619 ( 
.A(n_18172),
.B(n_9374),
.Y(n_18619)
);

INVx1_ASAP7_75t_L g18620 ( 
.A(n_18344),
.Y(n_18620)
);

NAND2x1_ASAP7_75t_L g18621 ( 
.A(n_18102),
.B(n_8995),
.Y(n_18621)
);

INVx2_ASAP7_75t_L g18622 ( 
.A(n_18370),
.Y(n_18622)
);

INVx2_ASAP7_75t_L g18623 ( 
.A(n_18426),
.Y(n_18623)
);

OAI22xp5_ASAP7_75t_SL g18624 ( 
.A1(n_18368),
.A2(n_18324),
.B1(n_18236),
.B2(n_18303),
.Y(n_18624)
);

CKINVDCx16_ASAP7_75t_R g18625 ( 
.A(n_18311),
.Y(n_18625)
);

OR2x2_ASAP7_75t_L g18626 ( 
.A(n_18342),
.B(n_9392),
.Y(n_18626)
);

NAND2xp5_ASAP7_75t_L g18627 ( 
.A(n_18246),
.B(n_9319),
.Y(n_18627)
);

OR2x2_ASAP7_75t_L g18628 ( 
.A(n_18495),
.B(n_9392),
.Y(n_18628)
);

NOR2xp33_ASAP7_75t_L g18629 ( 
.A(n_18454),
.B(n_9319),
.Y(n_18629)
);

INVx1_ASAP7_75t_SL g18630 ( 
.A(n_18126),
.Y(n_18630)
);

NOR2x1_ASAP7_75t_L g18631 ( 
.A(n_18242),
.B(n_9433),
.Y(n_18631)
);

HB1xp67_ASAP7_75t_L g18632 ( 
.A(n_18186),
.Y(n_18632)
);

AND2x4_ASAP7_75t_L g18633 ( 
.A(n_18234),
.B(n_9439),
.Y(n_18633)
);

INVx1_ASAP7_75t_L g18634 ( 
.A(n_18297),
.Y(n_18634)
);

INVx2_ASAP7_75t_L g18635 ( 
.A(n_18141),
.Y(n_18635)
);

AND2x4_ASAP7_75t_L g18636 ( 
.A(n_18385),
.B(n_9439),
.Y(n_18636)
);

INVx1_ASAP7_75t_L g18637 ( 
.A(n_18328),
.Y(n_18637)
);

INVx1_ASAP7_75t_L g18638 ( 
.A(n_18254),
.Y(n_18638)
);

NAND2xp5_ASAP7_75t_L g18639 ( 
.A(n_18411),
.B(n_18121),
.Y(n_18639)
);

AND2x4_ASAP7_75t_L g18640 ( 
.A(n_18184),
.B(n_9439),
.Y(n_18640)
);

NAND2xp5_ASAP7_75t_L g18641 ( 
.A(n_18224),
.B(n_9319),
.Y(n_18641)
);

NOR2xp33_ASAP7_75t_L g18642 ( 
.A(n_18163),
.B(n_9357),
.Y(n_18642)
);

AND2x2_ASAP7_75t_L g18643 ( 
.A(n_18295),
.B(n_9423),
.Y(n_18643)
);

INVx2_ASAP7_75t_L g18644 ( 
.A(n_18405),
.Y(n_18644)
);

NAND2xp5_ASAP7_75t_L g18645 ( 
.A(n_18408),
.B(n_9357),
.Y(n_18645)
);

OR2x2_ASAP7_75t_L g18646 ( 
.A(n_18283),
.B(n_9394),
.Y(n_18646)
);

INVx4_ASAP7_75t_L g18647 ( 
.A(n_18427),
.Y(n_18647)
);

INVx2_ASAP7_75t_L g18648 ( 
.A(n_18132),
.Y(n_18648)
);

AND2x2_ASAP7_75t_L g18649 ( 
.A(n_18252),
.B(n_9423),
.Y(n_18649)
);

AND2x2_ASAP7_75t_SL g18650 ( 
.A(n_18187),
.B(n_9218),
.Y(n_18650)
);

INVx1_ASAP7_75t_L g18651 ( 
.A(n_18353),
.Y(n_18651)
);

AO22x1_ASAP7_75t_L g18652 ( 
.A1(n_18274),
.A2(n_7355),
.B1(n_7543),
.B2(n_7232),
.Y(n_18652)
);

INVx1_ASAP7_75t_L g18653 ( 
.A(n_18375),
.Y(n_18653)
);

OAI22xp5_ASAP7_75t_L g18654 ( 
.A1(n_18143),
.A2(n_18230),
.B1(n_18214),
.B2(n_18263),
.Y(n_18654)
);

INVx1_ASAP7_75t_L g18655 ( 
.A(n_18223),
.Y(n_18655)
);

AND2x2_ASAP7_75t_L g18656 ( 
.A(n_18149),
.B(n_9423),
.Y(n_18656)
);

AND2x2_ASAP7_75t_L g18657 ( 
.A(n_18174),
.B(n_10990),
.Y(n_18657)
);

OR2x2_ASAP7_75t_L g18658 ( 
.A(n_18277),
.B(n_9394),
.Y(n_18658)
);

INVx1_ASAP7_75t_L g18659 ( 
.A(n_18192),
.Y(n_18659)
);

AND2x2_ASAP7_75t_L g18660 ( 
.A(n_18176),
.B(n_10990),
.Y(n_18660)
);

OAI22xp5_ASAP7_75t_L g18661 ( 
.A1(n_18319),
.A2(n_9335),
.B1(n_9336),
.B2(n_9315),
.Y(n_18661)
);

AND2x2_ASAP7_75t_L g18662 ( 
.A(n_18178),
.B(n_10998),
.Y(n_18662)
);

INVx1_ASAP7_75t_L g18663 ( 
.A(n_18193),
.Y(n_18663)
);

HB1xp67_ASAP7_75t_L g18664 ( 
.A(n_18265),
.Y(n_18664)
);

OAI22xp5_ASAP7_75t_L g18665 ( 
.A1(n_18336),
.A2(n_9335),
.B1(n_9336),
.B2(n_9315),
.Y(n_18665)
);

INVx2_ASAP7_75t_L g18666 ( 
.A(n_18265),
.Y(n_18666)
);

NOR2xp33_ASAP7_75t_L g18667 ( 
.A(n_18302),
.B(n_9357),
.Y(n_18667)
);

AND2x2_ASAP7_75t_L g18668 ( 
.A(n_18386),
.B(n_18357),
.Y(n_18668)
);

OR2x2_ASAP7_75t_L g18669 ( 
.A(n_18161),
.B(n_9408),
.Y(n_18669)
);

INVx1_ASAP7_75t_L g18670 ( 
.A(n_18397),
.Y(n_18670)
);

INVx1_ASAP7_75t_L g18671 ( 
.A(n_18410),
.Y(n_18671)
);

NOR2x1_ASAP7_75t_L g18672 ( 
.A(n_18329),
.B(n_9433),
.Y(n_18672)
);

INVx1_ASAP7_75t_SL g18673 ( 
.A(n_18422),
.Y(n_18673)
);

NAND2xp5_ASAP7_75t_L g18674 ( 
.A(n_18208),
.B(n_9357),
.Y(n_18674)
);

INVx2_ASAP7_75t_L g18675 ( 
.A(n_18292),
.Y(n_18675)
);

INVx2_ASAP7_75t_L g18676 ( 
.A(n_18292),
.Y(n_18676)
);

OR2x2_ASAP7_75t_L g18677 ( 
.A(n_18167),
.B(n_9408),
.Y(n_18677)
);

NAND2xp5_ASAP7_75t_L g18678 ( 
.A(n_18208),
.B(n_9357),
.Y(n_18678)
);

OR2x2_ASAP7_75t_L g18679 ( 
.A(n_18170),
.B(n_9409),
.Y(n_18679)
);

OR2x2_ASAP7_75t_L g18680 ( 
.A(n_18134),
.B(n_9409),
.Y(n_18680)
);

NAND2xp5_ASAP7_75t_L g18681 ( 
.A(n_18380),
.B(n_9373),
.Y(n_18681)
);

AOI22xp33_ASAP7_75t_L g18682 ( 
.A1(n_18441),
.A2(n_9335),
.B1(n_9336),
.B2(n_9315),
.Y(n_18682)
);

OR2x6_ASAP7_75t_L g18683 ( 
.A(n_18316),
.B(n_8544),
.Y(n_18683)
);

OR2x2_ASAP7_75t_L g18684 ( 
.A(n_18309),
.B(n_7255),
.Y(n_18684)
);

INVx2_ASAP7_75t_L g18685 ( 
.A(n_18262),
.Y(n_18685)
);

INVxp67_ASAP7_75t_L g18686 ( 
.A(n_18098),
.Y(n_18686)
);

HB1xp67_ASAP7_75t_L g18687 ( 
.A(n_18220),
.Y(n_18687)
);

NAND2x1_ASAP7_75t_SL g18688 ( 
.A(n_18420),
.B(n_7232),
.Y(n_18688)
);

AOI22xp33_ASAP7_75t_L g18689 ( 
.A1(n_18462),
.A2(n_9335),
.B1(n_9336),
.B2(n_9315),
.Y(n_18689)
);

INVx1_ASAP7_75t_SL g18690 ( 
.A(n_18421),
.Y(n_18690)
);

AND2x2_ASAP7_75t_L g18691 ( 
.A(n_18150),
.B(n_10998),
.Y(n_18691)
);

INVx1_ASAP7_75t_L g18692 ( 
.A(n_18388),
.Y(n_18692)
);

CKINVDCx16_ASAP7_75t_R g18693 ( 
.A(n_18112),
.Y(n_18693)
);

INVx1_ASAP7_75t_L g18694 ( 
.A(n_18391),
.Y(n_18694)
);

INVx1_ASAP7_75t_L g18695 ( 
.A(n_18412),
.Y(n_18695)
);

NAND2xp5_ASAP7_75t_L g18696 ( 
.A(n_18327),
.B(n_9373),
.Y(n_18696)
);

NAND2xp5_ASAP7_75t_L g18697 ( 
.A(n_18111),
.B(n_9373),
.Y(n_18697)
);

AND2x2_ASAP7_75t_L g18698 ( 
.A(n_18354),
.B(n_11001),
.Y(n_18698)
);

NAND2xp5_ASAP7_75t_SL g18699 ( 
.A(n_18189),
.B(n_9439),
.Y(n_18699)
);

INVx2_ASAP7_75t_L g18700 ( 
.A(n_18442),
.Y(n_18700)
);

INVx1_ASAP7_75t_L g18701 ( 
.A(n_18270),
.Y(n_18701)
);

INVx1_ASAP7_75t_SL g18702 ( 
.A(n_18259),
.Y(n_18702)
);

INVx1_ASAP7_75t_SL g18703 ( 
.A(n_18129),
.Y(n_18703)
);

NAND2xp5_ASAP7_75t_L g18704 ( 
.A(n_18289),
.B(n_9373),
.Y(n_18704)
);

CKINVDCx16_ASAP7_75t_R g18705 ( 
.A(n_18159),
.Y(n_18705)
);

BUFx2_ASAP7_75t_L g18706 ( 
.A(n_18393),
.Y(n_18706)
);

CKINVDCx16_ASAP7_75t_R g18707 ( 
.A(n_18399),
.Y(n_18707)
);

AND3x1_ASAP7_75t_L g18708 ( 
.A(n_18398),
.B(n_7258),
.C(n_7244),
.Y(n_18708)
);

NOR2x1_ASAP7_75t_L g18709 ( 
.A(n_18374),
.B(n_9380),
.Y(n_18709)
);

AND2x2_ASAP7_75t_L g18710 ( 
.A(n_18195),
.B(n_18428),
.Y(n_18710)
);

INVx1_ASAP7_75t_L g18711 ( 
.A(n_18284),
.Y(n_18711)
);

INVx1_ASAP7_75t_L g18712 ( 
.A(n_18286),
.Y(n_18712)
);

NAND2xp5_ASAP7_75t_L g18713 ( 
.A(n_18304),
.B(n_9373),
.Y(n_18713)
);

OR2x2_ASAP7_75t_L g18714 ( 
.A(n_18152),
.B(n_7271),
.Y(n_18714)
);

OR2x2_ASAP7_75t_L g18715 ( 
.A(n_18245),
.B(n_7271),
.Y(n_18715)
);

INVx1_ASAP7_75t_L g18716 ( 
.A(n_18135),
.Y(n_18716)
);

INVx1_ASAP7_75t_SL g18717 ( 
.A(n_18305),
.Y(n_18717)
);

INVx1_ASAP7_75t_L g18718 ( 
.A(n_18341),
.Y(n_18718)
);

AND2x2_ASAP7_75t_L g18719 ( 
.A(n_18423),
.B(n_11001),
.Y(n_18719)
);

INVx1_ASAP7_75t_L g18720 ( 
.A(n_18229),
.Y(n_18720)
);

AND2x2_ASAP7_75t_L g18721 ( 
.A(n_18203),
.B(n_18362),
.Y(n_18721)
);

INVx1_ASAP7_75t_L g18722 ( 
.A(n_18218),
.Y(n_18722)
);

INVx2_ASAP7_75t_L g18723 ( 
.A(n_18293),
.Y(n_18723)
);

INVx1_ASAP7_75t_L g18724 ( 
.A(n_18244),
.Y(n_18724)
);

AND2x2_ASAP7_75t_L g18725 ( 
.A(n_18417),
.B(n_11001),
.Y(n_18725)
);

INVx1_ASAP7_75t_L g18726 ( 
.A(n_18251),
.Y(n_18726)
);

INVx3_ASAP7_75t_L g18727 ( 
.A(n_18360),
.Y(n_18727)
);

NOR2x1_ASAP7_75t_L g18728 ( 
.A(n_18331),
.B(n_9380),
.Y(n_18728)
);

INVx1_ASAP7_75t_L g18729 ( 
.A(n_18253),
.Y(n_18729)
);

NOR2xp33_ASAP7_75t_L g18730 ( 
.A(n_18383),
.B(n_8341),
.Y(n_18730)
);

AND2x2_ASAP7_75t_L g18731 ( 
.A(n_18298),
.B(n_6946),
.Y(n_18731)
);

CKINVDCx16_ASAP7_75t_R g18732 ( 
.A(n_18402),
.Y(n_18732)
);

INVx1_ASAP7_75t_L g18733 ( 
.A(n_18330),
.Y(n_18733)
);

AND2x2_ASAP7_75t_L g18734 ( 
.A(n_18306),
.B(n_6946),
.Y(n_18734)
);

AOI222xp33_ASAP7_75t_L g18735 ( 
.A1(n_18099),
.A2(n_9507),
.B1(n_9336),
.B2(n_9404),
.C1(n_9335),
.C2(n_8186),
.Y(n_18735)
);

INVx2_ASAP7_75t_L g18736 ( 
.A(n_18452),
.Y(n_18736)
);

INVx2_ASAP7_75t_L g18737 ( 
.A(n_18345),
.Y(n_18737)
);

HB1xp67_ASAP7_75t_L g18738 ( 
.A(n_18300),
.Y(n_18738)
);

OR2x2_ASAP7_75t_L g18739 ( 
.A(n_18257),
.B(n_7287),
.Y(n_18739)
);

INVx1_ASAP7_75t_L g18740 ( 
.A(n_18240),
.Y(n_18740)
);

INVxp67_ASAP7_75t_L g18741 ( 
.A(n_18377),
.Y(n_18741)
);

INVx1_ASAP7_75t_SL g18742 ( 
.A(n_18416),
.Y(n_18742)
);

INVx2_ASAP7_75t_L g18743 ( 
.A(n_18356),
.Y(n_18743)
);

NAND2xp5_ASAP7_75t_SL g18744 ( 
.A(n_18088),
.B(n_18364),
.Y(n_18744)
);

INVx1_ASAP7_75t_SL g18745 ( 
.A(n_18348),
.Y(n_18745)
);

AND2x4_ASAP7_75t_L g18746 ( 
.A(n_18268),
.B(n_9439),
.Y(n_18746)
);

AND2x4_ASAP7_75t_L g18747 ( 
.A(n_18269),
.B(n_10474),
.Y(n_18747)
);

INVx1_ASAP7_75t_L g18748 ( 
.A(n_18379),
.Y(n_18748)
);

INVx2_ASAP7_75t_SL g18749 ( 
.A(n_18190),
.Y(n_18749)
);

NAND2xp5_ASAP7_75t_L g18750 ( 
.A(n_18352),
.B(n_8341),
.Y(n_18750)
);

AND2x2_ASAP7_75t_L g18751 ( 
.A(n_18313),
.B(n_6946),
.Y(n_18751)
);

INVx1_ASAP7_75t_L g18752 ( 
.A(n_18212),
.Y(n_18752)
);

OAI31xp33_ASAP7_75t_SL g18753 ( 
.A1(n_18173),
.A2(n_10160),
.A3(n_10459),
.B(n_10144),
.Y(n_18753)
);

INVx1_ASAP7_75t_SL g18754 ( 
.A(n_18361),
.Y(n_18754)
);

NAND2xp5_ASAP7_75t_L g18755 ( 
.A(n_18415),
.B(n_18222),
.Y(n_18755)
);

AND2x2_ASAP7_75t_L g18756 ( 
.A(n_18314),
.B(n_6946),
.Y(n_18756)
);

NAND2xp5_ASAP7_75t_L g18757 ( 
.A(n_18461),
.B(n_8341),
.Y(n_18757)
);

INVx2_ASAP7_75t_L g18758 ( 
.A(n_18355),
.Y(n_18758)
);

INVx1_ASAP7_75t_L g18759 ( 
.A(n_18239),
.Y(n_18759)
);

AND2x2_ASAP7_75t_L g18760 ( 
.A(n_18325),
.B(n_18332),
.Y(n_18760)
);

INVx1_ASAP7_75t_L g18761 ( 
.A(n_18337),
.Y(n_18761)
);

BUFx6f_ASAP7_75t_L g18762 ( 
.A(n_18376),
.Y(n_18762)
);

OR2x2_ASAP7_75t_L g18763 ( 
.A(n_18260),
.B(n_7287),
.Y(n_18763)
);

INVx1_ASAP7_75t_L g18764 ( 
.A(n_18241),
.Y(n_18764)
);

OAI22xp5_ASAP7_75t_L g18765 ( 
.A1(n_18467),
.A2(n_9336),
.B1(n_9507),
.B2(n_9404),
.Y(n_18765)
);

AND2x2_ASAP7_75t_L g18766 ( 
.A(n_18350),
.B(n_6979),
.Y(n_18766)
);

NOR2xp33_ASAP7_75t_L g18767 ( 
.A(n_18435),
.B(n_8341),
.Y(n_18767)
);

INVx1_ASAP7_75t_SL g18768 ( 
.A(n_18401),
.Y(n_18768)
);

NOR2xp33_ASAP7_75t_L g18769 ( 
.A(n_18449),
.B(n_8342),
.Y(n_18769)
);

AND2x2_ASAP7_75t_L g18770 ( 
.A(n_18264),
.B(n_6979),
.Y(n_18770)
);

NOR2xp67_ASAP7_75t_L g18771 ( 
.A(n_18290),
.B(n_18156),
.Y(n_18771)
);

INVx1_ASAP7_75t_L g18772 ( 
.A(n_18381),
.Y(n_18772)
);

INVx1_ASAP7_75t_L g18773 ( 
.A(n_18382),
.Y(n_18773)
);

INVx2_ASAP7_75t_L g18774 ( 
.A(n_18498),
.Y(n_18774)
);

AND2x2_ASAP7_75t_L g18775 ( 
.A(n_18363),
.B(n_18378),
.Y(n_18775)
);

OAI22xp5_ASAP7_75t_L g18776 ( 
.A1(n_18473),
.A2(n_9336),
.B1(n_9507),
.B2(n_9404),
.Y(n_18776)
);

NAND2xp5_ASAP7_75t_L g18777 ( 
.A(n_18310),
.B(n_8342),
.Y(n_18777)
);

NOR3xp33_ASAP7_75t_L g18778 ( 
.A(n_18106),
.B(n_8444),
.C(n_9307),
.Y(n_18778)
);

INVx1_ASAP7_75t_L g18779 ( 
.A(n_18261),
.Y(n_18779)
);

BUFx2_ASAP7_75t_L g18780 ( 
.A(n_18486),
.Y(n_18780)
);

NAND2xp5_ASAP7_75t_L g18781 ( 
.A(n_18205),
.B(n_18237),
.Y(n_18781)
);

INVx2_ASAP7_75t_SL g18782 ( 
.A(n_18271),
.Y(n_18782)
);

AND2x2_ASAP7_75t_L g18783 ( 
.A(n_18407),
.B(n_6979),
.Y(n_18783)
);

INVx1_ASAP7_75t_L g18784 ( 
.A(n_18272),
.Y(n_18784)
);

AND2x2_ASAP7_75t_L g18785 ( 
.A(n_18437),
.B(n_6979),
.Y(n_18785)
);

INVxp67_ASAP7_75t_L g18786 ( 
.A(n_18267),
.Y(n_18786)
);

INVx1_ASAP7_75t_SL g18787 ( 
.A(n_18468),
.Y(n_18787)
);

INVx1_ASAP7_75t_SL g18788 ( 
.A(n_18153),
.Y(n_18788)
);

INVx1_ASAP7_75t_SL g18789 ( 
.A(n_18210),
.Y(n_18789)
);

AND2x2_ASAP7_75t_L g18790 ( 
.A(n_18484),
.B(n_6981),
.Y(n_18790)
);

INVx1_ASAP7_75t_SL g18791 ( 
.A(n_18371),
.Y(n_18791)
);

NAND2xp5_ASAP7_75t_L g18792 ( 
.A(n_18179),
.B(n_8342),
.Y(n_18792)
);

NOR2xp33_ASAP7_75t_L g18793 ( 
.A(n_18448),
.B(n_18445),
.Y(n_18793)
);

INVx1_ASAP7_75t_L g18794 ( 
.A(n_18333),
.Y(n_18794)
);

AOI222xp33_ASAP7_75t_L g18795 ( 
.A1(n_18446),
.A2(n_9404),
.B1(n_9507),
.B2(n_9336),
.C1(n_8186),
.C2(n_8168),
.Y(n_18795)
);

OR2x2_ASAP7_75t_L g18796 ( 
.A(n_18291),
.B(n_7306),
.Y(n_18796)
);

AND2x2_ASAP7_75t_L g18797 ( 
.A(n_18487),
.B(n_6981),
.Y(n_18797)
);

INVx1_ASAP7_75t_L g18798 ( 
.A(n_18372),
.Y(n_18798)
);

INVx1_ASAP7_75t_L g18799 ( 
.A(n_18394),
.Y(n_18799)
);

AND2x2_ASAP7_75t_L g18800 ( 
.A(n_18463),
.B(n_6981),
.Y(n_18800)
);

INVx1_ASAP7_75t_SL g18801 ( 
.A(n_18243),
.Y(n_18801)
);

INVx3_ASAP7_75t_L g18802 ( 
.A(n_18433),
.Y(n_18802)
);

INVxp67_ASAP7_75t_L g18803 ( 
.A(n_18281),
.Y(n_18803)
);

INVx2_ASAP7_75t_L g18804 ( 
.A(n_18455),
.Y(n_18804)
);

AND2x2_ASAP7_75t_L g18805 ( 
.A(n_18444),
.B(n_18450),
.Y(n_18805)
);

INVx1_ASAP7_75t_L g18806 ( 
.A(n_18400),
.Y(n_18806)
);

AND2x4_ASAP7_75t_L g18807 ( 
.A(n_18466),
.B(n_10474),
.Y(n_18807)
);

AOI222xp33_ASAP7_75t_L g18808 ( 
.A1(n_18369),
.A2(n_9507),
.B1(n_9404),
.B2(n_8186),
.C1(n_8168),
.C2(n_8227),
.Y(n_18808)
);

INVx1_ASAP7_75t_L g18809 ( 
.A(n_18389),
.Y(n_18809)
);

OR2x2_ASAP7_75t_L g18810 ( 
.A(n_18177),
.B(n_7306),
.Y(n_18810)
);

INVx2_ASAP7_75t_L g18811 ( 
.A(n_18431),
.Y(n_18811)
);

INVx1_ASAP7_75t_L g18812 ( 
.A(n_18317),
.Y(n_18812)
);

AND2x2_ASAP7_75t_L g18813 ( 
.A(n_18396),
.B(n_6981),
.Y(n_18813)
);

INVx1_ASAP7_75t_L g18814 ( 
.A(n_18323),
.Y(n_18814)
);

OR2x2_ASAP7_75t_L g18815 ( 
.A(n_18322),
.B(n_7306),
.Y(n_18815)
);

INVx2_ASAP7_75t_L g18816 ( 
.A(n_18436),
.Y(n_18816)
);

OAI22xp5_ASAP7_75t_L g18817 ( 
.A1(n_18180),
.A2(n_9507),
.B1(n_9404),
.B2(n_9349),
.Y(n_18817)
);

OR2x6_ASAP7_75t_L g18818 ( 
.A(n_18471),
.B(n_8544),
.Y(n_18818)
);

INVx2_ASAP7_75t_L g18819 ( 
.A(n_18440),
.Y(n_18819)
);

INVx1_ASAP7_75t_L g18820 ( 
.A(n_18418),
.Y(n_18820)
);

INVx1_ASAP7_75t_SL g18821 ( 
.A(n_18139),
.Y(n_18821)
);

INVx2_ASAP7_75t_L g18822 ( 
.A(n_18447),
.Y(n_18822)
);

AND2x2_ASAP7_75t_L g18823 ( 
.A(n_18256),
.B(n_6986),
.Y(n_18823)
);

INVx1_ASAP7_75t_L g18824 ( 
.A(n_18221),
.Y(n_18824)
);

INVx2_ASAP7_75t_L g18825 ( 
.A(n_18429),
.Y(n_18825)
);

INVx2_ASAP7_75t_L g18826 ( 
.A(n_18457),
.Y(n_18826)
);

INVx2_ASAP7_75t_L g18827 ( 
.A(n_18432),
.Y(n_18827)
);

INVxp67_ASAP7_75t_L g18828 ( 
.A(n_18140),
.Y(n_18828)
);

INVx2_ASAP7_75t_L g18829 ( 
.A(n_18443),
.Y(n_18829)
);

AND2x4_ASAP7_75t_L g18830 ( 
.A(n_18465),
.B(n_10545),
.Y(n_18830)
);

INVx1_ASAP7_75t_SL g18831 ( 
.A(n_18359),
.Y(n_18831)
);

AND2x2_ASAP7_75t_L g18832 ( 
.A(n_18280),
.B(n_6986),
.Y(n_18832)
);

INVx1_ASAP7_75t_SL g18833 ( 
.A(n_18365),
.Y(n_18833)
);

INVx1_ASAP7_75t_SL g18834 ( 
.A(n_18367),
.Y(n_18834)
);

INVx2_ASAP7_75t_SL g18835 ( 
.A(n_18335),
.Y(n_18835)
);

INVxp67_ASAP7_75t_SL g18836 ( 
.A(n_18347),
.Y(n_18836)
);

HB1xp67_ASAP7_75t_L g18837 ( 
.A(n_18235),
.Y(n_18837)
);

AOI22xp33_ASAP7_75t_L g18838 ( 
.A1(n_18138),
.A2(n_9507),
.B1(n_9404),
.B2(n_8552),
.Y(n_18838)
);

AND2x2_ASAP7_75t_L g18839 ( 
.A(n_18478),
.B(n_6986),
.Y(n_18839)
);

INVx2_ASAP7_75t_L g18840 ( 
.A(n_18481),
.Y(n_18840)
);

OR2x2_ASAP7_75t_L g18841 ( 
.A(n_18226),
.B(n_18216),
.Y(n_18841)
);

INVx1_ASAP7_75t_L g18842 ( 
.A(n_18419),
.Y(n_18842)
);

NOR2xp33_ASAP7_75t_SL g18843 ( 
.A(n_18413),
.B(n_18258),
.Y(n_18843)
);

INVx2_ASAP7_75t_L g18844 ( 
.A(n_18439),
.Y(n_18844)
);

INVx1_ASAP7_75t_L g18845 ( 
.A(n_18340),
.Y(n_18845)
);

NOR2x1_ASAP7_75t_L g18846 ( 
.A(n_18349),
.B(n_9404),
.Y(n_18846)
);

NAND2xp5_ASAP7_75t_SL g18847 ( 
.A(n_18625),
.B(n_18338),
.Y(n_18847)
);

NAND2xp5_ASAP7_75t_L g18848 ( 
.A(n_18510),
.B(n_18403),
.Y(n_18848)
);

NOR3xp33_ASAP7_75t_L g18849 ( 
.A(n_18511),
.B(n_18384),
.C(n_18334),
.Y(n_18849)
);

AND2x4_ASAP7_75t_SL g18850 ( 
.A(n_18647),
.B(n_18204),
.Y(n_18850)
);

NOR2xp33_ASAP7_75t_L g18851 ( 
.A(n_18528),
.B(n_18603),
.Y(n_18851)
);

INVx1_ASAP7_75t_SL g18852 ( 
.A(n_18571),
.Y(n_18852)
);

AOI211x1_ASAP7_75t_SL g18853 ( 
.A1(n_18654),
.A2(n_18469),
.B(n_18460),
.C(n_18483),
.Y(n_18853)
);

OR2x2_ASAP7_75t_L g18854 ( 
.A(n_18525),
.B(n_18196),
.Y(n_18854)
);

INVx1_ASAP7_75t_L g18855 ( 
.A(n_18552),
.Y(n_18855)
);

AOI22xp5_ASAP7_75t_L g18856 ( 
.A1(n_18548),
.A2(n_18373),
.B1(n_18470),
.B2(n_18475),
.Y(n_18856)
);

AOI21xp33_ASAP7_75t_SL g18857 ( 
.A1(n_18693),
.A2(n_18339),
.B(n_18480),
.Y(n_18857)
);

INVx1_ASAP7_75t_L g18858 ( 
.A(n_18502),
.Y(n_18858)
);

INVx1_ASAP7_75t_SL g18859 ( 
.A(n_18513),
.Y(n_18859)
);

OAI221xp5_ASAP7_75t_SL g18860 ( 
.A1(n_18583),
.A2(n_18430),
.B1(n_18387),
.B2(n_18307),
.C(n_18154),
.Y(n_18860)
);

AND2x2_ASAP7_75t_L g18861 ( 
.A(n_18520),
.B(n_18464),
.Y(n_18861)
);

OAI22xp5_ASAP7_75t_L g18862 ( 
.A1(n_18596),
.A2(n_18145),
.B1(n_18200),
.B2(n_18301),
.Y(n_18862)
);

INVx2_ASAP7_75t_SL g18863 ( 
.A(n_18592),
.Y(n_18863)
);

NAND2x1p5_ASAP7_75t_L g18864 ( 
.A(n_18543),
.B(n_18434),
.Y(n_18864)
);

INVx1_ASAP7_75t_L g18865 ( 
.A(n_18574),
.Y(n_18865)
);

NAND2xp5_ASAP7_75t_L g18866 ( 
.A(n_18509),
.B(n_18133),
.Y(n_18866)
);

NAND3xp33_ASAP7_75t_L g18867 ( 
.A(n_18793),
.B(n_18227),
.C(n_18477),
.Y(n_18867)
);

NOR2xp33_ASAP7_75t_L g18868 ( 
.A(n_18630),
.B(n_18276),
.Y(n_18868)
);

INVx1_ASAP7_75t_L g18869 ( 
.A(n_18514),
.Y(n_18869)
);

NAND2xp5_ASAP7_75t_SL g18870 ( 
.A(n_18791),
.B(n_18491),
.Y(n_18870)
);

A2O1A1Ixp33_ASAP7_75t_L g18871 ( 
.A1(n_18629),
.A2(n_18459),
.B(n_18476),
.C(n_18472),
.Y(n_18871)
);

NAND2xp5_ASAP7_75t_L g18872 ( 
.A(n_18593),
.B(n_18299),
.Y(n_18872)
);

NAND2xp5_ASAP7_75t_L g18873 ( 
.A(n_18703),
.B(n_18479),
.Y(n_18873)
);

INVx1_ASAP7_75t_L g18874 ( 
.A(n_18515),
.Y(n_18874)
);

INVx2_ASAP7_75t_L g18875 ( 
.A(n_18537),
.Y(n_18875)
);

OAI22xp5_ASAP7_75t_L g18876 ( 
.A1(n_18575),
.A2(n_18451),
.B1(n_18494),
.B2(n_18424),
.Y(n_18876)
);

AOI21xp5_ASAP7_75t_L g18877 ( 
.A1(n_18639),
.A2(n_18182),
.B(n_18488),
.Y(n_18877)
);

AOI21xp33_ASAP7_75t_L g18878 ( 
.A1(n_18586),
.A2(n_18623),
.B(n_18516),
.Y(n_18878)
);

OAI22xp33_ASAP7_75t_L g18879 ( 
.A1(n_18707),
.A2(n_18732),
.B1(n_18544),
.B2(n_18519),
.Y(n_18879)
);

INVx2_ASAP7_75t_SL g18880 ( 
.A(n_18688),
.Y(n_18880)
);

NOR2xp33_ASAP7_75t_L g18881 ( 
.A(n_18584),
.B(n_18320),
.Y(n_18881)
);

AOI21x1_ASAP7_75t_L g18882 ( 
.A1(n_18744),
.A2(n_18451),
.B(n_18485),
.Y(n_18882)
);

AOI21xp5_ASAP7_75t_L g18883 ( 
.A1(n_18686),
.A2(n_18231),
.B(n_18191),
.Y(n_18883)
);

NOR3xp33_ASAP7_75t_SL g18884 ( 
.A(n_18705),
.B(n_18489),
.C(n_18490),
.Y(n_18884)
);

INVx1_ASAP7_75t_L g18885 ( 
.A(n_18709),
.Y(n_18885)
);

NAND2xp5_ASAP7_75t_L g18886 ( 
.A(n_18503),
.B(n_18233),
.Y(n_18886)
);

OAI22xp5_ASAP7_75t_L g18887 ( 
.A1(n_18545),
.A2(n_18414),
.B1(n_18248),
.B2(n_18275),
.Y(n_18887)
);

AOI21xp5_ASAP7_75t_L g18888 ( 
.A1(n_18624),
.A2(n_18249),
.B(n_18326),
.Y(n_18888)
);

NAND2x1_ASAP7_75t_L g18889 ( 
.A(n_18564),
.B(n_18482),
.Y(n_18889)
);

AOI21xp33_ASAP7_75t_SL g18890 ( 
.A1(n_18524),
.A2(n_18188),
.B(n_18458),
.Y(n_18890)
);

OAI221xp5_ASAP7_75t_SL g18891 ( 
.A1(n_18546),
.A2(n_18343),
.B1(n_9575),
.B2(n_9504),
.C(n_9497),
.Y(n_18891)
);

AOI221xp5_ASAP7_75t_L g18892 ( 
.A1(n_18837),
.A2(n_9507),
.B1(n_6955),
.B2(n_8128),
.C(n_8168),
.Y(n_18892)
);

NAND2xp5_ASAP7_75t_L g18893 ( 
.A(n_18604),
.B(n_8342),
.Y(n_18893)
);

OAI32xp33_ASAP7_75t_L g18894 ( 
.A1(n_18607),
.A2(n_9349),
.A3(n_9320),
.B1(n_7311),
.B2(n_7127),
.Y(n_18894)
);

AO221x1_ASAP7_75t_L g18895 ( 
.A1(n_18762),
.A2(n_9341),
.B1(n_9473),
.B2(n_9149),
.C(n_8995),
.Y(n_18895)
);

NAND2xp5_ASAP7_75t_L g18896 ( 
.A(n_18612),
.B(n_8344),
.Y(n_18896)
);

AOI211xp5_ASAP7_75t_L g18897 ( 
.A1(n_18632),
.A2(n_8128),
.B(n_8523),
.C(n_8519),
.Y(n_18897)
);

NAND2xp5_ASAP7_75t_L g18898 ( 
.A(n_18673),
.B(n_8344),
.Y(n_18898)
);

O2A1O1Ixp33_ASAP7_75t_L g18899 ( 
.A1(n_18733),
.A2(n_9320),
.B(n_9341),
.C(n_9149),
.Y(n_18899)
);

AOI21xp33_ASAP7_75t_L g18900 ( 
.A1(n_18687),
.A2(n_8168),
.B(n_8165),
.Y(n_18900)
);

NOR3xp33_ASAP7_75t_L g18901 ( 
.A(n_18538),
.B(n_9307),
.C(n_8444),
.Y(n_18901)
);

HB1xp67_ASAP7_75t_L g18902 ( 
.A(n_18664),
.Y(n_18902)
);

INVx1_ASAP7_75t_L g18903 ( 
.A(n_18728),
.Y(n_18903)
);

OR2x2_ASAP7_75t_L g18904 ( 
.A(n_18610),
.B(n_7311),
.Y(n_18904)
);

OAI221xp5_ASAP7_75t_L g18905 ( 
.A1(n_18780),
.A2(n_9575),
.B1(n_9504),
.B2(n_9497),
.C(n_9534),
.Y(n_18905)
);

AOI22xp33_ASAP7_75t_L g18906 ( 
.A1(n_18774),
.A2(n_8165),
.B1(n_8205),
.B2(n_8186),
.Y(n_18906)
);

INVxp67_ASAP7_75t_L g18907 ( 
.A(n_18566),
.Y(n_18907)
);

AOI221xp5_ASAP7_75t_L g18908 ( 
.A1(n_18590),
.A2(n_6955),
.B1(n_8165),
.B2(n_8227),
.C(n_8205),
.Y(n_18908)
);

INVx1_ASAP7_75t_L g18909 ( 
.A(n_18578),
.Y(n_18909)
);

AOI22xp5_ASAP7_75t_L g18910 ( 
.A1(n_18710),
.A2(n_9509),
.B1(n_8205),
.B2(n_8227),
.Y(n_18910)
);

O2A1O1Ixp33_ASAP7_75t_L g18911 ( 
.A1(n_18553),
.A2(n_9341),
.B(n_9473),
.C(n_9149),
.Y(n_18911)
);

AOI22xp5_ASAP7_75t_L g18912 ( 
.A1(n_18738),
.A2(n_9509),
.B1(n_8205),
.B2(n_8227),
.Y(n_18912)
);

INVx1_ASAP7_75t_L g18913 ( 
.A(n_18532),
.Y(n_18913)
);

OAI22xp33_ASAP7_75t_L g18914 ( 
.A1(n_18843),
.A2(n_7311),
.B1(n_7877),
.B2(n_7803),
.Y(n_18914)
);

NAND2xp5_ASAP7_75t_SL g18915 ( 
.A(n_18762),
.B(n_6955),
.Y(n_18915)
);

AO22x1_ASAP7_75t_L g18916 ( 
.A1(n_18569),
.A2(n_7232),
.B1(n_7543),
.B2(n_7355),
.Y(n_18916)
);

NAND2xp5_ASAP7_75t_L g18917 ( 
.A(n_18690),
.B(n_8344),
.Y(n_18917)
);

OAI22xp5_ASAP7_75t_L g18918 ( 
.A1(n_18508),
.A2(n_9028),
.B1(n_9033),
.B2(n_9018),
.Y(n_18918)
);

INVx2_ASAP7_75t_L g18919 ( 
.A(n_18589),
.Y(n_18919)
);

NOR2xp33_ASAP7_75t_L g18920 ( 
.A(n_18717),
.B(n_8165),
.Y(n_18920)
);

AND2x2_ASAP7_75t_L g18921 ( 
.A(n_18562),
.B(n_8098),
.Y(n_18921)
);

INVx1_ASAP7_75t_L g18922 ( 
.A(n_18634),
.Y(n_18922)
);

AOI221xp5_ASAP7_75t_L g18923 ( 
.A1(n_18787),
.A2(n_6955),
.B1(n_8244),
.B2(n_8247),
.C(n_8234),
.Y(n_18923)
);

HB1xp67_ASAP7_75t_L g18924 ( 
.A(n_18771),
.Y(n_18924)
);

AOI211xp5_ASAP7_75t_L g18925 ( 
.A1(n_18768),
.A2(n_18579),
.B(n_18804),
.C(n_18620),
.Y(n_18925)
);

INVx1_ASAP7_75t_L g18926 ( 
.A(n_18637),
.Y(n_18926)
);

INVxp67_ASAP7_75t_L g18927 ( 
.A(n_18638),
.Y(n_18927)
);

CKINVDCx14_ASAP7_75t_R g18928 ( 
.A(n_18527),
.Y(n_18928)
);

INVx2_ASAP7_75t_SL g18929 ( 
.A(n_18567),
.Y(n_18929)
);

AOI221xp5_ASAP7_75t_L g18930 ( 
.A1(n_18559),
.A2(n_18518),
.B1(n_18570),
.B2(n_18572),
.C(n_18667),
.Y(n_18930)
);

AND2x2_ASAP7_75t_L g18931 ( 
.A(n_18800),
.B(n_8098),
.Y(n_18931)
);

INVx1_ASAP7_75t_L g18932 ( 
.A(n_18500),
.Y(n_18932)
);

AOI22xp33_ASAP7_75t_L g18933 ( 
.A1(n_18778),
.A2(n_8234),
.B1(n_8247),
.B2(n_8244),
.Y(n_18933)
);

AOI22xp5_ASAP7_75t_L g18934 ( 
.A1(n_18721),
.A2(n_9509),
.B1(n_8244),
.B2(n_8247),
.Y(n_18934)
);

NOR2xp33_ASAP7_75t_L g18935 ( 
.A(n_18742),
.B(n_8234),
.Y(n_18935)
);

INVx1_ASAP7_75t_L g18936 ( 
.A(n_18839),
.Y(n_18936)
);

HB1xp67_ASAP7_75t_L g18937 ( 
.A(n_18618),
.Y(n_18937)
);

INVx1_ASAP7_75t_L g18938 ( 
.A(n_18651),
.Y(n_18938)
);

INVxp67_ASAP7_75t_L g18939 ( 
.A(n_18668),
.Y(n_18939)
);

INVx1_ASAP7_75t_SL g18940 ( 
.A(n_18745),
.Y(n_18940)
);

OAI21xp5_ASAP7_75t_SL g18941 ( 
.A1(n_18594),
.A2(n_18754),
.B(n_18702),
.Y(n_18941)
);

AND2x2_ASAP7_75t_L g18942 ( 
.A(n_18760),
.B(n_8098),
.Y(n_18942)
);

INVx2_ASAP7_75t_L g18943 ( 
.A(n_18597),
.Y(n_18943)
);

AOI31xp33_ASAP7_75t_L g18944 ( 
.A1(n_18670),
.A2(n_7818),
.A3(n_7806),
.B(n_7578),
.Y(n_18944)
);

AOI32xp33_ASAP7_75t_L g18945 ( 
.A1(n_18615),
.A2(n_8519),
.A3(n_8523),
.B1(n_8274),
.B2(n_8270),
.Y(n_18945)
);

INVx2_ASAP7_75t_L g18946 ( 
.A(n_18823),
.Y(n_18946)
);

OR2x2_ASAP7_75t_L g18947 ( 
.A(n_18749),
.B(n_7867),
.Y(n_18947)
);

OR2x2_ASAP7_75t_L g18948 ( 
.A(n_18558),
.B(n_7867),
.Y(n_18948)
);

INVx1_ASAP7_75t_L g18949 ( 
.A(n_18692),
.Y(n_18949)
);

NAND2xp5_ASAP7_75t_L g18950 ( 
.A(n_18821),
.B(n_8344),
.Y(n_18950)
);

NAND2xp5_ASAP7_75t_L g18951 ( 
.A(n_18801),
.B(n_8347),
.Y(n_18951)
);

AOI22xp5_ASAP7_75t_L g18952 ( 
.A1(n_18775),
.A2(n_9509),
.B1(n_8244),
.B2(n_8247),
.Y(n_18952)
);

OAI21xp33_ASAP7_75t_L g18953 ( 
.A1(n_18790),
.A2(n_8052),
.B(n_8035),
.Y(n_18953)
);

OAI21xp5_ASAP7_75t_L g18954 ( 
.A1(n_18741),
.A2(n_8270),
.B(n_8444),
.Y(n_18954)
);

INVxp67_ASAP7_75t_L g18955 ( 
.A(n_18694),
.Y(n_18955)
);

AOI31xp33_ASAP7_75t_L g18956 ( 
.A1(n_18671),
.A2(n_7818),
.A3(n_7806),
.B(n_7625),
.Y(n_18956)
);

OAI32xp33_ASAP7_75t_L g18957 ( 
.A1(n_18585),
.A2(n_7183),
.A3(n_7187),
.B1(n_7117),
.B2(n_7060),
.Y(n_18957)
);

OR2x2_ASAP7_75t_L g18958 ( 
.A(n_18723),
.B(n_7924),
.Y(n_18958)
);

NAND2xp5_ASAP7_75t_L g18959 ( 
.A(n_18789),
.B(n_8347),
.Y(n_18959)
);

OAI22xp5_ASAP7_75t_L g18960 ( 
.A1(n_18512),
.A2(n_9028),
.B1(n_9033),
.B2(n_9018),
.Y(n_18960)
);

OAI22xp5_ASAP7_75t_L g18961 ( 
.A1(n_18533),
.A2(n_9033),
.B1(n_9038),
.B2(n_9028),
.Y(n_18961)
);

AOI211xp5_ASAP7_75t_L g18962 ( 
.A1(n_18699),
.A2(n_9562),
.B(n_10160),
.C(n_10144),
.Y(n_18962)
);

NAND2xp5_ASAP7_75t_L g18963 ( 
.A(n_18831),
.B(n_8347),
.Y(n_18963)
);

AND2x2_ASAP7_75t_L g18964 ( 
.A(n_18561),
.B(n_8108),
.Y(n_18964)
);

INVx1_ASAP7_75t_L g18965 ( 
.A(n_18695),
.Y(n_18965)
);

INVx2_ASAP7_75t_L g18966 ( 
.A(n_18832),
.Y(n_18966)
);

OAI21xp33_ASAP7_75t_SL g18967 ( 
.A1(n_18672),
.A2(n_10459),
.B(n_10545),
.Y(n_18967)
);

NAND4xp75_ASAP7_75t_SL g18968 ( 
.A(n_18730),
.B(n_8016),
.C(n_8105),
.D(n_7073),
.Y(n_18968)
);

AND2x2_ASAP7_75t_L g18969 ( 
.A(n_18631),
.B(n_8108),
.Y(n_18969)
);

NAND2xp5_ASAP7_75t_L g18970 ( 
.A(n_18833),
.B(n_8347),
.Y(n_18970)
);

INVxp67_ASAP7_75t_L g18971 ( 
.A(n_18675),
.Y(n_18971)
);

INVx1_ASAP7_75t_L g18972 ( 
.A(n_18600),
.Y(n_18972)
);

OR2x2_ASAP7_75t_L g18973 ( 
.A(n_18737),
.B(n_7924),
.Y(n_18973)
);

INVx1_ASAP7_75t_SL g18974 ( 
.A(n_18834),
.Y(n_18974)
);

INVx2_ASAP7_75t_SL g18975 ( 
.A(n_18676),
.Y(n_18975)
);

OAI22xp5_ASAP7_75t_L g18976 ( 
.A1(n_18547),
.A2(n_9045),
.B1(n_9051),
.B2(n_9038),
.Y(n_18976)
);

INVx1_ASAP7_75t_L g18977 ( 
.A(n_18841),
.Y(n_18977)
);

AOI22xp33_ASAP7_75t_L g18978 ( 
.A1(n_18844),
.A2(n_8234),
.B1(n_8289),
.B2(n_8279),
.Y(n_18978)
);

INVx1_ASAP7_75t_L g18979 ( 
.A(n_18836),
.Y(n_18979)
);

AND2x2_ASAP7_75t_SL g18980 ( 
.A(n_18666),
.B(n_9397),
.Y(n_18980)
);

AOI22xp5_ASAP7_75t_L g18981 ( 
.A1(n_18635),
.A2(n_9509),
.B1(n_8289),
.B2(n_8300),
.Y(n_18981)
);

AND2x2_ASAP7_75t_L g18982 ( 
.A(n_18797),
.B(n_18727),
.Y(n_18982)
);

OAI21xp5_ASAP7_75t_L g18983 ( 
.A1(n_18587),
.A2(n_9236),
.B(n_9234),
.Y(n_18983)
);

NOR2xp67_ASAP7_75t_L g18984 ( 
.A(n_18712),
.B(n_7634),
.Y(n_18984)
);

OAI32xp33_ASAP7_75t_L g18985 ( 
.A1(n_18788),
.A2(n_7285),
.A3(n_7342),
.B1(n_7187),
.B2(n_7183),
.Y(n_18985)
);

INVx1_ASAP7_75t_L g18986 ( 
.A(n_18755),
.Y(n_18986)
);

O2A1O1Ixp5_ASAP7_75t_L g18987 ( 
.A1(n_18504),
.A2(n_9045),
.B(n_9051),
.C(n_9038),
.Y(n_18987)
);

NOR2xp33_ASAP7_75t_L g18988 ( 
.A(n_18507),
.B(n_8279),
.Y(n_18988)
);

INVx1_ASAP7_75t_L g18989 ( 
.A(n_18718),
.Y(n_18989)
);

NOR2xp33_ASAP7_75t_L g18990 ( 
.A(n_18822),
.B(n_8279),
.Y(n_18990)
);

AOI21xp33_ASAP7_75t_L g18991 ( 
.A1(n_18616),
.A2(n_18827),
.B(n_18782),
.Y(n_18991)
);

INVx1_ASAP7_75t_L g18992 ( 
.A(n_18521),
.Y(n_18992)
);

AND2x2_ASAP7_75t_L g18993 ( 
.A(n_18802),
.B(n_8108),
.Y(n_18993)
);

OAI22xp33_ASAP7_75t_L g18994 ( 
.A1(n_18697),
.A2(n_7877),
.B1(n_7894),
.B2(n_7803),
.Y(n_18994)
);

INVx1_ASAP7_75t_L g18995 ( 
.A(n_18663),
.Y(n_18995)
);

AND2x4_ASAP7_75t_L g18996 ( 
.A(n_18716),
.B(n_10634),
.Y(n_18996)
);

OAI221xp5_ASAP7_75t_L g18997 ( 
.A1(n_18736),
.A2(n_9534),
.B1(n_9415),
.B2(n_9127),
.C(n_8777),
.Y(n_18997)
);

INVx1_ASAP7_75t_L g18998 ( 
.A(n_18720),
.Y(n_18998)
);

A2O1A1Ixp33_ASAP7_75t_SL g18999 ( 
.A1(n_18653),
.A2(n_7637),
.B(n_7634),
.C(n_9045),
.Y(n_18999)
);

AOI22xp5_ASAP7_75t_L g19000 ( 
.A1(n_18655),
.A2(n_9509),
.B1(n_8289),
.B2(n_8300),
.Y(n_19000)
);

AND2x2_ASAP7_75t_L g19001 ( 
.A(n_18770),
.B(n_8108),
.Y(n_19001)
);

OA211x2_ASAP7_75t_L g19002 ( 
.A1(n_18786),
.A2(n_7637),
.B(n_7620),
.C(n_8724),
.Y(n_19002)
);

OAI22xp33_ASAP7_75t_L g19003 ( 
.A1(n_18816),
.A2(n_7877),
.B1(n_7894),
.B2(n_7803),
.Y(n_19003)
);

OR2x2_ASAP7_75t_L g19004 ( 
.A(n_18811),
.B(n_7941),
.Y(n_19004)
);

AOI211xp5_ASAP7_75t_SL g19005 ( 
.A1(n_18803),
.A2(n_7818),
.B(n_7533),
.C(n_7444),
.Y(n_19005)
);

AOI31xp33_ASAP7_75t_SL g19006 ( 
.A1(n_18828),
.A2(n_7620),
.A3(n_7500),
.B(n_7524),
.Y(n_19006)
);

INVx1_ASAP7_75t_L g19007 ( 
.A(n_18722),
.Y(n_19007)
);

INVx1_ASAP7_75t_L g19008 ( 
.A(n_18758),
.Y(n_19008)
);

OAI22xp33_ASAP7_75t_L g19009 ( 
.A1(n_18819),
.A2(n_7877),
.B1(n_7894),
.B2(n_7803),
.Y(n_19009)
);

NAND2x1_ASAP7_75t_L g19010 ( 
.A(n_18818),
.B(n_9473),
.Y(n_19010)
);

NAND2xp5_ASAP7_75t_L g19011 ( 
.A(n_18743),
.B(n_8352),
.Y(n_19011)
);

NAND2xp5_ASAP7_75t_L g19012 ( 
.A(n_18701),
.B(n_8352),
.Y(n_19012)
);

INVx1_ASAP7_75t_L g19013 ( 
.A(n_18711),
.Y(n_19013)
);

OA33x2_ASAP7_75t_L g19014 ( 
.A1(n_18781),
.A2(n_7620),
.A3(n_7539),
.B1(n_7548),
.B2(n_7538),
.B3(n_7567),
.Y(n_19014)
);

INVx1_ASAP7_75t_L g19015 ( 
.A(n_18506),
.Y(n_19015)
);

AND2x2_ASAP7_75t_L g19016 ( 
.A(n_18636),
.B(n_10634),
.Y(n_19016)
);

AOI22xp5_ASAP7_75t_L g19017 ( 
.A1(n_18725),
.A2(n_8289),
.B1(n_8300),
.B2(n_8279),
.Y(n_19017)
);

INVx1_ASAP7_75t_L g19018 ( 
.A(n_18601),
.Y(n_19018)
);

INVx1_ASAP7_75t_L g19019 ( 
.A(n_18658),
.Y(n_19019)
);

INVx4_ASAP7_75t_L g19020 ( 
.A(n_18706),
.Y(n_19020)
);

INVx1_ASAP7_75t_L g19021 ( 
.A(n_18669),
.Y(n_19021)
);

OAI21xp5_ASAP7_75t_L g19022 ( 
.A1(n_18764),
.A2(n_9236),
.B(n_9234),
.Y(n_19022)
);

NAND2xp5_ASAP7_75t_L g19023 ( 
.A(n_18650),
.B(n_8352),
.Y(n_19023)
);

NOR2xp33_ASAP7_75t_L g19024 ( 
.A(n_18759),
.B(n_8300),
.Y(n_19024)
);

NAND2xp5_ASAP7_75t_L g19025 ( 
.A(n_18835),
.B(n_8352),
.Y(n_19025)
);

AOI21xp5_ASAP7_75t_L g19026 ( 
.A1(n_18501),
.A2(n_9078),
.B(n_9051),
.Y(n_19026)
);

OAI22xp5_ASAP7_75t_L g19027 ( 
.A1(n_18708),
.A2(n_18565),
.B1(n_18700),
.B2(n_18644),
.Y(n_19027)
);

INVx1_ASAP7_75t_L g19028 ( 
.A(n_18677),
.Y(n_19028)
);

AOI221xp5_ASAP7_75t_L g19029 ( 
.A1(n_18642),
.A2(n_6955),
.B1(n_8328),
.B2(n_9553),
.C(n_8380),
.Y(n_19029)
);

INVxp67_ASAP7_75t_L g19030 ( 
.A(n_18761),
.Y(n_19030)
);

AND2x2_ASAP7_75t_L g19031 ( 
.A(n_18731),
.B(n_6986),
.Y(n_19031)
);

INVxp67_ASAP7_75t_L g19032 ( 
.A(n_18724),
.Y(n_19032)
);

NAND3xp33_ASAP7_75t_L g19033 ( 
.A(n_18599),
.B(n_18729),
.C(n_18726),
.Y(n_19033)
);

A2O1A1Ixp33_ASAP7_75t_L g19034 ( 
.A1(n_18554),
.A2(n_8178),
.B(n_8136),
.C(n_8132),
.Y(n_19034)
);

INVx2_ASAP7_75t_L g19035 ( 
.A(n_18535),
.Y(n_19035)
);

NAND2xp33_ASAP7_75t_SL g19036 ( 
.A(n_18577),
.B(n_7232),
.Y(n_19036)
);

AOI22xp5_ASAP7_75t_L g19037 ( 
.A1(n_18808),
.A2(n_8328),
.B1(n_8380),
.B2(n_8367),
.Y(n_19037)
);

OAI22xp5_ASAP7_75t_L g19038 ( 
.A1(n_18659),
.A2(n_9078),
.B1(n_9083),
.B2(n_9080),
.Y(n_19038)
);

OAI221xp5_ASAP7_75t_L g19039 ( 
.A1(n_18580),
.A2(n_8777),
.B1(n_9477),
.B2(n_9454),
.C(n_9340),
.Y(n_19039)
);

NAND2xp5_ASAP7_75t_SL g19040 ( 
.A(n_18825),
.B(n_6955),
.Y(n_19040)
);

XOR2xp5_ASAP7_75t_L g19041 ( 
.A(n_18685),
.B(n_8172),
.Y(n_19041)
);

INVx1_ASAP7_75t_L g19042 ( 
.A(n_18679),
.Y(n_19042)
);

NOR2xp67_ASAP7_75t_L g19043 ( 
.A(n_18794),
.B(n_7941),
.Y(n_19043)
);

AOI22xp5_ASAP7_75t_L g19044 ( 
.A1(n_18698),
.A2(n_8328),
.B1(n_8380),
.B2(n_8367),
.Y(n_19044)
);

NAND2xp5_ASAP7_75t_L g19045 ( 
.A(n_18748),
.B(n_8367),
.Y(n_19045)
);

AO21x1_ASAP7_75t_L g19046 ( 
.A1(n_18752),
.A2(n_7625),
.B(n_7533),
.Y(n_19046)
);

INVx1_ASAP7_75t_L g19047 ( 
.A(n_18680),
.Y(n_19047)
);

NAND2xp5_ASAP7_75t_L g19048 ( 
.A(n_18767),
.B(n_8367),
.Y(n_19048)
);

OAI31xp33_ASAP7_75t_L g19049 ( 
.A1(n_18769),
.A2(n_18531),
.A3(n_18523),
.B(n_18598),
.Y(n_19049)
);

OAI22xp5_ASAP7_75t_L g19050 ( 
.A1(n_18829),
.A2(n_9078),
.B1(n_9083),
.B2(n_9080),
.Y(n_19050)
);

INVx1_ASAP7_75t_L g19051 ( 
.A(n_18619),
.Y(n_19051)
);

NAND2x1_ASAP7_75t_L g19052 ( 
.A(n_18818),
.B(n_9490),
.Y(n_19052)
);

INVx1_ASAP7_75t_L g19053 ( 
.A(n_18626),
.Y(n_19053)
);

O2A1O1Ixp33_ASAP7_75t_SL g19054 ( 
.A1(n_18591),
.A2(n_7945),
.B(n_8032),
.C(n_7992),
.Y(n_19054)
);

AND2x2_ASAP7_75t_L g19055 ( 
.A(n_18734),
.B(n_6995),
.Y(n_19055)
);

INVx1_ASAP7_75t_L g19056 ( 
.A(n_18517),
.Y(n_19056)
);

INVx1_ASAP7_75t_L g19057 ( 
.A(n_18582),
.Y(n_19057)
);

OAI22xp5_ASAP7_75t_L g19058 ( 
.A1(n_18840),
.A2(n_9080),
.B1(n_9084),
.B2(n_9083),
.Y(n_19058)
);

O2A1O1Ixp33_ASAP7_75t_L g19059 ( 
.A1(n_18826),
.A2(n_9537),
.B(n_9490),
.C(n_9562),
.Y(n_19059)
);

NAND2xp5_ASAP7_75t_L g19060 ( 
.A(n_18845),
.B(n_8380),
.Y(n_19060)
);

INVx1_ASAP7_75t_L g19061 ( 
.A(n_18646),
.Y(n_19061)
);

NAND3x1_ASAP7_75t_L g19062 ( 
.A(n_18824),
.B(n_9086),
.C(n_9084),
.Y(n_19062)
);

INVxp67_ASAP7_75t_L g19063 ( 
.A(n_18812),
.Y(n_19063)
);

NAND3xp33_ASAP7_75t_L g19064 ( 
.A(n_18799),
.B(n_8328),
.C(n_8402),
.Y(n_19064)
);

AOI22xp33_ASAP7_75t_SL g19065 ( 
.A1(n_18540),
.A2(n_9361),
.B1(n_9511),
.B2(n_9193),
.Y(n_19065)
);

NOR2xp33_ASAP7_75t_L g19066 ( 
.A(n_18796),
.B(n_18806),
.Y(n_19066)
);

INVx2_ASAP7_75t_L g19067 ( 
.A(n_18535),
.Y(n_19067)
);

NAND3xp33_ASAP7_75t_L g19068 ( 
.A(n_18809),
.B(n_8409),
.C(n_8402),
.Y(n_19068)
);

OAI221xp5_ASAP7_75t_L g19069 ( 
.A1(n_18581),
.A2(n_9477),
.B1(n_9454),
.B2(n_9293),
.C(n_8330),
.Y(n_19069)
);

AOI21xp5_ASAP7_75t_SL g19070 ( 
.A1(n_18740),
.A2(n_7877),
.B(n_7803),
.Y(n_19070)
);

OR2x2_ASAP7_75t_L g19071 ( 
.A(n_18628),
.B(n_7945),
.Y(n_19071)
);

AND2x2_ASAP7_75t_L g19072 ( 
.A(n_18751),
.B(n_6995),
.Y(n_19072)
);

OAI21xp33_ASAP7_75t_SL g19073 ( 
.A1(n_18753),
.A2(n_8739),
.B(n_8736),
.Y(n_19073)
);

INVx1_ASAP7_75t_L g19074 ( 
.A(n_18602),
.Y(n_19074)
);

INVx1_ASAP7_75t_L g19075 ( 
.A(n_18814),
.Y(n_19075)
);

INVx1_ASAP7_75t_L g19076 ( 
.A(n_18820),
.Y(n_19076)
);

AOI21xp5_ASAP7_75t_L g19077 ( 
.A1(n_18505),
.A2(n_9086),
.B(n_9084),
.Y(n_19077)
);

OAI21xp33_ASAP7_75t_L g19078 ( 
.A1(n_18805),
.A2(n_8052),
.B(n_7539),
.Y(n_19078)
);

INVx1_ASAP7_75t_L g19079 ( 
.A(n_18842),
.Y(n_19079)
);

NAND2xp5_ASAP7_75t_L g19080 ( 
.A(n_18779),
.B(n_8402),
.Y(n_19080)
);

AOI32xp33_ASAP7_75t_L g19081 ( 
.A1(n_18539),
.A2(n_18798),
.A3(n_18772),
.B1(n_18773),
.B2(n_18784),
.Y(n_19081)
);

INVx2_ASAP7_75t_L g19082 ( 
.A(n_18621),
.Y(n_19082)
);

INVxp67_ASAP7_75t_SL g19083 ( 
.A(n_18648),
.Y(n_19083)
);

NAND2xp5_ASAP7_75t_L g19084 ( 
.A(n_18573),
.B(n_8402),
.Y(n_19084)
);

OAI22xp33_ASAP7_75t_L g19085 ( 
.A1(n_18757),
.A2(n_18529),
.B1(n_18551),
.B2(n_18549),
.Y(n_19085)
);

OR2x2_ASAP7_75t_L g19086 ( 
.A(n_18756),
.B(n_7992),
.Y(n_19086)
);

OAI21xp5_ASAP7_75t_L g19087 ( 
.A1(n_18750),
.A2(n_9236),
.B(n_9234),
.Y(n_19087)
);

INVx1_ASAP7_75t_L g19088 ( 
.A(n_18684),
.Y(n_19088)
);

OAI221xp5_ASAP7_75t_L g19089 ( 
.A1(n_18622),
.A2(n_8330),
.B1(n_8357),
.B2(n_8197),
.C(n_8172),
.Y(n_19089)
);

INVx1_ASAP7_75t_SL g19090 ( 
.A(n_18608),
.Y(n_19090)
);

NOR3xp33_ASAP7_75t_L g19091 ( 
.A(n_18627),
.B(n_8708),
.C(n_8513),
.Y(n_19091)
);

INVx1_ASAP7_75t_L g19092 ( 
.A(n_18714),
.Y(n_19092)
);

NAND3xp33_ASAP7_75t_SL g19093 ( 
.A(n_18609),
.B(n_8197),
.C(n_8172),
.Y(n_19093)
);

O2A1O1Ixp5_ASAP7_75t_L g19094 ( 
.A1(n_18652),
.A2(n_9092),
.B(n_9094),
.C(n_9086),
.Y(n_19094)
);

OAI21xp5_ASAP7_75t_L g19095 ( 
.A1(n_18645),
.A2(n_8513),
.B(n_8429),
.Y(n_19095)
);

INVx1_ASAP7_75t_L g19096 ( 
.A(n_18715),
.Y(n_19096)
);

NOR2xp33_ASAP7_75t_L g19097 ( 
.A(n_18807),
.B(n_8409),
.Y(n_19097)
);

INVx1_ASAP7_75t_L g19098 ( 
.A(n_18739),
.Y(n_19098)
);

INVx1_ASAP7_75t_SL g19099 ( 
.A(n_18526),
.Y(n_19099)
);

OAI22xp5_ASAP7_75t_L g19100 ( 
.A1(n_18838),
.A2(n_9092),
.B1(n_9101),
.B2(n_9094),
.Y(n_19100)
);

INVxp67_ASAP7_75t_L g19101 ( 
.A(n_18704),
.Y(n_19101)
);

NOR2xp33_ASAP7_75t_L g19102 ( 
.A(n_18763),
.B(n_8409),
.Y(n_19102)
);

NAND2xp5_ASAP7_75t_L g19103 ( 
.A(n_18785),
.B(n_8409),
.Y(n_19103)
);

AOI222xp33_ASAP7_75t_L g19104 ( 
.A1(n_18719),
.A2(n_8212),
.B1(n_8421),
.B2(n_8425),
.C1(n_8420),
.C2(n_8414),
.Y(n_19104)
);

INVx1_ASAP7_75t_L g19105 ( 
.A(n_18815),
.Y(n_19105)
);

INVx2_ASAP7_75t_L g19106 ( 
.A(n_18536),
.Y(n_19106)
);

INVxp67_ASAP7_75t_L g19107 ( 
.A(n_18713),
.Y(n_19107)
);

INVx1_ASAP7_75t_L g19108 ( 
.A(n_18810),
.Y(n_19108)
);

NAND2xp5_ASAP7_75t_L g19109 ( 
.A(n_18563),
.B(n_8414),
.Y(n_19109)
);

AND2x2_ASAP7_75t_L g19110 ( 
.A(n_18766),
.B(n_6995),
.Y(n_19110)
);

NAND2xp5_ASAP7_75t_L g19111 ( 
.A(n_18556),
.B(n_8414),
.Y(n_19111)
);

INVx1_ASAP7_75t_L g19112 ( 
.A(n_18777),
.Y(n_19112)
);

NOR4xp25_ASAP7_75t_SL g19113 ( 
.A(n_18683),
.B(n_8028),
.C(n_8045),
.D(n_8025),
.Y(n_19113)
);

NAND2xp5_ASAP7_75t_SL g19114 ( 
.A(n_18830),
.B(n_18633),
.Y(n_19114)
);

OAI22xp33_ASAP7_75t_SL g19115 ( 
.A1(n_18696),
.A2(n_8197),
.B1(n_8330),
.B2(n_8172),
.Y(n_19115)
);

AND2x2_ASAP7_75t_L g19116 ( 
.A(n_18783),
.B(n_6995),
.Y(n_19116)
);

NAND2xp5_ASAP7_75t_L g19117 ( 
.A(n_18522),
.B(n_8414),
.Y(n_19117)
);

INVx1_ASAP7_75t_L g19118 ( 
.A(n_18792),
.Y(n_19118)
);

INVx1_ASAP7_75t_L g19119 ( 
.A(n_18681),
.Y(n_19119)
);

INVx1_ASAP7_75t_L g19120 ( 
.A(n_18846),
.Y(n_19120)
);

OAI21xp33_ASAP7_75t_L g19121 ( 
.A1(n_18683),
.A2(n_7539),
.B(n_7538),
.Y(n_19121)
);

OAI22xp33_ASAP7_75t_L g19122 ( 
.A1(n_18641),
.A2(n_8056),
.B1(n_8057),
.B2(n_7894),
.Y(n_19122)
);

AND2x2_ASAP7_75t_L g19123 ( 
.A(n_18813),
.B(n_8694),
.Y(n_19123)
);

NAND2xp5_ASAP7_75t_L g19124 ( 
.A(n_18747),
.B(n_8420),
.Y(n_19124)
);

INVx1_ASAP7_75t_L g19125 ( 
.A(n_18674),
.Y(n_19125)
);

OAI22xp5_ASAP7_75t_L g19126 ( 
.A1(n_18588),
.A2(n_18746),
.B1(n_18542),
.B2(n_18530),
.Y(n_19126)
);

OAI21xp33_ASAP7_75t_L g19127 ( 
.A1(n_18640),
.A2(n_7548),
.B(n_7538),
.Y(n_19127)
);

NOR2xp33_ASAP7_75t_L g19128 ( 
.A(n_18691),
.B(n_8420),
.Y(n_19128)
);

INVx2_ASAP7_75t_SL g19129 ( 
.A(n_18657),
.Y(n_19129)
);

INVx1_ASAP7_75t_L g19130 ( 
.A(n_18678),
.Y(n_19130)
);

INVx1_ASAP7_75t_L g19131 ( 
.A(n_18660),
.Y(n_19131)
);

INVxp67_ASAP7_75t_L g19132 ( 
.A(n_18662),
.Y(n_19132)
);

OAI22xp33_ASAP7_75t_L g19133 ( 
.A1(n_18568),
.A2(n_18776),
.B1(n_18576),
.B2(n_18605),
.Y(n_19133)
);

INVx1_ASAP7_75t_L g19134 ( 
.A(n_18614),
.Y(n_19134)
);

INVx1_ASAP7_75t_L g19135 ( 
.A(n_18595),
.Y(n_19135)
);

AOI22xp33_ASAP7_75t_L g19136 ( 
.A1(n_18649),
.A2(n_8550),
.B1(n_8552),
.B2(n_8914),
.Y(n_19136)
);

INVx1_ASAP7_75t_L g19137 ( 
.A(n_18606),
.Y(n_19137)
);

INVx1_ASAP7_75t_L g19138 ( 
.A(n_18611),
.Y(n_19138)
);

NOR2xp33_ASAP7_75t_L g19139 ( 
.A(n_18613),
.B(n_8420),
.Y(n_19139)
);

INVxp67_ASAP7_75t_L g19140 ( 
.A(n_18617),
.Y(n_19140)
);

A2O1A1Ixp33_ASAP7_75t_L g19141 ( 
.A1(n_18643),
.A2(n_8136),
.B(n_8132),
.C(n_8277),
.Y(n_19141)
);

INVxp67_ASAP7_75t_L g19142 ( 
.A(n_18557),
.Y(n_19142)
);

AOI322xp5_ASAP7_75t_L g19143 ( 
.A1(n_18879),
.A2(n_18656),
.A3(n_18550),
.B1(n_18541),
.B2(n_18689),
.C1(n_18682),
.C2(n_18560),
.Y(n_19143)
);

INVx2_ASAP7_75t_SL g19144 ( 
.A(n_18902),
.Y(n_19144)
);

INVx1_ASAP7_75t_SL g19145 ( 
.A(n_18852),
.Y(n_19145)
);

INVxp67_ASAP7_75t_L g19146 ( 
.A(n_18924),
.Y(n_19146)
);

OR2x2_ASAP7_75t_L g19147 ( 
.A(n_18885),
.B(n_18555),
.Y(n_19147)
);

NAND3xp33_ASAP7_75t_L g19148 ( 
.A(n_18925),
.B(n_18735),
.C(n_18795),
.Y(n_19148)
);

AOI22xp5_ASAP7_75t_L g19149 ( 
.A1(n_19099),
.A2(n_18661),
.B1(n_18665),
.B2(n_18765),
.Y(n_19149)
);

INVx1_ASAP7_75t_L g19150 ( 
.A(n_19083),
.Y(n_19150)
);

AND2x2_ASAP7_75t_L g19151 ( 
.A(n_18907),
.B(n_18534),
.Y(n_19151)
);

OAI322xp33_ASAP7_75t_L g19152 ( 
.A1(n_18928),
.A2(n_18817),
.A3(n_9101),
.B1(n_9107),
.B2(n_9092),
.C1(n_9114),
.C2(n_9112),
.Y(n_19152)
);

AOI221xp5_ASAP7_75t_L g19153 ( 
.A1(n_18878),
.A2(n_6955),
.B1(n_8425),
.B2(n_8433),
.C(n_8421),
.Y(n_19153)
);

INVx1_ASAP7_75t_L g19154 ( 
.A(n_18903),
.Y(n_19154)
);

OAI21xp33_ASAP7_75t_SL g19155 ( 
.A1(n_18940),
.A2(n_8739),
.B(n_8736),
.Y(n_19155)
);

OAI22xp5_ASAP7_75t_L g19156 ( 
.A1(n_18855),
.A2(n_18865),
.B1(n_18858),
.B2(n_18955),
.Y(n_19156)
);

INVx1_ASAP7_75t_L g19157 ( 
.A(n_18937),
.Y(n_19157)
);

A2O1A1Ixp33_ASAP7_75t_L g19158 ( 
.A1(n_18868),
.A2(n_8515),
.B(n_8136),
.C(n_8132),
.Y(n_19158)
);

NAND2xp5_ASAP7_75t_L g19159 ( 
.A(n_18859),
.B(n_8421),
.Y(n_19159)
);

AOI22xp5_ASAP7_75t_L g19160 ( 
.A1(n_19140),
.A2(n_8425),
.B1(n_8433),
.B2(n_8421),
.Y(n_19160)
);

AND2x2_ASAP7_75t_L g19161 ( 
.A(n_18982),
.B(n_8694),
.Y(n_19161)
);

INVx1_ASAP7_75t_L g19162 ( 
.A(n_18875),
.Y(n_19162)
);

AND2x2_ASAP7_75t_L g19163 ( 
.A(n_18969),
.B(n_8694),
.Y(n_19163)
);

INVx1_ASAP7_75t_L g19164 ( 
.A(n_18851),
.Y(n_19164)
);

INVx1_ASAP7_75t_L g19165 ( 
.A(n_18854),
.Y(n_19165)
);

INVx1_ASAP7_75t_L g19166 ( 
.A(n_18975),
.Y(n_19166)
);

OAI22xp5_ASAP7_75t_L g19167 ( 
.A1(n_18939),
.A2(n_9094),
.B1(n_9107),
.B2(n_9101),
.Y(n_19167)
);

OAI221xp5_ASAP7_75t_L g19168 ( 
.A1(n_18884),
.A2(n_8330),
.B1(n_8357),
.B2(n_8197),
.C(n_8172),
.Y(n_19168)
);

INVx1_ASAP7_75t_L g19169 ( 
.A(n_19008),
.Y(n_19169)
);

AOI211x1_ASAP7_75t_L g19170 ( 
.A1(n_18882),
.A2(n_9553),
.B(n_7548),
.C(n_9112),
.Y(n_19170)
);

AOI22xp33_ASAP7_75t_L g19171 ( 
.A1(n_19129),
.A2(n_8552),
.B1(n_8550),
.B2(n_8914),
.Y(n_19171)
);

AOI22xp5_ASAP7_75t_L g19172 ( 
.A1(n_19142),
.A2(n_8433),
.B1(n_8440),
.B2(n_8425),
.Y(n_19172)
);

NAND2xp5_ASAP7_75t_L g19173 ( 
.A(n_18974),
.B(n_8433),
.Y(n_19173)
);

AOI22xp33_ASAP7_75t_L g19174 ( 
.A1(n_19135),
.A2(n_8550),
.B1(n_8916),
.B2(n_8914),
.Y(n_19174)
);

INVx1_ASAP7_75t_L g19175 ( 
.A(n_18909),
.Y(n_19175)
);

OAI21xp33_ASAP7_75t_L g19176 ( 
.A1(n_18881),
.A2(n_7734),
.B(n_7727),
.Y(n_19176)
);

INVx1_ASAP7_75t_SL g19177 ( 
.A(n_18848),
.Y(n_19177)
);

OAI22xp5_ASAP7_75t_L g19178 ( 
.A1(n_18949),
.A2(n_9107),
.B1(n_9114),
.B2(n_9112),
.Y(n_19178)
);

INVx1_ASAP7_75t_L g19179 ( 
.A(n_18919),
.Y(n_19179)
);

OAI32xp33_ASAP7_75t_L g19180 ( 
.A1(n_18853),
.A2(n_7285),
.A3(n_7369),
.B1(n_7342),
.B2(n_7187),
.Y(n_19180)
);

INVx2_ASAP7_75t_L g19181 ( 
.A(n_19020),
.Y(n_19181)
);

NAND3xp33_ASAP7_75t_L g19182 ( 
.A(n_18857),
.B(n_8457),
.C(n_8440),
.Y(n_19182)
);

OAI322xp33_ASAP7_75t_L g19183 ( 
.A1(n_19132),
.A2(n_9129),
.A3(n_9119),
.B1(n_9153),
.B2(n_9157),
.C1(n_9122),
.C2(n_9114),
.Y(n_19183)
);

INVx1_ASAP7_75t_L g19184 ( 
.A(n_18863),
.Y(n_19184)
);

OR2x2_ASAP7_75t_L g19185 ( 
.A(n_19020),
.B(n_8032),
.Y(n_19185)
);

INVxp67_ASAP7_75t_L g19186 ( 
.A(n_18847),
.Y(n_19186)
);

OAI222xp33_ASAP7_75t_L g19187 ( 
.A1(n_18927),
.A2(n_9103),
.B1(n_9032),
.B2(n_9126),
.C1(n_9064),
.C2(n_9001),
.Y(n_19187)
);

O2A1O1Ixp33_ASAP7_75t_L g19188 ( 
.A1(n_18880),
.A2(n_9537),
.B(n_9490),
.C(n_7720),
.Y(n_19188)
);

INVx1_ASAP7_75t_L g19189 ( 
.A(n_18922),
.Y(n_19189)
);

INVx1_ASAP7_75t_L g19190 ( 
.A(n_18926),
.Y(n_19190)
);

INVx2_ASAP7_75t_L g19191 ( 
.A(n_18977),
.Y(n_19191)
);

INVx1_ASAP7_75t_L g19192 ( 
.A(n_18913),
.Y(n_19192)
);

OAI22xp5_ASAP7_75t_L g19193 ( 
.A1(n_18965),
.A2(n_19033),
.B1(n_18938),
.B2(n_18867),
.Y(n_19193)
);

AND2x2_ASAP7_75t_SL g19194 ( 
.A(n_18849),
.B(n_9238),
.Y(n_19194)
);

NAND3xp33_ASAP7_75t_L g19195 ( 
.A(n_18971),
.B(n_8457),
.C(n_8440),
.Y(n_19195)
);

INVx1_ASAP7_75t_SL g19196 ( 
.A(n_18873),
.Y(n_19196)
);

OAI21xp33_ASAP7_75t_L g19197 ( 
.A1(n_18869),
.A2(n_7734),
.B(n_7727),
.Y(n_19197)
);

OAI21xp33_ASAP7_75t_L g19198 ( 
.A1(n_18874),
.A2(n_7734),
.B(n_7727),
.Y(n_19198)
);

NAND2xp5_ASAP7_75t_L g19199 ( 
.A(n_18980),
.B(n_8440),
.Y(n_19199)
);

BUFx2_ASAP7_75t_L g19200 ( 
.A(n_18864),
.Y(n_19200)
);

AOI22xp5_ASAP7_75t_SL g19201 ( 
.A1(n_19030),
.A2(n_19032),
.B1(n_18872),
.B2(n_19063),
.Y(n_19201)
);

INVx1_ASAP7_75t_L g19202 ( 
.A(n_18946),
.Y(n_19202)
);

NOR2xp33_ASAP7_75t_SL g19203 ( 
.A(n_18991),
.B(n_7232),
.Y(n_19203)
);

INVx1_ASAP7_75t_L g19204 ( 
.A(n_18966),
.Y(n_19204)
);

OAI32xp33_ASAP7_75t_L g19205 ( 
.A1(n_18866),
.A2(n_7342),
.A3(n_7369),
.B1(n_7285),
.B2(n_7894),
.Y(n_19205)
);

A2O1A1Ixp33_ASAP7_75t_L g19206 ( 
.A1(n_18972),
.A2(n_8515),
.B(n_8513),
.C(n_8212),
.Y(n_19206)
);

NAND2xp33_ASAP7_75t_L g19207 ( 
.A(n_18932),
.B(n_7355),
.Y(n_19207)
);

OAI22xp33_ASAP7_75t_L g19208 ( 
.A1(n_18856),
.A2(n_8057),
.B1(n_8076),
.B2(n_8056),
.Y(n_19208)
);

NAND2xp5_ASAP7_75t_L g19209 ( 
.A(n_18942),
.B(n_8457),
.Y(n_19209)
);

AOI22xp5_ASAP7_75t_L g19210 ( 
.A1(n_19137),
.A2(n_8458),
.B1(n_8459),
.B2(n_8457),
.Y(n_19210)
);

OAI22xp5_ASAP7_75t_L g19211 ( 
.A1(n_18979),
.A2(n_9119),
.B1(n_9129),
.B2(n_9122),
.Y(n_19211)
);

INVx1_ASAP7_75t_SL g19212 ( 
.A(n_18861),
.Y(n_19212)
);

OR2x2_ASAP7_75t_L g19213 ( 
.A(n_18936),
.B(n_8040),
.Y(n_19213)
);

INVx1_ASAP7_75t_L g19214 ( 
.A(n_19013),
.Y(n_19214)
);

INVx2_ASAP7_75t_L g19215 ( 
.A(n_18964),
.Y(n_19215)
);

OAI22xp5_ASAP7_75t_L g19216 ( 
.A1(n_18989),
.A2(n_9119),
.B1(n_9129),
.B2(n_9122),
.Y(n_19216)
);

AND2x2_ASAP7_75t_L g19217 ( 
.A(n_18921),
.B(n_18993),
.Y(n_19217)
);

NOR3xp33_ASAP7_75t_L g19218 ( 
.A(n_18941),
.B(n_8515),
.C(n_8708),
.Y(n_19218)
);

AOI21xp33_ASAP7_75t_L g19219 ( 
.A1(n_19090),
.A2(n_8916),
.B(n_8914),
.Y(n_19219)
);

OAI21xp33_ASAP7_75t_L g19220 ( 
.A1(n_18986),
.A2(n_7762),
.B(n_7755),
.Y(n_19220)
);

NAND2xp5_ASAP7_75t_L g19221 ( 
.A(n_18992),
.B(n_19043),
.Y(n_19221)
);

AOI221xp5_ASAP7_75t_L g19222 ( 
.A1(n_18994),
.A2(n_6955),
.B1(n_8459),
.B2(n_8497),
.C(n_8458),
.Y(n_19222)
);

NOR2x1_ASAP7_75t_L g19223 ( 
.A(n_18870),
.B(n_18995),
.Y(n_19223)
);

INVx2_ASAP7_75t_L g19224 ( 
.A(n_19061),
.Y(n_19224)
);

HB1xp67_ASAP7_75t_L g19225 ( 
.A(n_18984),
.Y(n_19225)
);

AOI211xp5_ASAP7_75t_L g19226 ( 
.A1(n_19027),
.A2(n_8655),
.B(n_8650),
.C(n_7355),
.Y(n_19226)
);

NAND2xp5_ASAP7_75t_L g19227 ( 
.A(n_19074),
.B(n_8458),
.Y(n_19227)
);

NAND2xp5_ASAP7_75t_L g19228 ( 
.A(n_19018),
.B(n_8458),
.Y(n_19228)
);

AOI222xp33_ASAP7_75t_L g19229 ( 
.A1(n_18967),
.A2(n_8212),
.B1(n_8508),
.B2(n_8531),
.C1(n_8497),
.C2(n_8459),
.Y(n_19229)
);

INVx1_ASAP7_75t_SL g19230 ( 
.A(n_18850),
.Y(n_19230)
);

AOI22xp33_ASAP7_75t_L g19231 ( 
.A1(n_19138),
.A2(n_8916),
.B1(n_8914),
.B2(n_8459),
.Y(n_19231)
);

AOI21xp33_ASAP7_75t_L g19232 ( 
.A1(n_19131),
.A2(n_8916),
.B(n_8729),
.Y(n_19232)
);

A2O1A1Ixp33_ASAP7_75t_L g19233 ( 
.A1(n_19049),
.A2(n_8277),
.B(n_8220),
.C(n_8237),
.Y(n_19233)
);

OAI21xp5_ASAP7_75t_L g19234 ( 
.A1(n_18877),
.A2(n_8277),
.B(n_8429),
.Y(n_19234)
);

AOI21xp33_ASAP7_75t_L g19235 ( 
.A1(n_18929),
.A2(n_8916),
.B(n_8729),
.Y(n_19235)
);

INVx1_ASAP7_75t_L g19236 ( 
.A(n_18998),
.Y(n_19236)
);

INVx2_ASAP7_75t_L g19237 ( 
.A(n_19057),
.Y(n_19237)
);

INVx1_ASAP7_75t_SL g19238 ( 
.A(n_19007),
.Y(n_19238)
);

NAND3xp33_ASAP7_75t_L g19239 ( 
.A(n_19081),
.B(n_8508),
.C(n_8497),
.Y(n_19239)
);

NAND2xp5_ASAP7_75t_L g19240 ( 
.A(n_19019),
.B(n_8497),
.Y(n_19240)
);

INVx1_ASAP7_75t_L g19241 ( 
.A(n_19062),
.Y(n_19241)
);

NAND2xp5_ASAP7_75t_L g19242 ( 
.A(n_19021),
.B(n_8508),
.Y(n_19242)
);

AND2x2_ASAP7_75t_L g19243 ( 
.A(n_18931),
.B(n_8694),
.Y(n_19243)
);

OR2x2_ASAP7_75t_L g19244 ( 
.A(n_18893),
.B(n_8040),
.Y(n_19244)
);

INVx1_ASAP7_75t_L g19245 ( 
.A(n_19028),
.Y(n_19245)
);

AOI22xp33_ASAP7_75t_L g19246 ( 
.A1(n_19139),
.A2(n_8508),
.B1(n_8546),
.B2(n_8531),
.Y(n_19246)
);

INVx2_ASAP7_75t_L g19247 ( 
.A(n_19042),
.Y(n_19247)
);

INVx1_ASAP7_75t_L g19248 ( 
.A(n_19047),
.Y(n_19248)
);

O2A1O1Ixp5_ASAP7_75t_L g19249 ( 
.A1(n_18889),
.A2(n_9157),
.B(n_9158),
.C(n_9153),
.Y(n_19249)
);

INVx2_ASAP7_75t_SL g19250 ( 
.A(n_18948),
.Y(n_19250)
);

NOR2xp33_ASAP7_75t_SL g19251 ( 
.A(n_19015),
.B(n_7355),
.Y(n_19251)
);

INVx1_ASAP7_75t_L g19252 ( 
.A(n_19051),
.Y(n_19252)
);

AND2x2_ASAP7_75t_L g19253 ( 
.A(n_19076),
.B(n_8694),
.Y(n_19253)
);

INVx1_ASAP7_75t_L g19254 ( 
.A(n_19053),
.Y(n_19254)
);

OAI21xp33_ASAP7_75t_L g19255 ( 
.A1(n_19066),
.A2(n_7762),
.B(n_7755),
.Y(n_19255)
);

A2O1A1Ixp33_ASAP7_75t_L g19256 ( 
.A1(n_18920),
.A2(n_8220),
.B(n_8237),
.C(n_8650),
.Y(n_19256)
);

INVx1_ASAP7_75t_L g19257 ( 
.A(n_19056),
.Y(n_19257)
);

AND2x2_ASAP7_75t_L g19258 ( 
.A(n_19079),
.B(n_8694),
.Y(n_19258)
);

NAND2xp5_ASAP7_75t_L g19259 ( 
.A(n_19088),
.B(n_8531),
.Y(n_19259)
);

OAI21xp5_ASAP7_75t_L g19260 ( 
.A1(n_18935),
.A2(n_8429),
.B(n_8220),
.Y(n_19260)
);

AND4x1_ASAP7_75t_L g19261 ( 
.A(n_18930),
.B(n_8924),
.C(n_8724),
.D(n_7520),
.Y(n_19261)
);

NAND2xp5_ASAP7_75t_L g19262 ( 
.A(n_19096),
.B(n_8531),
.Y(n_19262)
);

INVx1_ASAP7_75t_L g19263 ( 
.A(n_19134),
.Y(n_19263)
);

NOR2x1_ASAP7_75t_L g19264 ( 
.A(n_19075),
.B(n_19035),
.Y(n_19264)
);

AOI211xp5_ASAP7_75t_L g19265 ( 
.A1(n_18860),
.A2(n_8650),
.B(n_8655),
.C(n_7543),
.Y(n_19265)
);

NAND2xp5_ASAP7_75t_L g19266 ( 
.A(n_19098),
.B(n_8546),
.Y(n_19266)
);

INVx1_ASAP7_75t_L g19267 ( 
.A(n_18958),
.Y(n_19267)
);

NOR2xp33_ASAP7_75t_L g19268 ( 
.A(n_19114),
.B(n_18896),
.Y(n_19268)
);

INVx1_ASAP7_75t_L g19269 ( 
.A(n_19120),
.Y(n_19269)
);

OAI21xp5_ASAP7_75t_L g19270 ( 
.A1(n_18898),
.A2(n_8237),
.B(n_8541),
.Y(n_19270)
);

OR2x2_ASAP7_75t_L g19271 ( 
.A(n_18917),
.B(n_8060),
.Y(n_19271)
);

OAI21xp5_ASAP7_75t_SL g19272 ( 
.A1(n_18883),
.A2(n_9032),
.B(n_9001),
.Y(n_19272)
);

INVx1_ASAP7_75t_L g19273 ( 
.A(n_18950),
.Y(n_19273)
);

INVx1_ASAP7_75t_L g19274 ( 
.A(n_18951),
.Y(n_19274)
);

INVx1_ASAP7_75t_L g19275 ( 
.A(n_18959),
.Y(n_19275)
);

INVx2_ASAP7_75t_L g19276 ( 
.A(n_19002),
.Y(n_19276)
);

OAI22x1_ASAP7_75t_L g19277 ( 
.A1(n_19067),
.A2(n_7543),
.B1(n_7931),
.B2(n_7906),
.Y(n_19277)
);

AND2x2_ASAP7_75t_L g19278 ( 
.A(n_19116),
.B(n_8694),
.Y(n_19278)
);

NAND3xp33_ASAP7_75t_L g19279 ( 
.A(n_19101),
.B(n_8631),
.C(n_8546),
.Y(n_19279)
);

AOI221xp5_ASAP7_75t_L g19280 ( 
.A1(n_19133),
.A2(n_19085),
.B1(n_19107),
.B2(n_18871),
.C(n_19119),
.Y(n_19280)
);

NAND2xp5_ASAP7_75t_L g19281 ( 
.A(n_19105),
.B(n_8546),
.Y(n_19281)
);

NOR2xp33_ASAP7_75t_L g19282 ( 
.A(n_19092),
.B(n_8631),
.Y(n_19282)
);

NOR2xp33_ASAP7_75t_SL g19283 ( 
.A(n_19082),
.B(n_7543),
.Y(n_19283)
);

NOR2xp33_ASAP7_75t_L g19284 ( 
.A(n_19108),
.B(n_8631),
.Y(n_19284)
);

INVx1_ASAP7_75t_L g19285 ( 
.A(n_18963),
.Y(n_19285)
);

INVx1_ASAP7_75t_L g19286 ( 
.A(n_18970),
.Y(n_19286)
);

OAI22xp5_ASAP7_75t_L g19287 ( 
.A1(n_18943),
.A2(n_9153),
.B1(n_9158),
.B2(n_9157),
.Y(n_19287)
);

INVx1_ASAP7_75t_L g19288 ( 
.A(n_19004),
.Y(n_19288)
);

NAND2xp5_ASAP7_75t_L g19289 ( 
.A(n_18990),
.B(n_8631),
.Y(n_19289)
);

NAND2x1_ASAP7_75t_L g19290 ( 
.A(n_19070),
.B(n_9537),
.Y(n_19290)
);

AND2x4_ASAP7_75t_L g19291 ( 
.A(n_19106),
.B(n_8060),
.Y(n_19291)
);

INVx1_ASAP7_75t_L g19292 ( 
.A(n_18973),
.Y(n_19292)
);

NOR2xp33_ASAP7_75t_L g19293 ( 
.A(n_19112),
.B(n_8639),
.Y(n_19293)
);

INVx1_ASAP7_75t_L g19294 ( 
.A(n_18947),
.Y(n_19294)
);

NAND2xp5_ASAP7_75t_L g19295 ( 
.A(n_19024),
.B(n_8639),
.Y(n_19295)
);

INVx1_ASAP7_75t_L g19296 ( 
.A(n_19011),
.Y(n_19296)
);

OAI221xp5_ASAP7_75t_L g19297 ( 
.A1(n_18915),
.A2(n_8357),
.B1(n_8428),
.B2(n_8330),
.C(n_8197),
.Y(n_19297)
);

INVxp67_ASAP7_75t_L g19298 ( 
.A(n_19118),
.Y(n_19298)
);

INVx1_ASAP7_75t_L g19299 ( 
.A(n_19025),
.Y(n_19299)
);

AND2x2_ASAP7_75t_L g19300 ( 
.A(n_19031),
.B(n_8694),
.Y(n_19300)
);

INVx1_ASAP7_75t_SL g19301 ( 
.A(n_19036),
.Y(n_19301)
);

AOI222xp33_ASAP7_75t_L g19302 ( 
.A1(n_19073),
.A2(n_8712),
.B1(n_8699),
.B2(n_8714),
.C1(n_8705),
.C2(n_8639),
.Y(n_19302)
);

OAI221xp5_ASAP7_75t_L g19303 ( 
.A1(n_19040),
.A2(n_8564),
.B1(n_8597),
.B2(n_8428),
.C(n_8357),
.Y(n_19303)
);

BUFx2_ASAP7_75t_L g19304 ( 
.A(n_19045),
.Y(n_19304)
);

NAND2xp5_ASAP7_75t_L g19305 ( 
.A(n_19041),
.B(n_8639),
.Y(n_19305)
);

OAI22xp33_ASAP7_75t_L g19306 ( 
.A1(n_19117),
.A2(n_8057),
.B1(n_8076),
.B2(n_8056),
.Y(n_19306)
);

NOR2x1p5_ASAP7_75t_L g19307 ( 
.A(n_18886),
.B(n_8056),
.Y(n_19307)
);

AOI21xp5_ASAP7_75t_L g19308 ( 
.A1(n_18888),
.A2(n_9181),
.B(n_9158),
.Y(n_19308)
);

OAI221xp5_ASAP7_75t_L g19309 ( 
.A1(n_18876),
.A2(n_8564),
.B1(n_8597),
.B2(n_8428),
.C(n_8357),
.Y(n_19309)
);

OAI221xp5_ASAP7_75t_L g19310 ( 
.A1(n_18862),
.A2(n_8597),
.B1(n_8610),
.B2(n_8564),
.C(n_8428),
.Y(n_19310)
);

OAI211xp5_ASAP7_75t_SL g19311 ( 
.A1(n_19125),
.A2(n_7910),
.B(n_7943),
.C(n_7916),
.Y(n_19311)
);

AND2x2_ASAP7_75t_L g19312 ( 
.A(n_19055),
.B(n_8123),
.Y(n_19312)
);

NOR2xp33_ASAP7_75t_L g19313 ( 
.A(n_19012),
.B(n_8699),
.Y(n_19313)
);

OAI22xp33_ASAP7_75t_SL g19314 ( 
.A1(n_19080),
.A2(n_9032),
.B1(n_9064),
.B2(n_9001),
.Y(n_19314)
);

INVx1_ASAP7_75t_L g19315 ( 
.A(n_19060),
.Y(n_19315)
);

OAI22xp5_ASAP7_75t_L g19316 ( 
.A1(n_19065),
.A2(n_9181),
.B1(n_9189),
.B2(n_9188),
.Y(n_19316)
);

OAI31xp33_ASAP7_75t_L g19317 ( 
.A1(n_18914),
.A2(n_9032),
.A3(n_9064),
.B(n_9001),
.Y(n_19317)
);

INVx1_ASAP7_75t_L g19318 ( 
.A(n_18904),
.Y(n_19318)
);

NAND2xp5_ASAP7_75t_L g19319 ( 
.A(n_18890),
.B(n_8699),
.Y(n_19319)
);

OAI21xp5_ASAP7_75t_SL g19320 ( 
.A1(n_18887),
.A2(n_9032),
.B(n_9001),
.Y(n_19320)
);

OAI221xp5_ASAP7_75t_L g19321 ( 
.A1(n_19097),
.A2(n_19126),
.B1(n_18923),
.B2(n_18999),
.C(n_18908),
.Y(n_19321)
);

AND2x2_ASAP7_75t_L g19322 ( 
.A(n_19072),
.B(n_7967),
.Y(n_19322)
);

OAI221xp5_ASAP7_75t_L g19323 ( 
.A1(n_19130),
.A2(n_18933),
.B1(n_19109),
.B2(n_18987),
.C(n_19023),
.Y(n_19323)
);

OR2x2_ASAP7_75t_L g19324 ( 
.A(n_19086),
.B(n_8066),
.Y(n_19324)
);

NAND2xp33_ASAP7_75t_SL g19325 ( 
.A(n_19113),
.B(n_7906),
.Y(n_19325)
);

NOR2xp33_ASAP7_75t_L g19326 ( 
.A(n_19046),
.B(n_8699),
.Y(n_19326)
);

O2A1O1Ixp33_ASAP7_75t_L g19327 ( 
.A1(n_19054),
.A2(n_7934),
.B(n_8712),
.C(n_8705),
.Y(n_19327)
);

AOI21xp33_ASAP7_75t_L g19328 ( 
.A1(n_19128),
.A2(n_8729),
.B(n_8690),
.Y(n_19328)
);

AND2x2_ASAP7_75t_L g19329 ( 
.A(n_19110),
.B(n_7967),
.Y(n_19329)
);

OAI21xp5_ASAP7_75t_L g19330 ( 
.A1(n_19068),
.A2(n_8541),
.B(n_8390),
.Y(n_19330)
);

NAND2xp5_ASAP7_75t_L g19331 ( 
.A(n_19078),
.B(n_8705),
.Y(n_19331)
);

INVx1_ASAP7_75t_SL g19332 ( 
.A(n_19071),
.Y(n_19332)
);

NAND2xp33_ASAP7_75t_R g19333 ( 
.A(n_19084),
.B(n_8655),
.Y(n_19333)
);

HB1xp67_ASAP7_75t_L g19334 ( 
.A(n_19010),
.Y(n_19334)
);

AND2x2_ASAP7_75t_L g19335 ( 
.A(n_19001),
.B(n_19005),
.Y(n_19335)
);

AND2x2_ASAP7_75t_L g19336 ( 
.A(n_18916),
.B(n_7967),
.Y(n_19336)
);

O2A1O1Ixp33_ASAP7_75t_L g19337 ( 
.A1(n_19094),
.A2(n_7934),
.B(n_8712),
.C(n_8705),
.Y(n_19337)
);

AND2x2_ASAP7_75t_SL g19338 ( 
.A(n_19048),
.B(n_9238),
.Y(n_19338)
);

OAI221xp5_ASAP7_75t_L g19339 ( 
.A1(n_18962),
.A2(n_8597),
.B1(n_8610),
.B2(n_8564),
.C(n_8428),
.Y(n_19339)
);

NAND2xp5_ASAP7_75t_L g19340 ( 
.A(n_18988),
.B(n_8712),
.Y(n_19340)
);

AOI22xp5_ASAP7_75t_L g19341 ( 
.A1(n_19111),
.A2(n_8732),
.B1(n_8751),
.B2(n_8714),
.Y(n_19341)
);

OAI22xp5_ASAP7_75t_L g19342 ( 
.A1(n_19103),
.A2(n_9181),
.B1(n_9189),
.B2(n_9188),
.Y(n_19342)
);

OR2x2_ASAP7_75t_L g19343 ( 
.A(n_19124),
.B(n_8066),
.Y(n_19343)
);

OAI21xp33_ASAP7_75t_L g19344 ( 
.A1(n_18905),
.A2(n_7762),
.B(n_7755),
.Y(n_19344)
);

INVx1_ASAP7_75t_SL g19345 ( 
.A(n_18968),
.Y(n_19345)
);

AND2x2_ASAP7_75t_L g19346 ( 
.A(n_18953),
.B(n_19123),
.Y(n_19346)
);

AOI221xp5_ASAP7_75t_L g19347 ( 
.A1(n_19122),
.A2(n_6955),
.B1(n_8732),
.B2(n_8751),
.C(n_8714),
.Y(n_19347)
);

NAND2xp33_ASAP7_75t_SL g19348 ( 
.A(n_19052),
.B(n_7906),
.Y(n_19348)
);

AND2x2_ASAP7_75t_L g19349 ( 
.A(n_18895),
.B(n_7967),
.Y(n_19349)
);

INVxp67_ASAP7_75t_L g19350 ( 
.A(n_19102),
.Y(n_19350)
);

NAND2xp5_ASAP7_75t_L g19351 ( 
.A(n_19016),
.B(n_8714),
.Y(n_19351)
);

O2A1O1Ixp33_ASAP7_75t_SL g19352 ( 
.A1(n_18899),
.A2(n_7394),
.B(n_7017),
.C(n_7034),
.Y(n_19352)
);

INVx1_ASAP7_75t_L g19353 ( 
.A(n_19050),
.Y(n_19353)
);

OAI211xp5_ASAP7_75t_SL g19354 ( 
.A1(n_18945),
.A2(n_7910),
.B(n_7943),
.C(n_7916),
.Y(n_19354)
);

O2A1O1Ixp5_ASAP7_75t_L g19355 ( 
.A1(n_18957),
.A2(n_9189),
.B(n_9192),
.C(n_9188),
.Y(n_19355)
);

AOI21xp33_ASAP7_75t_L g19356 ( 
.A1(n_19100),
.A2(n_8729),
.B(n_8690),
.Y(n_19356)
);

INVxp67_ASAP7_75t_SL g19357 ( 
.A(n_19026),
.Y(n_19357)
);

OAI21xp5_ASAP7_75t_L g19358 ( 
.A1(n_19064),
.A2(n_8541),
.B(n_8390),
.Y(n_19358)
);

NAND2xp5_ASAP7_75t_L g19359 ( 
.A(n_18944),
.B(n_8732),
.Y(n_19359)
);

INVx1_ASAP7_75t_L g19360 ( 
.A(n_19058),
.Y(n_19360)
);

AOI21xp33_ASAP7_75t_SL g19361 ( 
.A1(n_18900),
.A2(n_8597),
.B(n_8564),
.Y(n_19361)
);

OAI322xp33_ASAP7_75t_L g19362 ( 
.A1(n_19077),
.A2(n_9217),
.A3(n_9203),
.B1(n_9227),
.B2(n_9268),
.C1(n_9211),
.C2(n_9192),
.Y(n_19362)
);

INVx2_ASAP7_75t_L g19363 ( 
.A(n_18996),
.Y(n_19363)
);

AOI21xp5_ASAP7_75t_L g19364 ( 
.A1(n_19003),
.A2(n_9203),
.B(n_9192),
.Y(n_19364)
);

HB1xp67_ASAP7_75t_L g19365 ( 
.A(n_18918),
.Y(n_19365)
);

AND2x2_ASAP7_75t_L g19366 ( 
.A(n_18910),
.B(n_8038),
.Y(n_19366)
);

INVxp67_ASAP7_75t_SL g19367 ( 
.A(n_19009),
.Y(n_19367)
);

INVx1_ASAP7_75t_L g19368 ( 
.A(n_19006),
.Y(n_19368)
);

INVx1_ASAP7_75t_L g19369 ( 
.A(n_19038),
.Y(n_19369)
);

AOI21xp5_ASAP7_75t_L g19370 ( 
.A1(n_18956),
.A2(n_9211),
.B(n_9203),
.Y(n_19370)
);

INVx1_ASAP7_75t_L g19371 ( 
.A(n_18961),
.Y(n_19371)
);

OAI22xp5_ASAP7_75t_L g19372 ( 
.A1(n_18891),
.A2(n_9211),
.B1(n_9227),
.B2(n_9217),
.Y(n_19372)
);

INVx1_ASAP7_75t_L g19373 ( 
.A(n_18976),
.Y(n_19373)
);

NAND2xp5_ASAP7_75t_L g19374 ( 
.A(n_19121),
.B(n_8732),
.Y(n_19374)
);

OAI22xp5_ASAP7_75t_L g19375 ( 
.A1(n_19136),
.A2(n_9217),
.B1(n_9268),
.B2(n_9227),
.Y(n_19375)
);

NAND2xp5_ASAP7_75t_SL g19376 ( 
.A(n_19115),
.B(n_6955),
.Y(n_19376)
);

NOR2xp33_ASAP7_75t_L g19377 ( 
.A(n_19093),
.B(n_19069),
.Y(n_19377)
);

INVx1_ASAP7_75t_L g19378 ( 
.A(n_18960),
.Y(n_19378)
);

OAI33xp33_ASAP7_75t_L g19379 ( 
.A1(n_19059),
.A2(n_9282),
.A3(n_9269),
.B1(n_9289),
.B2(n_9272),
.B3(n_9268),
.Y(n_19379)
);

INVx2_ASAP7_75t_L g19380 ( 
.A(n_18996),
.Y(n_19380)
);

AOI21xp5_ASAP7_75t_L g19381 ( 
.A1(n_18894),
.A2(n_9272),
.B(n_9269),
.Y(n_19381)
);

NAND2xp5_ASAP7_75t_L g19382 ( 
.A(n_19104),
.B(n_8751),
.Y(n_19382)
);

INVx1_ASAP7_75t_L g19383 ( 
.A(n_18985),
.Y(n_19383)
);

NOR3xp33_ASAP7_75t_L g19384 ( 
.A(n_19029),
.B(n_8708),
.C(n_8333),
.Y(n_19384)
);

AND2x2_ASAP7_75t_L g19385 ( 
.A(n_18911),
.B(n_8038),
.Y(n_19385)
);

OAI22xp33_ASAP7_75t_L g19386 ( 
.A1(n_18912),
.A2(n_8057),
.B1(n_8076),
.B2(n_8056),
.Y(n_19386)
);

INVx1_ASAP7_75t_L g19387 ( 
.A(n_19091),
.Y(n_19387)
);

INVx2_ASAP7_75t_L g19388 ( 
.A(n_18997),
.Y(n_19388)
);

INVx2_ASAP7_75t_L g19389 ( 
.A(n_19039),
.Y(n_19389)
);

AOI21xp5_ASAP7_75t_L g19390 ( 
.A1(n_19095),
.A2(n_9272),
.B(n_9269),
.Y(n_19390)
);

NAND2xp33_ASAP7_75t_L g19391 ( 
.A(n_19127),
.B(n_6977),
.Y(n_19391)
);

NOR2xp33_ASAP7_75t_L g19392 ( 
.A(n_18981),
.B(n_8751),
.Y(n_19392)
);

INVx1_ASAP7_75t_L g19393 ( 
.A(n_19022),
.Y(n_19393)
);

INVx1_ASAP7_75t_L g19394 ( 
.A(n_19044),
.Y(n_19394)
);

NAND2xp5_ASAP7_75t_L g19395 ( 
.A(n_18978),
.B(n_8752),
.Y(n_19395)
);

INVx1_ASAP7_75t_L g19396 ( 
.A(n_18901),
.Y(n_19396)
);

OAI32xp33_ASAP7_75t_L g19397 ( 
.A1(n_18954),
.A2(n_7369),
.A3(n_8057),
.B1(n_8104),
.B2(n_8076),
.Y(n_19397)
);

INVx1_ASAP7_75t_L g19398 ( 
.A(n_19017),
.Y(n_19398)
);

O2A1O1Ixp33_ASAP7_75t_L g19399 ( 
.A1(n_19034),
.A2(n_8752),
.B(n_8782),
.C(n_8770),
.Y(n_19399)
);

NAND2xp5_ASAP7_75t_SL g19400 ( 
.A(n_18892),
.B(n_19000),
.Y(n_19400)
);

AOI22xp5_ASAP7_75t_L g19401 ( 
.A1(n_18934),
.A2(n_8770),
.B1(n_8782),
.B2(n_8752),
.Y(n_19401)
);

NAND2xp5_ASAP7_75t_L g19402 ( 
.A(n_18906),
.B(n_8752),
.Y(n_19402)
);

INVx2_ASAP7_75t_L g19403 ( 
.A(n_18952),
.Y(n_19403)
);

NAND2xp5_ASAP7_75t_L g19404 ( 
.A(n_19141),
.B(n_8770),
.Y(n_19404)
);

AOI211xp5_ASAP7_75t_L g19405 ( 
.A1(n_18983),
.A2(n_9224),
.B(n_7371),
.C(n_8539),
.Y(n_19405)
);

OAI211xp5_ASAP7_75t_L g19406 ( 
.A1(n_18897),
.A2(n_7730),
.B(n_7164),
.C(n_8025),
.Y(n_19406)
);

AOI222xp33_ASAP7_75t_L g19407 ( 
.A1(n_19087),
.A2(n_8788),
.B1(n_8782),
.B2(n_8825),
.C1(n_8794),
.C2(n_8770),
.Y(n_19407)
);

AOI22xp5_ASAP7_75t_L g19408 ( 
.A1(n_19345),
.A2(n_19037),
.B1(n_19089),
.B2(n_19014),
.Y(n_19408)
);

OR2x2_ASAP7_75t_L g19409 ( 
.A(n_19145),
.B(n_8353),
.Y(n_19409)
);

INVx1_ASAP7_75t_L g19410 ( 
.A(n_19200),
.Y(n_19410)
);

INVx1_ASAP7_75t_L g19411 ( 
.A(n_19144),
.Y(n_19411)
);

OR2x2_ASAP7_75t_L g19412 ( 
.A(n_19157),
.B(n_8353),
.Y(n_19412)
);

INVx1_ASAP7_75t_L g19413 ( 
.A(n_19150),
.Y(n_19413)
);

INVx1_ASAP7_75t_SL g19414 ( 
.A(n_19177),
.Y(n_19414)
);

HB1xp67_ASAP7_75t_L g19415 ( 
.A(n_19165),
.Y(n_19415)
);

INVx2_ASAP7_75t_SL g19416 ( 
.A(n_19223),
.Y(n_19416)
);

NOR2xp33_ASAP7_75t_L g19417 ( 
.A(n_19146),
.B(n_8782),
.Y(n_19417)
);

OR2x2_ASAP7_75t_L g19418 ( 
.A(n_19181),
.B(n_8353),
.Y(n_19418)
);

OR2x2_ASAP7_75t_L g19419 ( 
.A(n_19230),
.B(n_8353),
.Y(n_19419)
);

NAND2xp5_ASAP7_75t_L g19420 ( 
.A(n_19238),
.B(n_8788),
.Y(n_19420)
);

AND2x2_ASAP7_75t_L g19421 ( 
.A(n_19191),
.B(n_9224),
.Y(n_19421)
);

INVx1_ASAP7_75t_L g19422 ( 
.A(n_19162),
.Y(n_19422)
);

AND2x2_ASAP7_75t_L g19423 ( 
.A(n_19264),
.B(n_9224),
.Y(n_19423)
);

AND2x2_ASAP7_75t_L g19424 ( 
.A(n_19196),
.B(n_9558),
.Y(n_19424)
);

INVx1_ASAP7_75t_L g19425 ( 
.A(n_19166),
.Y(n_19425)
);

INVx2_ASAP7_75t_L g19426 ( 
.A(n_19237),
.Y(n_19426)
);

INVxp67_ASAP7_75t_L g19427 ( 
.A(n_19225),
.Y(n_19427)
);

NAND2x1_ASAP7_75t_L g19428 ( 
.A(n_19179),
.B(n_8711),
.Y(n_19428)
);

INVx1_ASAP7_75t_L g19429 ( 
.A(n_19169),
.Y(n_19429)
);

INVx1_ASAP7_75t_L g19430 ( 
.A(n_19247),
.Y(n_19430)
);

INVx1_ASAP7_75t_L g19431 ( 
.A(n_19224),
.Y(n_19431)
);

NAND2xp5_ASAP7_75t_SL g19432 ( 
.A(n_19186),
.B(n_8788),
.Y(n_19432)
);

INVx2_ASAP7_75t_L g19433 ( 
.A(n_19307),
.Y(n_19433)
);

AND2x2_ASAP7_75t_L g19434 ( 
.A(n_19212),
.B(n_19201),
.Y(n_19434)
);

INVx3_ASAP7_75t_L g19435 ( 
.A(n_19291),
.Y(n_19435)
);

INVx2_ASAP7_75t_L g19436 ( 
.A(n_19194),
.Y(n_19436)
);

NAND2xp5_ASAP7_75t_L g19437 ( 
.A(n_19335),
.B(n_8788),
.Y(n_19437)
);

CKINVDCx16_ASAP7_75t_R g19438 ( 
.A(n_19193),
.Y(n_19438)
);

NAND2xp5_ASAP7_75t_SL g19439 ( 
.A(n_19154),
.B(n_8794),
.Y(n_19439)
);

AOI22xp33_ASAP7_75t_L g19440 ( 
.A1(n_19304),
.A2(n_8825),
.B1(n_8842),
.B2(n_8794),
.Y(n_19440)
);

INVx1_ASAP7_75t_L g19441 ( 
.A(n_19245),
.Y(n_19441)
);

INVx1_ASAP7_75t_L g19442 ( 
.A(n_19248),
.Y(n_19442)
);

NOR2x1p5_ASAP7_75t_L g19443 ( 
.A(n_19164),
.B(n_19175),
.Y(n_19443)
);

AOI222xp33_ASAP7_75t_L g19444 ( 
.A1(n_19325),
.A2(n_8842),
.B1(n_8825),
.B2(n_8863),
.C1(n_8857),
.C2(n_8794),
.Y(n_19444)
);

NAND2xp5_ASAP7_75t_L g19445 ( 
.A(n_19334),
.B(n_8825),
.Y(n_19445)
);

AND2x2_ASAP7_75t_L g19446 ( 
.A(n_19349),
.B(n_19214),
.Y(n_19446)
);

NAND2xp5_ASAP7_75t_L g19447 ( 
.A(n_19368),
.B(n_8842),
.Y(n_19447)
);

INVx1_ASAP7_75t_L g19448 ( 
.A(n_19252),
.Y(n_19448)
);

INVxp67_ASAP7_75t_L g19449 ( 
.A(n_19203),
.Y(n_19449)
);

NAND2xp33_ASAP7_75t_SL g19450 ( 
.A(n_19250),
.B(n_7906),
.Y(n_19450)
);

INVx1_ASAP7_75t_L g19451 ( 
.A(n_19254),
.Y(n_19451)
);

NAND2xp5_ASAP7_75t_L g19452 ( 
.A(n_19276),
.B(n_8842),
.Y(n_19452)
);

AOI22xp33_ASAP7_75t_L g19453 ( 
.A1(n_19396),
.A2(n_8863),
.B1(n_8874),
.B2(n_8857),
.Y(n_19453)
);

INVx1_ASAP7_75t_L g19454 ( 
.A(n_19257),
.Y(n_19454)
);

AND2x2_ASAP7_75t_L g19455 ( 
.A(n_19236),
.B(n_9558),
.Y(n_19455)
);

OR2x2_ASAP7_75t_L g19456 ( 
.A(n_19221),
.B(n_8353),
.Y(n_19456)
);

INVx1_ASAP7_75t_L g19457 ( 
.A(n_19189),
.Y(n_19457)
);

AND2x2_ASAP7_75t_SL g19458 ( 
.A(n_19190),
.B(n_19192),
.Y(n_19458)
);

AND2x4_ASAP7_75t_L g19459 ( 
.A(n_19217),
.B(n_8076),
.Y(n_19459)
);

AND2x2_ASAP7_75t_L g19460 ( 
.A(n_19184),
.B(n_9558),
.Y(n_19460)
);

NAND2xp5_ASAP7_75t_L g19461 ( 
.A(n_19318),
.B(n_8857),
.Y(n_19461)
);

INVx1_ASAP7_75t_L g19462 ( 
.A(n_19156),
.Y(n_19462)
);

NOR2xp33_ASAP7_75t_L g19463 ( 
.A(n_19332),
.B(n_8857),
.Y(n_19463)
);

INVx1_ASAP7_75t_L g19464 ( 
.A(n_19185),
.Y(n_19464)
);

NAND2xp5_ASAP7_75t_L g19465 ( 
.A(n_19363),
.B(n_8863),
.Y(n_19465)
);

INVx1_ASAP7_75t_L g19466 ( 
.A(n_19199),
.Y(n_19466)
);

INVx1_ASAP7_75t_L g19467 ( 
.A(n_19269),
.Y(n_19467)
);

INVx1_ASAP7_75t_L g19468 ( 
.A(n_19357),
.Y(n_19468)
);

AND2x2_ASAP7_75t_L g19469 ( 
.A(n_19215),
.B(n_8038),
.Y(n_19469)
);

INVx2_ASAP7_75t_L g19470 ( 
.A(n_19290),
.Y(n_19470)
);

NOR2xp33_ASAP7_75t_L g19471 ( 
.A(n_19380),
.B(n_8863),
.Y(n_19471)
);

INVx1_ASAP7_75t_L g19472 ( 
.A(n_19365),
.Y(n_19472)
);

INVx1_ASAP7_75t_SL g19473 ( 
.A(n_19151),
.Y(n_19473)
);

AND2x4_ASAP7_75t_L g19474 ( 
.A(n_19298),
.B(n_6977),
.Y(n_19474)
);

NAND2xp5_ASAP7_75t_L g19475 ( 
.A(n_19202),
.B(n_8874),
.Y(n_19475)
);

NAND2xp33_ASAP7_75t_SL g19476 ( 
.A(n_19147),
.B(n_7906),
.Y(n_19476)
);

OR2x2_ASAP7_75t_L g19477 ( 
.A(n_19204),
.B(n_8353),
.Y(n_19477)
);

NAND2xp5_ASAP7_75t_L g19478 ( 
.A(n_19253),
.B(n_8874),
.Y(n_19478)
);

INVx1_ASAP7_75t_L g19479 ( 
.A(n_19159),
.Y(n_19479)
);

INVx2_ASAP7_75t_L g19480 ( 
.A(n_19258),
.Y(n_19480)
);

AND2x2_ASAP7_75t_L g19481 ( 
.A(n_19288),
.B(n_8038),
.Y(n_19481)
);

AND2x2_ASAP7_75t_L g19482 ( 
.A(n_19292),
.B(n_8062),
.Y(n_19482)
);

INVx2_ASAP7_75t_SL g19483 ( 
.A(n_19291),
.Y(n_19483)
);

INVx2_ASAP7_75t_L g19484 ( 
.A(n_19249),
.Y(n_19484)
);

INVx2_ASAP7_75t_SL g19485 ( 
.A(n_19213),
.Y(n_19485)
);

NAND2xp5_ASAP7_75t_L g19486 ( 
.A(n_19268),
.B(n_8874),
.Y(n_19486)
);

AOI21xp5_ASAP7_75t_SL g19487 ( 
.A1(n_19294),
.A2(n_8104),
.B(n_7258),
.Y(n_19487)
);

AOI222xp33_ASAP7_75t_L g19488 ( 
.A1(n_19280),
.A2(n_8919),
.B1(n_8902),
.B2(n_8961),
.C1(n_8946),
.C2(n_8894),
.Y(n_19488)
);

INVx1_ASAP7_75t_L g19489 ( 
.A(n_19173),
.Y(n_19489)
);

INVxp67_ASAP7_75t_L g19490 ( 
.A(n_19267),
.Y(n_19490)
);

INVx2_ASAP7_75t_L g19491 ( 
.A(n_19338),
.Y(n_19491)
);

NOR2x1_ASAP7_75t_L g19492 ( 
.A(n_19241),
.B(n_8104),
.Y(n_19492)
);

NAND2xp5_ASAP7_75t_SL g19493 ( 
.A(n_19251),
.B(n_8894),
.Y(n_19493)
);

NAND2xp5_ASAP7_75t_L g19494 ( 
.A(n_19170),
.B(n_8894),
.Y(n_19494)
);

INVx1_ASAP7_75t_SL g19495 ( 
.A(n_19301),
.Y(n_19495)
);

AND2x2_ASAP7_75t_L g19496 ( 
.A(n_19385),
.B(n_8062),
.Y(n_19496)
);

INVxp67_ASAP7_75t_L g19497 ( 
.A(n_19367),
.Y(n_19497)
);

AND2x2_ASAP7_75t_L g19498 ( 
.A(n_19346),
.B(n_8062),
.Y(n_19498)
);

INVx1_ASAP7_75t_L g19499 ( 
.A(n_19262),
.Y(n_19499)
);

NAND2xp5_ASAP7_75t_L g19500 ( 
.A(n_19350),
.B(n_8894),
.Y(n_19500)
);

INVx1_ASAP7_75t_SL g19501 ( 
.A(n_19383),
.Y(n_19501)
);

AND2x2_ASAP7_75t_L g19502 ( 
.A(n_19336),
.B(n_8062),
.Y(n_19502)
);

NAND2xp5_ASAP7_75t_L g19503 ( 
.A(n_19273),
.B(n_8902),
.Y(n_19503)
);

INVx1_ASAP7_75t_SL g19504 ( 
.A(n_19274),
.Y(n_19504)
);

INVx2_ASAP7_75t_SL g19505 ( 
.A(n_19266),
.Y(n_19505)
);

OAI22xp5_ASAP7_75t_L g19506 ( 
.A1(n_19148),
.A2(n_9289),
.B1(n_9297),
.B2(n_9282),
.Y(n_19506)
);

NAND2xp5_ASAP7_75t_L g19507 ( 
.A(n_19275),
.B(n_8902),
.Y(n_19507)
);

AND2x2_ASAP7_75t_L g19508 ( 
.A(n_19312),
.B(n_9533),
.Y(n_19508)
);

NOR2x1_ASAP7_75t_L g19509 ( 
.A(n_19263),
.B(n_8104),
.Y(n_19509)
);

INVx3_ASAP7_75t_L g19510 ( 
.A(n_19244),
.Y(n_19510)
);

AND2x4_ASAP7_75t_L g19511 ( 
.A(n_19315),
.B(n_7017),
.Y(n_19511)
);

INVx1_ASAP7_75t_L g19512 ( 
.A(n_19281),
.Y(n_19512)
);

AND2x2_ASAP7_75t_L g19513 ( 
.A(n_19322),
.B(n_9541),
.Y(n_19513)
);

OAI222xp33_ASAP7_75t_L g19514 ( 
.A1(n_19321),
.A2(n_9138),
.B1(n_9103),
.B2(n_9147),
.C1(n_9126),
.C2(n_9064),
.Y(n_19514)
);

INVx1_ASAP7_75t_SL g19515 ( 
.A(n_19285),
.Y(n_19515)
);

NAND2x1_ASAP7_75t_L g19516 ( 
.A(n_19371),
.B(n_8711),
.Y(n_19516)
);

OR2x2_ASAP7_75t_L g19517 ( 
.A(n_19319),
.B(n_19359),
.Y(n_19517)
);

NAND2xp5_ASAP7_75t_L g19518 ( 
.A(n_19286),
.B(n_8902),
.Y(n_19518)
);

AOI222xp33_ASAP7_75t_L g19519 ( 
.A1(n_19326),
.A2(n_8961),
.B1(n_8946),
.B2(n_8973),
.C1(n_8963),
.C2(n_8919),
.Y(n_19519)
);

INVx1_ASAP7_75t_L g19520 ( 
.A(n_19227),
.Y(n_19520)
);

AOI222xp33_ASAP7_75t_L g19521 ( 
.A1(n_19376),
.A2(n_8961),
.B1(n_8946),
.B2(n_8973),
.C1(n_8963),
.C2(n_8919),
.Y(n_19521)
);

NOR2xp33_ASAP7_75t_L g19522 ( 
.A(n_19323),
.B(n_8919),
.Y(n_19522)
);

NOR2xp33_ASAP7_75t_L g19523 ( 
.A(n_19296),
.B(n_8946),
.Y(n_19523)
);

OAI22xp5_ASAP7_75t_L g19524 ( 
.A1(n_19158),
.A2(n_9289),
.B1(n_9297),
.B2(n_9282),
.Y(n_19524)
);

INVx1_ASAP7_75t_L g19525 ( 
.A(n_19228),
.Y(n_19525)
);

AND2x2_ASAP7_75t_L g19526 ( 
.A(n_19329),
.B(n_9541),
.Y(n_19526)
);

OR2x2_ASAP7_75t_L g19527 ( 
.A(n_19271),
.B(n_8353),
.Y(n_19527)
);

NAND2xp5_ASAP7_75t_L g19528 ( 
.A(n_19284),
.B(n_19282),
.Y(n_19528)
);

AND2x4_ASAP7_75t_L g19529 ( 
.A(n_19403),
.B(n_8104),
.Y(n_19529)
);

NAND2xp5_ASAP7_75t_L g19530 ( 
.A(n_19293),
.B(n_8961),
.Y(n_19530)
);

NAND2xp5_ASAP7_75t_L g19531 ( 
.A(n_19299),
.B(n_8963),
.Y(n_19531)
);

AND2x2_ASAP7_75t_L g19532 ( 
.A(n_19161),
.B(n_9542),
.Y(n_19532)
);

INVx1_ASAP7_75t_SL g19533 ( 
.A(n_19389),
.Y(n_19533)
);

INVx1_ASAP7_75t_L g19534 ( 
.A(n_19259),
.Y(n_19534)
);

NOR2x1_ASAP7_75t_L g19535 ( 
.A(n_19387),
.B(n_7694),
.Y(n_19535)
);

INVx1_ASAP7_75t_L g19536 ( 
.A(n_19240),
.Y(n_19536)
);

INVx1_ASAP7_75t_L g19537 ( 
.A(n_19242),
.Y(n_19537)
);

CKINVDCx16_ASAP7_75t_R g19538 ( 
.A(n_19388),
.Y(n_19538)
);

INVx2_ASAP7_75t_SL g19539 ( 
.A(n_19398),
.Y(n_19539)
);

INVx1_ASAP7_75t_L g19540 ( 
.A(n_19180),
.Y(n_19540)
);

HB1xp67_ASAP7_75t_L g19541 ( 
.A(n_19373),
.Y(n_19541)
);

INVx1_ASAP7_75t_L g19542 ( 
.A(n_19369),
.Y(n_19542)
);

AND2x2_ASAP7_75t_L g19543 ( 
.A(n_19283),
.B(n_9542),
.Y(n_19543)
);

NOR2xp33_ASAP7_75t_L g19544 ( 
.A(n_19393),
.B(n_8963),
.Y(n_19544)
);

INVxp67_ASAP7_75t_L g19545 ( 
.A(n_19394),
.Y(n_19545)
);

NAND2xp5_ASAP7_75t_L g19546 ( 
.A(n_19143),
.B(n_8973),
.Y(n_19546)
);

AOI22xp33_ASAP7_75t_L g19547 ( 
.A1(n_19163),
.A2(n_8976),
.B1(n_8990),
.B2(n_8973),
.Y(n_19547)
);

INVx1_ASAP7_75t_L g19548 ( 
.A(n_19353),
.Y(n_19548)
);

NAND2xp5_ASAP7_75t_L g19549 ( 
.A(n_19261),
.B(n_8976),
.Y(n_19549)
);

INVx1_ASAP7_75t_L g19550 ( 
.A(n_19360),
.Y(n_19550)
);

NOR2xp67_ASAP7_75t_L g19551 ( 
.A(n_19149),
.B(n_7034),
.Y(n_19551)
);

AND2x2_ASAP7_75t_L g19552 ( 
.A(n_19272),
.B(n_9542),
.Y(n_19552)
);

NOR2xp33_ASAP7_75t_L g19553 ( 
.A(n_19208),
.B(n_8976),
.Y(n_19553)
);

INVx1_ASAP7_75t_L g19554 ( 
.A(n_19378),
.Y(n_19554)
);

AND2x2_ASAP7_75t_L g19555 ( 
.A(n_19377),
.B(n_9546),
.Y(n_19555)
);

INVx1_ASAP7_75t_L g19556 ( 
.A(n_19239),
.Y(n_19556)
);

INVx1_ASAP7_75t_L g19557 ( 
.A(n_19324),
.Y(n_19557)
);

NAND2xp33_ASAP7_75t_L g19558 ( 
.A(n_19348),
.B(n_7075),
.Y(n_19558)
);

INVx1_ASAP7_75t_L g19559 ( 
.A(n_19343),
.Y(n_19559)
);

OR2x2_ASAP7_75t_L g19560 ( 
.A(n_19351),
.B(n_8353),
.Y(n_19560)
);

INVx1_ASAP7_75t_L g19561 ( 
.A(n_19308),
.Y(n_19561)
);

NAND2xp33_ASAP7_75t_R g19562 ( 
.A(n_19209),
.B(n_8025),
.Y(n_19562)
);

NOR2xp33_ASAP7_75t_L g19563 ( 
.A(n_19372),
.B(n_8976),
.Y(n_19563)
);

AND2x2_ASAP7_75t_L g19564 ( 
.A(n_19255),
.B(n_9546),
.Y(n_19564)
);

NAND2xp5_ASAP7_75t_L g19565 ( 
.A(n_19313),
.B(n_8990),
.Y(n_19565)
);

INVx1_ASAP7_75t_L g19566 ( 
.A(n_19352),
.Y(n_19566)
);

AND2x2_ASAP7_75t_L g19567 ( 
.A(n_19220),
.B(n_9546),
.Y(n_19567)
);

INVx3_ASAP7_75t_L g19568 ( 
.A(n_19289),
.Y(n_19568)
);

NAND2xp5_ASAP7_75t_SL g19569 ( 
.A(n_19182),
.B(n_8990),
.Y(n_19569)
);

BUFx2_ASAP7_75t_L g19570 ( 
.A(n_19295),
.Y(n_19570)
);

INVx1_ASAP7_75t_L g19571 ( 
.A(n_19391),
.Y(n_19571)
);

INVx1_ASAP7_75t_L g19572 ( 
.A(n_19355),
.Y(n_19572)
);

NOR2xp33_ASAP7_75t_L g19573 ( 
.A(n_19379),
.B(n_8990),
.Y(n_19573)
);

NAND2xp5_ASAP7_75t_L g19574 ( 
.A(n_19370),
.B(n_9014),
.Y(n_19574)
);

INVx1_ASAP7_75t_L g19575 ( 
.A(n_19305),
.Y(n_19575)
);

AND2x2_ASAP7_75t_L g19576 ( 
.A(n_19197),
.B(n_9547),
.Y(n_19576)
);

NAND2xp5_ASAP7_75t_L g19577 ( 
.A(n_19229),
.B(n_9014),
.Y(n_19577)
);

AND2x2_ASAP7_75t_L g19578 ( 
.A(n_19198),
.B(n_9547),
.Y(n_19578)
);

NAND2xp5_ASAP7_75t_L g19579 ( 
.A(n_19176),
.B(n_9014),
.Y(n_19579)
);

NOR2xp33_ASAP7_75t_L g19580 ( 
.A(n_19400),
.B(n_9014),
.Y(n_19580)
);

XNOR2xp5_ASAP7_75t_L g19581 ( 
.A(n_19406),
.B(n_19265),
.Y(n_19581)
);

AND2x2_ASAP7_75t_L g19582 ( 
.A(n_19243),
.B(n_9547),
.Y(n_19582)
);

OR2x2_ASAP7_75t_L g19583 ( 
.A(n_19340),
.B(n_8364),
.Y(n_19583)
);

NAND2xp5_ASAP7_75t_L g19584 ( 
.A(n_19327),
.B(n_9029),
.Y(n_19584)
);

NAND2xp5_ASAP7_75t_L g19585 ( 
.A(n_19218),
.B(n_9029),
.Y(n_19585)
);

NAND2xp5_ASAP7_75t_L g19586 ( 
.A(n_19331),
.B(n_9029),
.Y(n_19586)
);

AND2x2_ASAP7_75t_L g19587 ( 
.A(n_19207),
.B(n_9551),
.Y(n_19587)
);

NOR2xp33_ASAP7_75t_L g19588 ( 
.A(n_19205),
.B(n_9029),
.Y(n_19588)
);

AND2x2_ASAP7_75t_L g19589 ( 
.A(n_19277),
.B(n_9551),
.Y(n_19589)
);

NAND2xp5_ASAP7_75t_L g19590 ( 
.A(n_19382),
.B(n_9096),
.Y(n_19590)
);

INVx1_ASAP7_75t_L g19591 ( 
.A(n_19404),
.Y(n_19591)
);

NOR2xp33_ASAP7_75t_L g19592 ( 
.A(n_19354),
.B(n_9096),
.Y(n_19592)
);

NOR2xp33_ASAP7_75t_L g19593 ( 
.A(n_19397),
.B(n_9096),
.Y(n_19593)
);

AND2x2_ASAP7_75t_L g19594 ( 
.A(n_19278),
.B(n_9551),
.Y(n_19594)
);

NOR2xp33_ASAP7_75t_SL g19595 ( 
.A(n_19320),
.B(n_7164),
.Y(n_19595)
);

INVx1_ASAP7_75t_L g19596 ( 
.A(n_19195),
.Y(n_19596)
);

INVx1_ASAP7_75t_L g19597 ( 
.A(n_19316),
.Y(n_19597)
);

INVx3_ASAP7_75t_L g19598 ( 
.A(n_19366),
.Y(n_19598)
);

INVx1_ASAP7_75t_L g19599 ( 
.A(n_19375),
.Y(n_19599)
);

AND2x2_ASAP7_75t_L g19600 ( 
.A(n_19300),
.B(n_9552),
.Y(n_19600)
);

AND2x2_ASAP7_75t_L g19601 ( 
.A(n_19344),
.B(n_9552),
.Y(n_19601)
);

NAND2xp5_ASAP7_75t_L g19602 ( 
.A(n_19153),
.B(n_9096),
.Y(n_19602)
);

INVx1_ASAP7_75t_L g19603 ( 
.A(n_19152),
.Y(n_19603)
);

NOR2xp33_ASAP7_75t_SL g19604 ( 
.A(n_19317),
.B(n_7164),
.Y(n_19604)
);

INVx1_ASAP7_75t_L g19605 ( 
.A(n_19402),
.Y(n_19605)
);

NAND2xp5_ASAP7_75t_L g19606 ( 
.A(n_19234),
.B(n_9106),
.Y(n_19606)
);

INVx1_ASAP7_75t_SL g19607 ( 
.A(n_19395),
.Y(n_19607)
);

CKINVDCx20_ASAP7_75t_R g19608 ( 
.A(n_19374),
.Y(n_19608)
);

NAND2xp5_ASAP7_75t_L g19609 ( 
.A(n_19390),
.B(n_9106),
.Y(n_19609)
);

AOI22xp33_ASAP7_75t_L g19610 ( 
.A1(n_19384),
.A2(n_9116),
.B1(n_9123),
.B2(n_9106),
.Y(n_19610)
);

NOR2xp33_ASAP7_75t_L g19611 ( 
.A(n_19219),
.B(n_19232),
.Y(n_19611)
);

INVx1_ASAP7_75t_SL g19612 ( 
.A(n_19356),
.Y(n_19612)
);

OR2x2_ASAP7_75t_L g19613 ( 
.A(n_19279),
.B(n_8364),
.Y(n_19613)
);

NOR2xp33_ASAP7_75t_L g19614 ( 
.A(n_19155),
.B(n_9106),
.Y(n_19614)
);

NOR2xp33_ASAP7_75t_L g19615 ( 
.A(n_19235),
.B(n_9116),
.Y(n_19615)
);

OR2x2_ASAP7_75t_L g19616 ( 
.A(n_19339),
.B(n_8364),
.Y(n_19616)
);

INVx1_ASAP7_75t_SL g19617 ( 
.A(n_19328),
.Y(n_19617)
);

NOR3x1_ASAP7_75t_L g19618 ( 
.A(n_19168),
.B(n_9046),
.C(n_8648),
.Y(n_19618)
);

AND2x4_ASAP7_75t_L g19619 ( 
.A(n_19210),
.B(n_7075),
.Y(n_19619)
);

INVx1_ASAP7_75t_L g19620 ( 
.A(n_19337),
.Y(n_19620)
);

INVx1_ASAP7_75t_L g19621 ( 
.A(n_19216),
.Y(n_19621)
);

NAND2xp5_ASAP7_75t_L g19622 ( 
.A(n_19392),
.B(n_9116),
.Y(n_19622)
);

NOR2x1_ASAP7_75t_L g19623 ( 
.A(n_19362),
.B(n_7694),
.Y(n_19623)
);

CKINVDCx20_ASAP7_75t_R g19624 ( 
.A(n_19160),
.Y(n_19624)
);

INVx1_ASAP7_75t_L g19625 ( 
.A(n_19287),
.Y(n_19625)
);

AND2x2_ASAP7_75t_L g19626 ( 
.A(n_19226),
.B(n_19361),
.Y(n_19626)
);

OR2x2_ASAP7_75t_L g19627 ( 
.A(n_19306),
.B(n_8364),
.Y(n_19627)
);

INVx1_ASAP7_75t_L g19628 ( 
.A(n_19399),
.Y(n_19628)
);

AND2x2_ASAP7_75t_L g19629 ( 
.A(n_19302),
.B(n_9552),
.Y(n_19629)
);

OR2x2_ASAP7_75t_L g19630 ( 
.A(n_19233),
.B(n_8364),
.Y(n_19630)
);

NAND2x1p5_ASAP7_75t_L g19631 ( 
.A(n_19172),
.B(n_7394),
.Y(n_19631)
);

NOR2xp33_ASAP7_75t_L g19632 ( 
.A(n_19386),
.B(n_9116),
.Y(n_19632)
);

OR2x2_ASAP7_75t_L g19633 ( 
.A(n_19342),
.B(n_19330),
.Y(n_19633)
);

INVx3_ASAP7_75t_L g19634 ( 
.A(n_19222),
.Y(n_19634)
);

AOI222xp33_ASAP7_75t_L g19635 ( 
.A1(n_19347),
.A2(n_9151),
.B1(n_9145),
.B2(n_9168),
.C1(n_9155),
.C2(n_9123),
.Y(n_19635)
);

INVx1_ASAP7_75t_L g19636 ( 
.A(n_19183),
.Y(n_19636)
);

NOR2xp33_ASAP7_75t_L g19637 ( 
.A(n_19311),
.B(n_9123),
.Y(n_19637)
);

OR2x2_ASAP7_75t_L g19638 ( 
.A(n_19358),
.B(n_8364),
.Y(n_19638)
);

INVxp67_ASAP7_75t_L g19639 ( 
.A(n_19333),
.Y(n_19639)
);

OAI31xp33_ASAP7_75t_SL g19640 ( 
.A1(n_19178),
.A2(n_8641),
.A3(n_8648),
.B(n_8499),
.Y(n_19640)
);

INVx1_ASAP7_75t_L g19641 ( 
.A(n_19211),
.Y(n_19641)
);

NAND2xp5_ASAP7_75t_L g19642 ( 
.A(n_19231),
.B(n_9123),
.Y(n_19642)
);

OR2x6_ASAP7_75t_L g19643 ( 
.A(n_19364),
.B(n_9193),
.Y(n_19643)
);

AND2x2_ASAP7_75t_L g19644 ( 
.A(n_19405),
.B(n_9557),
.Y(n_19644)
);

NAND2xp5_ASAP7_75t_L g19645 ( 
.A(n_19171),
.B(n_9145),
.Y(n_19645)
);

OAI22xp5_ASAP7_75t_L g19646 ( 
.A1(n_19174),
.A2(n_9302),
.B1(n_9309),
.B2(n_9297),
.Y(n_19646)
);

OR2x2_ASAP7_75t_L g19647 ( 
.A(n_19381),
.B(n_8364),
.Y(n_19647)
);

INVx1_ASAP7_75t_L g19648 ( 
.A(n_19167),
.Y(n_19648)
);

INVx1_ASAP7_75t_SL g19649 ( 
.A(n_19401),
.Y(n_19649)
);

INVx1_ASAP7_75t_L g19650 ( 
.A(n_19341),
.Y(n_19650)
);

AOI22xp5_ASAP7_75t_L g19651 ( 
.A1(n_19407),
.A2(n_9151),
.B1(n_9155),
.B2(n_9145),
.Y(n_19651)
);

AOI221xp5_ASAP7_75t_L g19652 ( 
.A1(n_19270),
.A2(n_9155),
.B1(n_9168),
.B2(n_9151),
.C(n_9145),
.Y(n_19652)
);

NOR2xp33_ASAP7_75t_L g19653 ( 
.A(n_19309),
.B(n_9151),
.Y(n_19653)
);

AND2x2_ASAP7_75t_L g19654 ( 
.A(n_19188),
.B(n_9557),
.Y(n_19654)
);

NAND2xp5_ASAP7_75t_L g19655 ( 
.A(n_19246),
.B(n_19260),
.Y(n_19655)
);

HB1xp67_ASAP7_75t_L g19656 ( 
.A(n_19310),
.Y(n_19656)
);

NAND2xp5_ASAP7_75t_L g19657 ( 
.A(n_19314),
.B(n_9155),
.Y(n_19657)
);

NAND3x1_ASAP7_75t_L g19658 ( 
.A(n_19187),
.B(n_9309),
.C(n_9302),
.Y(n_19658)
);

INVx1_ASAP7_75t_SL g19659 ( 
.A(n_19303),
.Y(n_19659)
);

HB1xp67_ASAP7_75t_L g19660 ( 
.A(n_19297),
.Y(n_19660)
);

INVx1_ASAP7_75t_L g19661 ( 
.A(n_19206),
.Y(n_19661)
);

INVx1_ASAP7_75t_L g19662 ( 
.A(n_19256),
.Y(n_19662)
);

INVx2_ASAP7_75t_L g19663 ( 
.A(n_19200),
.Y(n_19663)
);

NAND2xp5_ASAP7_75t_L g19664 ( 
.A(n_19144),
.B(n_9168),
.Y(n_19664)
);

INVx1_ASAP7_75t_L g19665 ( 
.A(n_19200),
.Y(n_19665)
);

INVx1_ASAP7_75t_L g19666 ( 
.A(n_19200),
.Y(n_19666)
);

INVx1_ASAP7_75t_SL g19667 ( 
.A(n_19200),
.Y(n_19667)
);

INVx1_ASAP7_75t_SL g19668 ( 
.A(n_19200),
.Y(n_19668)
);

AOI222xp33_ASAP7_75t_L g19669 ( 
.A1(n_19146),
.A2(n_9200),
.B1(n_9178),
.B2(n_9212),
.C1(n_9208),
.C2(n_9168),
.Y(n_19669)
);

INVx2_ASAP7_75t_L g19670 ( 
.A(n_19416),
.Y(n_19670)
);

NAND2xp5_ASAP7_75t_L g19671 ( 
.A(n_19438),
.B(n_9178),
.Y(n_19671)
);

NAND2xp5_ASAP7_75t_SL g19672 ( 
.A(n_19667),
.B(n_9178),
.Y(n_19672)
);

INVx1_ASAP7_75t_L g19673 ( 
.A(n_19415),
.Y(n_19673)
);

AO22x2_ASAP7_75t_L g19674 ( 
.A1(n_19668),
.A2(n_9178),
.B1(n_9208),
.B2(n_9200),
.Y(n_19674)
);

AND2x2_ASAP7_75t_L g19675 ( 
.A(n_19434),
.B(n_9535),
.Y(n_19675)
);

XNOR2x1_ASAP7_75t_L g19676 ( 
.A(n_19473),
.B(n_8610),
.Y(n_19676)
);

NAND2xp5_ASAP7_75t_L g19677 ( 
.A(n_19414),
.B(n_9200),
.Y(n_19677)
);

INVx1_ASAP7_75t_L g19678 ( 
.A(n_19663),
.Y(n_19678)
);

NOR2xp33_ASAP7_75t_L g19679 ( 
.A(n_19497),
.B(n_9200),
.Y(n_19679)
);

INVx1_ASAP7_75t_L g19680 ( 
.A(n_19410),
.Y(n_19680)
);

INVx1_ASAP7_75t_SL g19681 ( 
.A(n_19458),
.Y(n_19681)
);

NAND2xp5_ASAP7_75t_L g19682 ( 
.A(n_19533),
.B(n_9208),
.Y(n_19682)
);

INVx1_ASAP7_75t_SL g19683 ( 
.A(n_19665),
.Y(n_19683)
);

INVx1_ASAP7_75t_L g19684 ( 
.A(n_19666),
.Y(n_19684)
);

CKINVDCx5p33_ASAP7_75t_R g19685 ( 
.A(n_19538),
.Y(n_19685)
);

OR2x2_ASAP7_75t_L g19686 ( 
.A(n_19501),
.B(n_8364),
.Y(n_19686)
);

INVx1_ASAP7_75t_L g19687 ( 
.A(n_19541),
.Y(n_19687)
);

INVx1_ASAP7_75t_L g19688 ( 
.A(n_19472),
.Y(n_19688)
);

NAND2xp5_ASAP7_75t_L g19689 ( 
.A(n_19639),
.B(n_9208),
.Y(n_19689)
);

NOR2xp33_ASAP7_75t_L g19690 ( 
.A(n_19427),
.B(n_9212),
.Y(n_19690)
);

AND2x2_ASAP7_75t_L g19691 ( 
.A(n_19498),
.B(n_9535),
.Y(n_19691)
);

NAND2xp5_ASAP7_75t_L g19692 ( 
.A(n_19435),
.B(n_19483),
.Y(n_19692)
);

INVx2_ASAP7_75t_L g19693 ( 
.A(n_19443),
.Y(n_19693)
);

INVx1_ASAP7_75t_L g19694 ( 
.A(n_19426),
.Y(n_19694)
);

XNOR2x1_ASAP7_75t_L g19695 ( 
.A(n_19495),
.B(n_8610),
.Y(n_19695)
);

INVx1_ASAP7_75t_L g19696 ( 
.A(n_19462),
.Y(n_19696)
);

NOR2xp33_ASAP7_75t_L g19697 ( 
.A(n_19490),
.B(n_9212),
.Y(n_19697)
);

NAND2xp5_ASAP7_75t_L g19698 ( 
.A(n_19423),
.B(n_9212),
.Y(n_19698)
);

INVx1_ASAP7_75t_L g19699 ( 
.A(n_19430),
.Y(n_19699)
);

OR2x2_ASAP7_75t_L g19700 ( 
.A(n_19431),
.B(n_9292),
.Y(n_19700)
);

NAND2xp5_ASAP7_75t_SL g19701 ( 
.A(n_19422),
.B(n_9231),
.Y(n_19701)
);

INVx2_ASAP7_75t_L g19702 ( 
.A(n_19428),
.Y(n_19702)
);

NAND2xp5_ASAP7_75t_L g19703 ( 
.A(n_19468),
.B(n_9231),
.Y(n_19703)
);

HB1xp67_ASAP7_75t_L g19704 ( 
.A(n_19509),
.Y(n_19704)
);

INVx1_ASAP7_75t_L g19705 ( 
.A(n_19539),
.Y(n_19705)
);

NAND2xp33_ASAP7_75t_R g19706 ( 
.A(n_19446),
.B(n_8028),
.Y(n_19706)
);

AND2x2_ASAP7_75t_L g19707 ( 
.A(n_19459),
.B(n_9535),
.Y(n_19707)
);

INVx1_ASAP7_75t_L g19708 ( 
.A(n_19411),
.Y(n_19708)
);

OR2x2_ASAP7_75t_L g19709 ( 
.A(n_19504),
.B(n_19515),
.Y(n_19709)
);

XOR2xp5_ASAP7_75t_L g19710 ( 
.A(n_19581),
.B(n_8610),
.Y(n_19710)
);

INVxp67_ASAP7_75t_SL g19711 ( 
.A(n_19441),
.Y(n_19711)
);

INVx1_ASAP7_75t_SL g19712 ( 
.A(n_19442),
.Y(n_19712)
);

INVx1_ASAP7_75t_L g19713 ( 
.A(n_19448),
.Y(n_19713)
);

NAND2xp33_ASAP7_75t_L g19714 ( 
.A(n_19467),
.B(n_7078),
.Y(n_19714)
);

HB1xp67_ASAP7_75t_L g19715 ( 
.A(n_19545),
.Y(n_19715)
);

NAND2xp5_ASAP7_75t_SL g19716 ( 
.A(n_19451),
.B(n_9231),
.Y(n_19716)
);

INVx1_ASAP7_75t_L g19717 ( 
.A(n_19454),
.Y(n_19717)
);

NAND2xp5_ASAP7_75t_L g19718 ( 
.A(n_19505),
.B(n_9231),
.Y(n_19718)
);

NAND2xp5_ASAP7_75t_L g19719 ( 
.A(n_19466),
.B(n_9241),
.Y(n_19719)
);

NAND2xp5_ASAP7_75t_L g19720 ( 
.A(n_19529),
.B(n_9241),
.Y(n_19720)
);

AOI21xp33_ASAP7_75t_L g19721 ( 
.A1(n_19429),
.A2(n_8729),
.B(n_8690),
.Y(n_19721)
);

INVx1_ASAP7_75t_L g19722 ( 
.A(n_19457),
.Y(n_19722)
);

NAND2xp5_ASAP7_75t_L g19723 ( 
.A(n_19570),
.B(n_9241),
.Y(n_19723)
);

INVx1_ASAP7_75t_L g19724 ( 
.A(n_19413),
.Y(n_19724)
);

OAI21xp5_ASAP7_75t_SL g19725 ( 
.A1(n_19546),
.A2(n_7274),
.B(n_9064),
.Y(n_19725)
);

INVx1_ASAP7_75t_L g19726 ( 
.A(n_19437),
.Y(n_19726)
);

NOR2xp33_ASAP7_75t_L g19727 ( 
.A(n_19607),
.B(n_9241),
.Y(n_19727)
);

INVx1_ASAP7_75t_L g19728 ( 
.A(n_19542),
.Y(n_19728)
);

NAND2xp5_ASAP7_75t_L g19729 ( 
.A(n_19568),
.B(n_9243),
.Y(n_19729)
);

INVx1_ASAP7_75t_L g19730 ( 
.A(n_19535),
.Y(n_19730)
);

INVx1_ASAP7_75t_L g19731 ( 
.A(n_19492),
.Y(n_19731)
);

INVx1_ASAP7_75t_L g19732 ( 
.A(n_19420),
.Y(n_19732)
);

XOR2x2_ASAP7_75t_L g19733 ( 
.A(n_19516),
.B(n_8697),
.Y(n_19733)
);

AOI322xp5_ASAP7_75t_L g19734 ( 
.A1(n_19548),
.A2(n_7041),
.A3(n_8798),
.B1(n_7520),
.B2(n_9308),
.C1(n_9311),
.C2(n_9243),
.Y(n_19734)
);

NAND2xp5_ASAP7_75t_L g19735 ( 
.A(n_19424),
.B(n_9243),
.Y(n_19735)
);

NOR4xp25_ASAP7_75t_SL g19736 ( 
.A(n_19425),
.B(n_19464),
.C(n_19559),
.D(n_19557),
.Y(n_19736)
);

INVx1_ASAP7_75t_L g19737 ( 
.A(n_19474),
.Y(n_19737)
);

NAND2xp5_ASAP7_75t_L g19738 ( 
.A(n_19551),
.B(n_9243),
.Y(n_19738)
);

INVx1_ASAP7_75t_L g19739 ( 
.A(n_19474),
.Y(n_19739)
);

AOI21xp33_ASAP7_75t_L g19740 ( 
.A1(n_19517),
.A2(n_8690),
.B(n_9308),
.Y(n_19740)
);

INVx1_ASAP7_75t_L g19741 ( 
.A(n_19419),
.Y(n_19741)
);

AND2x2_ASAP7_75t_L g19742 ( 
.A(n_19481),
.B(n_9535),
.Y(n_19742)
);

AND2x2_ASAP7_75t_L g19743 ( 
.A(n_19482),
.B(n_9535),
.Y(n_19743)
);

OAI21xp5_ASAP7_75t_SL g19744 ( 
.A1(n_19449),
.A2(n_7274),
.B(n_9103),
.Y(n_19744)
);

INVx1_ASAP7_75t_L g19745 ( 
.A(n_19554),
.Y(n_19745)
);

OAI22xp5_ASAP7_75t_L g19746 ( 
.A1(n_19485),
.A2(n_9309),
.B1(n_9314),
.B2(n_9302),
.Y(n_19746)
);

NAND2xp5_ASAP7_75t_L g19747 ( 
.A(n_19491),
.B(n_9308),
.Y(n_19747)
);

AND2x2_ASAP7_75t_L g19748 ( 
.A(n_19469),
.B(n_9535),
.Y(n_19748)
);

AND2x2_ASAP7_75t_L g19749 ( 
.A(n_19496),
.B(n_19460),
.Y(n_19749)
);

INVx1_ASAP7_75t_L g19750 ( 
.A(n_19550),
.Y(n_19750)
);

NAND2xp5_ASAP7_75t_L g19751 ( 
.A(n_19510),
.B(n_9308),
.Y(n_19751)
);

AND3x1_ASAP7_75t_L g19752 ( 
.A(n_19470),
.B(n_8924),
.C(n_7259),
.Y(n_19752)
);

NOR2xp33_ASAP7_75t_L g19753 ( 
.A(n_19540),
.B(n_9311),
.Y(n_19753)
);

NAND2xp5_ASAP7_75t_SL g19754 ( 
.A(n_19436),
.B(n_9311),
.Y(n_19754)
);

INVx1_ASAP7_75t_L g19755 ( 
.A(n_19409),
.Y(n_19755)
);

XNOR2x2_ASAP7_75t_L g19756 ( 
.A(n_19566),
.B(n_9046),
.Y(n_19756)
);

INVx2_ASAP7_75t_L g19757 ( 
.A(n_19484),
.Y(n_19757)
);

XOR2xp5_ASAP7_75t_L g19758 ( 
.A(n_19608),
.B(n_8697),
.Y(n_19758)
);

XNOR2xp5_ASAP7_75t_L g19759 ( 
.A(n_19660),
.B(n_8697),
.Y(n_19759)
);

OAI32xp33_ASAP7_75t_L g19760 ( 
.A1(n_19456),
.A2(n_7725),
.A3(n_7773),
.B1(n_7758),
.B2(n_7694),
.Y(n_19760)
);

AND2x2_ASAP7_75t_L g19761 ( 
.A(n_19502),
.B(n_9535),
.Y(n_19761)
);

AND2x2_ASAP7_75t_L g19762 ( 
.A(n_19598),
.B(n_9535),
.Y(n_19762)
);

INVx2_ASAP7_75t_L g19763 ( 
.A(n_19561),
.Y(n_19763)
);

AND2x2_ASAP7_75t_L g19764 ( 
.A(n_19421),
.B(n_9576),
.Y(n_19764)
);

INVxp67_ASAP7_75t_L g19765 ( 
.A(n_19528),
.Y(n_19765)
);

AND2x2_ASAP7_75t_L g19766 ( 
.A(n_19480),
.B(n_9576),
.Y(n_19766)
);

AND2x2_ASAP7_75t_L g19767 ( 
.A(n_19433),
.B(n_19455),
.Y(n_19767)
);

XNOR2xp5_ASAP7_75t_L g19768 ( 
.A(n_19656),
.B(n_8697),
.Y(n_19768)
);

AOI22xp33_ASAP7_75t_L g19769 ( 
.A1(n_19603),
.A2(n_9311),
.B1(n_9351),
.B2(n_9323),
.Y(n_19769)
);

INVx1_ASAP7_75t_L g19770 ( 
.A(n_19475),
.Y(n_19770)
);

OR2x2_ASAP7_75t_L g19771 ( 
.A(n_19549),
.B(n_9292),
.Y(n_19771)
);

AOI21xp33_ASAP7_75t_L g19772 ( 
.A1(n_19617),
.A2(n_8690),
.B(n_9323),
.Y(n_19772)
);

OAI22xp5_ASAP7_75t_L g19773 ( 
.A1(n_19572),
.A2(n_9322),
.B1(n_9360),
.B2(n_9314),
.Y(n_19773)
);

NAND2xp5_ASAP7_75t_L g19774 ( 
.A(n_19662),
.B(n_19463),
.Y(n_19774)
);

NAND2xp5_ASAP7_75t_SL g19775 ( 
.A(n_19571),
.B(n_9323),
.Y(n_19775)
);

AND2x2_ASAP7_75t_L g19776 ( 
.A(n_19623),
.B(n_9576),
.Y(n_19776)
);

AND2x2_ASAP7_75t_L g19777 ( 
.A(n_19555),
.B(n_19511),
.Y(n_19777)
);

CKINVDCx20_ASAP7_75t_L g19778 ( 
.A(n_19643),
.Y(n_19778)
);

INVx1_ASAP7_75t_L g19779 ( 
.A(n_19486),
.Y(n_19779)
);

NAND2xp5_ASAP7_75t_L g19780 ( 
.A(n_19605),
.B(n_9323),
.Y(n_19780)
);

NAND2xp5_ASAP7_75t_L g19781 ( 
.A(n_19479),
.B(n_9351),
.Y(n_19781)
);

INVx1_ASAP7_75t_L g19782 ( 
.A(n_19477),
.Y(n_19782)
);

NAND2xp5_ASAP7_75t_L g19783 ( 
.A(n_19489),
.B(n_9351),
.Y(n_19783)
);

NAND2xp5_ASAP7_75t_L g19784 ( 
.A(n_19499),
.B(n_9351),
.Y(n_19784)
);

INVxp67_ASAP7_75t_L g19785 ( 
.A(n_19512),
.Y(n_19785)
);

INVx1_ASAP7_75t_SL g19786 ( 
.A(n_19649),
.Y(n_19786)
);

XOR2xp5_ASAP7_75t_L g19787 ( 
.A(n_19624),
.B(n_8697),
.Y(n_19787)
);

INVx1_ASAP7_75t_L g19788 ( 
.A(n_19658),
.Y(n_19788)
);

OAI21xp5_ASAP7_75t_L g19789 ( 
.A1(n_19522),
.A2(n_8432),
.B(n_9226),
.Y(n_19789)
);

XNOR2x1_ASAP7_75t_L g19790 ( 
.A(n_19659),
.B(n_8785),
.Y(n_19790)
);

OAI22xp5_ASAP7_75t_L g19791 ( 
.A1(n_19636),
.A2(n_9322),
.B1(n_9360),
.B2(n_9314),
.Y(n_19791)
);

OR2x2_ASAP7_75t_L g19792 ( 
.A(n_19664),
.B(n_9292),
.Y(n_19792)
);

AOI322xp5_ASAP7_75t_L g19793 ( 
.A1(n_19580),
.A2(n_9359),
.A3(n_9385),
.B1(n_9366),
.B2(n_9419),
.C1(n_9389),
.C2(n_9376),
.Y(n_19793)
);

INVx1_ASAP7_75t_L g19794 ( 
.A(n_19461),
.Y(n_19794)
);

INVx1_ASAP7_75t_L g19795 ( 
.A(n_19445),
.Y(n_19795)
);

INVx1_ASAP7_75t_L g19796 ( 
.A(n_19511),
.Y(n_19796)
);

INVx1_ASAP7_75t_L g19797 ( 
.A(n_19531),
.Y(n_19797)
);

NOR2x1_ASAP7_75t_L g19798 ( 
.A(n_19520),
.B(n_19525),
.Y(n_19798)
);

INVx1_ASAP7_75t_L g19799 ( 
.A(n_19432),
.Y(n_19799)
);

INVx1_ASAP7_75t_L g19800 ( 
.A(n_19503),
.Y(n_19800)
);

XNOR2x2_ASAP7_75t_L g19801 ( 
.A(n_19612),
.B(n_9046),
.Y(n_19801)
);

A2O1A1Ixp33_ASAP7_75t_L g19802 ( 
.A1(n_19611),
.A2(n_8539),
.B(n_9360),
.C(n_9322),
.Y(n_19802)
);

INVx1_ASAP7_75t_L g19803 ( 
.A(n_19507),
.Y(n_19803)
);

AND2x4_ASAP7_75t_L g19804 ( 
.A(n_19534),
.B(n_9359),
.Y(n_19804)
);

INVx1_ASAP7_75t_L g19805 ( 
.A(n_19518),
.Y(n_19805)
);

INVx1_ASAP7_75t_L g19806 ( 
.A(n_19439),
.Y(n_19806)
);

NAND2xp5_ASAP7_75t_L g19807 ( 
.A(n_19536),
.B(n_9359),
.Y(n_19807)
);

INVx1_ASAP7_75t_L g19808 ( 
.A(n_19523),
.Y(n_19808)
);

NOR3xp33_ASAP7_75t_SL g19809 ( 
.A(n_19537),
.B(n_7371),
.C(n_7444),
.Y(n_19809)
);

OR2x2_ASAP7_75t_L g19810 ( 
.A(n_19412),
.B(n_9292),
.Y(n_19810)
);

OAI21xp33_ASAP7_75t_L g19811 ( 
.A1(n_19595),
.A2(n_7219),
.B(n_7210),
.Y(n_19811)
);

INVxp67_ASAP7_75t_L g19812 ( 
.A(n_19596),
.Y(n_19812)
);

INVx2_ASAP7_75t_SL g19813 ( 
.A(n_19626),
.Y(n_19813)
);

AND2x2_ASAP7_75t_L g19814 ( 
.A(n_19417),
.B(n_9576),
.Y(n_19814)
);

INVx1_ASAP7_75t_L g19815 ( 
.A(n_19465),
.Y(n_19815)
);

HAxp5_ASAP7_75t_SL g19816 ( 
.A(n_19575),
.B(n_8720),
.CON(n_19816),
.SN(n_19816)
);

BUFx3_ASAP7_75t_L g19817 ( 
.A(n_19650),
.Y(n_19817)
);

NOR4xp25_ASAP7_75t_SL g19818 ( 
.A(n_19661),
.B(n_8045),
.C(n_8054),
.D(n_8028),
.Y(n_19818)
);

NAND2xp5_ASAP7_75t_L g19819 ( 
.A(n_19573),
.B(n_9359),
.Y(n_19819)
);

NAND2xp5_ASAP7_75t_L g19820 ( 
.A(n_19544),
.B(n_9366),
.Y(n_19820)
);

INVx1_ASAP7_75t_L g19821 ( 
.A(n_19500),
.Y(n_19821)
);

AND2x2_ASAP7_75t_L g19822 ( 
.A(n_19631),
.B(n_9576),
.Y(n_19822)
);

NAND2xp5_ASAP7_75t_L g19823 ( 
.A(n_19591),
.B(n_9366),
.Y(n_19823)
);

AND2x2_ASAP7_75t_L g19824 ( 
.A(n_19408),
.B(n_9576),
.Y(n_19824)
);

NOR2xp33_ASAP7_75t_L g19825 ( 
.A(n_19620),
.B(n_9366),
.Y(n_19825)
);

INVxp67_ASAP7_75t_L g19826 ( 
.A(n_19556),
.Y(n_19826)
);

NAND2xp5_ASAP7_75t_L g19827 ( 
.A(n_19471),
.B(n_19628),
.Y(n_19827)
);

INVx2_ASAP7_75t_L g19828 ( 
.A(n_19643),
.Y(n_19828)
);

INVx1_ASAP7_75t_L g19829 ( 
.A(n_19633),
.Y(n_19829)
);

INVx1_ASAP7_75t_L g19830 ( 
.A(n_19655),
.Y(n_19830)
);

HB1xp67_ASAP7_75t_L g19831 ( 
.A(n_19452),
.Y(n_19831)
);

OAI21xp5_ASAP7_75t_L g19832 ( 
.A1(n_19447),
.A2(n_8432),
.B(n_9226),
.Y(n_19832)
);

INVxp67_ASAP7_75t_L g19833 ( 
.A(n_19625),
.Y(n_19833)
);

AOI22xp33_ASAP7_75t_SL g19834 ( 
.A1(n_19634),
.A2(n_8773),
.B1(n_9330),
.B2(n_8711),
.Y(n_19834)
);

BUFx2_ASAP7_75t_L g19835 ( 
.A(n_19476),
.Y(n_19835)
);

BUFx2_ASAP7_75t_L g19836 ( 
.A(n_19450),
.Y(n_19836)
);

INVxp67_ASAP7_75t_L g19837 ( 
.A(n_19621),
.Y(n_19837)
);

CKINVDCx5p33_ASAP7_75t_R g19838 ( 
.A(n_19641),
.Y(n_19838)
);

OAI211xp5_ASAP7_75t_L g19839 ( 
.A1(n_19597),
.A2(n_7730),
.B(n_7164),
.C(n_7097),
.Y(n_19839)
);

OAI221xp5_ASAP7_75t_L g19840 ( 
.A1(n_19558),
.A2(n_8785),
.B1(n_8982),
.B2(n_8893),
.C(n_9103),
.Y(n_19840)
);

INVx1_ASAP7_75t_L g19841 ( 
.A(n_19648),
.Y(n_19841)
);

NAND2xp5_ASAP7_75t_L g19842 ( 
.A(n_19614),
.B(n_9376),
.Y(n_19842)
);

INVx1_ASAP7_75t_L g19843 ( 
.A(n_19647),
.Y(n_19843)
);

NOR3xp33_ASAP7_75t_SL g19844 ( 
.A(n_19562),
.B(n_7371),
.C(n_7444),
.Y(n_19844)
);

INVx1_ASAP7_75t_L g19845 ( 
.A(n_19506),
.Y(n_19845)
);

XNOR2x2_ASAP7_75t_L g19846 ( 
.A(n_19599),
.B(n_8641),
.Y(n_19846)
);

INVx1_ASAP7_75t_L g19847 ( 
.A(n_19574),
.Y(n_19847)
);

AND2x2_ASAP7_75t_L g19848 ( 
.A(n_19527),
.B(n_9576),
.Y(n_19848)
);

NAND2xp33_ASAP7_75t_SL g19849 ( 
.A(n_19630),
.B(n_7931),
.Y(n_19849)
);

INVx2_ASAP7_75t_L g19850 ( 
.A(n_19583),
.Y(n_19850)
);

NAND2xp33_ASAP7_75t_R g19851 ( 
.A(n_19638),
.B(n_8045),
.Y(n_19851)
);

INVx1_ASAP7_75t_L g19852 ( 
.A(n_19560),
.Y(n_19852)
);

INVx1_ASAP7_75t_L g19853 ( 
.A(n_19590),
.Y(n_19853)
);

INVx1_ASAP7_75t_L g19854 ( 
.A(n_19494),
.Y(n_19854)
);

NAND2xp5_ASAP7_75t_L g19855 ( 
.A(n_19444),
.B(n_9376),
.Y(n_19855)
);

BUFx2_ASAP7_75t_L g19856 ( 
.A(n_19657),
.Y(n_19856)
);

INVxp67_ASAP7_75t_SL g19857 ( 
.A(n_19493),
.Y(n_19857)
);

NOR4xp25_ASAP7_75t_SL g19858 ( 
.A(n_19569),
.B(n_8078),
.C(n_8101),
.D(n_8054),
.Y(n_19858)
);

NAND2xp5_ASAP7_75t_L g19859 ( 
.A(n_19478),
.B(n_9376),
.Y(n_19859)
);

OR2x6_ASAP7_75t_L g19860 ( 
.A(n_19487),
.B(n_9193),
.Y(n_19860)
);

OAI22xp5_ASAP7_75t_L g19861 ( 
.A1(n_19627),
.A2(n_9403),
.B1(n_9412),
.B2(n_9365),
.Y(n_19861)
);

INVx1_ASAP7_75t_L g19862 ( 
.A(n_19530),
.Y(n_19862)
);

BUFx3_ASAP7_75t_L g19863 ( 
.A(n_19593),
.Y(n_19863)
);

INVx1_ASAP7_75t_L g19864 ( 
.A(n_19565),
.Y(n_19864)
);

OAI22xp5_ASAP7_75t_L g19865 ( 
.A1(n_19547),
.A2(n_19616),
.B1(n_19610),
.B2(n_19418),
.Y(n_19865)
);

NOR2xp33_ASAP7_75t_L g19866 ( 
.A(n_19613),
.B(n_9385),
.Y(n_19866)
);

OAI311xp33_ASAP7_75t_L g19867 ( 
.A1(n_19585),
.A2(n_7219),
.A3(n_7210),
.B1(n_7567),
.C1(n_7560),
.Y(n_19867)
);

INVx1_ASAP7_75t_L g19868 ( 
.A(n_19588),
.Y(n_19868)
);

INVx1_ASAP7_75t_L g19869 ( 
.A(n_19609),
.Y(n_19869)
);

AOI211xp5_ASAP7_75t_L g19870 ( 
.A1(n_19632),
.A2(n_8539),
.B(n_7423),
.C(n_9226),
.Y(n_19870)
);

NAND2xp5_ASAP7_75t_L g19871 ( 
.A(n_19587),
.B(n_9385),
.Y(n_19871)
);

INVxp67_ASAP7_75t_L g19872 ( 
.A(n_19604),
.Y(n_19872)
);

OR2x2_ASAP7_75t_L g19873 ( 
.A(n_19577),
.B(n_9292),
.Y(n_19873)
);

NOR3xp33_ASAP7_75t_SL g19874 ( 
.A(n_19615),
.B(n_7470),
.C(n_7423),
.Y(n_19874)
);

OAI22xp5_ASAP7_75t_L g19875 ( 
.A1(n_19606),
.A2(n_9403),
.B1(n_9412),
.B2(n_9365),
.Y(n_19875)
);

AND2x2_ASAP7_75t_L g19876 ( 
.A(n_19644),
.B(n_9576),
.Y(n_19876)
);

AND2x2_ASAP7_75t_L g19877 ( 
.A(n_19552),
.B(n_9579),
.Y(n_19877)
);

INVx1_ASAP7_75t_L g19878 ( 
.A(n_19586),
.Y(n_19878)
);

INVx1_ASAP7_75t_L g19879 ( 
.A(n_19584),
.Y(n_19879)
);

NOR2xp33_ASAP7_75t_R g19880 ( 
.A(n_19589),
.B(n_19543),
.Y(n_19880)
);

INVx1_ASAP7_75t_L g19881 ( 
.A(n_19622),
.Y(n_19881)
);

O2A1O1Ixp33_ASAP7_75t_L g19882 ( 
.A1(n_19642),
.A2(n_9126),
.B(n_9138),
.C(n_9103),
.Y(n_19882)
);

AOI221x1_ASAP7_75t_SL g19883 ( 
.A1(n_19646),
.A2(n_7210),
.B1(n_7219),
.B2(n_9389),
.C(n_9385),
.Y(n_19883)
);

INVx1_ASAP7_75t_L g19884 ( 
.A(n_19563),
.Y(n_19884)
);

INVx1_ASAP7_75t_L g19885 ( 
.A(n_19645),
.Y(n_19885)
);

AND2x2_ASAP7_75t_L g19886 ( 
.A(n_19618),
.B(n_9579),
.Y(n_19886)
);

NAND2xp5_ASAP7_75t_L g19887 ( 
.A(n_19619),
.B(n_9389),
.Y(n_19887)
);

INVx1_ASAP7_75t_L g19888 ( 
.A(n_19619),
.Y(n_19888)
);

INVx1_ASAP7_75t_L g19889 ( 
.A(n_19553),
.Y(n_19889)
);

OR2x2_ASAP7_75t_L g19890 ( 
.A(n_19579),
.B(n_9292),
.Y(n_19890)
);

AOI211xp5_ASAP7_75t_SL g19891 ( 
.A1(n_19653),
.A2(n_19514),
.B(n_19524),
.C(n_19654),
.Y(n_19891)
);

NAND2xp33_ASAP7_75t_R g19892 ( 
.A(n_19601),
.B(n_8054),
.Y(n_19892)
);

OA22x2_ASAP7_75t_SL g19893 ( 
.A1(n_19711),
.A2(n_19640),
.B1(n_19592),
.B2(n_19602),
.Y(n_19893)
);

INVx1_ASAP7_75t_L g19894 ( 
.A(n_19715),
.Y(n_19894)
);

OAI21xp5_ASAP7_75t_L g19895 ( 
.A1(n_19681),
.A2(n_19629),
.B(n_19582),
.Y(n_19895)
);

INVx1_ASAP7_75t_L g19896 ( 
.A(n_19685),
.Y(n_19896)
);

AOI211x1_ASAP7_75t_L g19897 ( 
.A1(n_19673),
.A2(n_19672),
.B(n_19678),
.C(n_19687),
.Y(n_19897)
);

INVx1_ASAP7_75t_L g19898 ( 
.A(n_19709),
.Y(n_19898)
);

NAND2xp5_ASAP7_75t_L g19899 ( 
.A(n_19683),
.B(n_19637),
.Y(n_19899)
);

NAND3xp33_ASAP7_75t_L g19900 ( 
.A(n_19688),
.B(n_19488),
.C(n_19453),
.Y(n_19900)
);

NAND2xp5_ASAP7_75t_SL g19901 ( 
.A(n_19670),
.B(n_19669),
.Y(n_19901)
);

NOR4xp25_ASAP7_75t_L g19902 ( 
.A(n_19712),
.B(n_19532),
.C(n_19600),
.D(n_19594),
.Y(n_19902)
);

NAND3xp33_ASAP7_75t_L g19903 ( 
.A(n_19680),
.B(n_19578),
.C(n_19576),
.Y(n_19903)
);

NAND3xp33_ASAP7_75t_SL g19904 ( 
.A(n_19736),
.B(n_19521),
.C(n_19567),
.Y(n_19904)
);

AOI211x1_ASAP7_75t_SL g19905 ( 
.A1(n_19791),
.A2(n_19564),
.B(n_19635),
.C(n_19508),
.Y(n_19905)
);

AOI21xp5_ASAP7_75t_L g19906 ( 
.A1(n_19704),
.A2(n_19526),
.B(n_19513),
.Y(n_19906)
);

NAND2xp5_ASAP7_75t_SL g19907 ( 
.A(n_19684),
.B(n_19440),
.Y(n_19907)
);

AOI21xp5_ASAP7_75t_L g19908 ( 
.A1(n_19813),
.A2(n_19652),
.B(n_19651),
.Y(n_19908)
);

NAND2xp5_ASAP7_75t_SL g19909 ( 
.A(n_19705),
.B(n_19519),
.Y(n_19909)
);

NAND2xp5_ASAP7_75t_L g19910 ( 
.A(n_19786),
.B(n_9389),
.Y(n_19910)
);

INVx1_ASAP7_75t_L g19911 ( 
.A(n_19817),
.Y(n_19911)
);

AOI21xp5_ASAP7_75t_L g19912 ( 
.A1(n_19857),
.A2(n_9403),
.B(n_9365),
.Y(n_19912)
);

NOR2x1_ASAP7_75t_L g19913 ( 
.A(n_19708),
.B(n_9361),
.Y(n_19913)
);

AND2x2_ASAP7_75t_L g19914 ( 
.A(n_19757),
.B(n_9361),
.Y(n_19914)
);

NAND2xp5_ASAP7_75t_L g19915 ( 
.A(n_19830),
.B(n_9419),
.Y(n_19915)
);

NOR3xp33_ASAP7_75t_L g19916 ( 
.A(n_19692),
.B(n_7181),
.C(n_7144),
.Y(n_19916)
);

INVxp67_ASAP7_75t_L g19917 ( 
.A(n_19798),
.Y(n_19917)
);

AOI21xp5_ASAP7_75t_L g19918 ( 
.A1(n_19731),
.A2(n_9435),
.B(n_9412),
.Y(n_19918)
);

INVx1_ASAP7_75t_L g19919 ( 
.A(n_19728),
.Y(n_19919)
);

AOI211xp5_ASAP7_75t_L g19920 ( 
.A1(n_19829),
.A2(n_7423),
.B(n_8499),
.C(n_7470),
.Y(n_19920)
);

OA22x2_ASAP7_75t_L g19921 ( 
.A1(n_19724),
.A2(n_7078),
.B1(n_7158),
.B2(n_7097),
.Y(n_19921)
);

OAI211xp5_ASAP7_75t_L g19922 ( 
.A1(n_19812),
.A2(n_7730),
.B(n_7265),
.C(n_7294),
.Y(n_19922)
);

OAI22xp5_ASAP7_75t_L g19923 ( 
.A1(n_19693),
.A2(n_9441),
.B1(n_9447),
.B2(n_9435),
.Y(n_19923)
);

A2O1A1Ixp33_ASAP7_75t_SL g19924 ( 
.A1(n_19694),
.A2(n_9441),
.B(n_9447),
.C(n_9435),
.Y(n_19924)
);

OAI21xp33_ASAP7_75t_SL g19925 ( 
.A1(n_19860),
.A2(n_8739),
.B(n_8736),
.Y(n_19925)
);

OAI21xp33_ASAP7_75t_L g19926 ( 
.A1(n_19699),
.A2(n_7916),
.B(n_7910),
.Y(n_19926)
);

OAI211xp5_ASAP7_75t_SL g19927 ( 
.A1(n_19826),
.A2(n_7394),
.B(n_7730),
.C(n_9441),
.Y(n_19927)
);

NAND2xp5_ASAP7_75t_SL g19928 ( 
.A(n_19713),
.B(n_9419),
.Y(n_19928)
);

INVx1_ASAP7_75t_SL g19929 ( 
.A(n_19745),
.Y(n_19929)
);

AOI21xp33_ASAP7_75t_SL g19930 ( 
.A1(n_19696),
.A2(n_9138),
.B(n_9126),
.Y(n_19930)
);

INVx1_ASAP7_75t_L g19931 ( 
.A(n_19750),
.Y(n_19931)
);

INVx1_ASAP7_75t_L g19932 ( 
.A(n_19671),
.Y(n_19932)
);

AOI211x1_ASAP7_75t_L g19933 ( 
.A1(n_19775),
.A2(n_19819),
.B(n_19716),
.C(n_19730),
.Y(n_19933)
);

NOR2xp67_ASAP7_75t_L g19934 ( 
.A(n_19717),
.B(n_19722),
.Y(n_19934)
);

INVx1_ASAP7_75t_L g19935 ( 
.A(n_19676),
.Y(n_19935)
);

OAI21xp33_ASAP7_75t_L g19936 ( 
.A1(n_19695),
.A2(n_7960),
.B(n_7943),
.Y(n_19936)
);

AOI21xp5_ASAP7_75t_L g19937 ( 
.A1(n_19835),
.A2(n_9455),
.B(n_9447),
.Y(n_19937)
);

OAI21xp33_ASAP7_75t_L g19938 ( 
.A1(n_19765),
.A2(n_7963),
.B(n_7960),
.Y(n_19938)
);

INVx3_ASAP7_75t_L g19939 ( 
.A(n_19763),
.Y(n_19939)
);

NAND3xp33_ASAP7_75t_L g19940 ( 
.A(n_19837),
.B(n_19838),
.C(n_19833),
.Y(n_19940)
);

HB1xp67_ASAP7_75t_L g19941 ( 
.A(n_19706),
.Y(n_19941)
);

NOR2x1_ASAP7_75t_SL g19942 ( 
.A(n_19702),
.B(n_19796),
.Y(n_19942)
);

NOR3xp33_ASAP7_75t_L g19943 ( 
.A(n_19785),
.B(n_7217),
.C(n_7181),
.Y(n_19943)
);

AO22x2_ASAP7_75t_L g19944 ( 
.A1(n_19788),
.A2(n_9419),
.B1(n_9422),
.B2(n_9420),
.Y(n_19944)
);

NAND2xp5_ASAP7_75t_L g19945 ( 
.A(n_19749),
.B(n_19856),
.Y(n_19945)
);

OR2x2_ASAP7_75t_L g19946 ( 
.A(n_19686),
.B(n_19682),
.Y(n_19946)
);

INVx1_ASAP7_75t_L g19947 ( 
.A(n_19723),
.Y(n_19947)
);

AOI22xp5_ASAP7_75t_L g19948 ( 
.A1(n_19851),
.A2(n_9422),
.B1(n_9452),
.B2(n_9420),
.Y(n_19948)
);

NAND2xp5_ASAP7_75t_SL g19949 ( 
.A(n_19841),
.B(n_9420),
.Y(n_19949)
);

AOI221xp5_ASAP7_75t_L g19950 ( 
.A1(n_19849),
.A2(n_9469),
.B1(n_9480),
.B2(n_9456),
.C(n_9455),
.Y(n_19950)
);

AOI22xp33_ASAP7_75t_L g19951 ( 
.A1(n_19850),
.A2(n_9422),
.B1(n_9452),
.B2(n_9420),
.Y(n_19951)
);

NAND2xp5_ASAP7_75t_L g19952 ( 
.A(n_19675),
.B(n_9422),
.Y(n_19952)
);

NOR2x1_ASAP7_75t_SL g19953 ( 
.A(n_19737),
.B(n_9511),
.Y(n_19953)
);

AOI221xp5_ASAP7_75t_L g19954 ( 
.A1(n_19753),
.A2(n_9456),
.B1(n_9480),
.B2(n_9469),
.C(n_9455),
.Y(n_19954)
);

AOI22x1_ASAP7_75t_L g19955 ( 
.A1(n_19836),
.A2(n_7265),
.B1(n_7294),
.B2(n_7158),
.Y(n_19955)
);

INVx2_ASAP7_75t_L g19956 ( 
.A(n_19674),
.Y(n_19956)
);

AOI21xp5_ASAP7_75t_L g19957 ( 
.A1(n_19774),
.A2(n_9469),
.B(n_9456),
.Y(n_19957)
);

AOI21xp5_ASAP7_75t_L g19958 ( 
.A1(n_19739),
.A2(n_9481),
.B(n_9480),
.Y(n_19958)
);

NAND4xp25_ASAP7_75t_SL g19959 ( 
.A(n_19769),
.B(n_7933),
.C(n_7940),
.D(n_7911),
.Y(n_19959)
);

NOR2xp33_ASAP7_75t_L g19960 ( 
.A(n_19843),
.B(n_9452),
.Y(n_19960)
);

INVx1_ASAP7_75t_L g19961 ( 
.A(n_19831),
.Y(n_19961)
);

NAND2xp5_ASAP7_75t_L g19962 ( 
.A(n_19886),
.B(n_9452),
.Y(n_19962)
);

OAI21xp5_ASAP7_75t_L g19963 ( 
.A1(n_19827),
.A2(n_9493),
.B(n_9459),
.Y(n_19963)
);

NAND2xp5_ASAP7_75t_L g19964 ( 
.A(n_19767),
.B(n_19741),
.Y(n_19964)
);

OAI21xp5_ASAP7_75t_SL g19965 ( 
.A1(n_19777),
.A2(n_9138),
.B(n_9126),
.Y(n_19965)
);

NAND3xp33_ASAP7_75t_L g19966 ( 
.A(n_19854),
.B(n_9493),
.C(n_9459),
.Y(n_19966)
);

BUFx2_ASAP7_75t_L g19967 ( 
.A(n_19880),
.Y(n_19967)
);

AOI211xp5_ASAP7_75t_L g19968 ( 
.A1(n_19865),
.A2(n_8499),
.B(n_7470),
.C(n_7567),
.Y(n_19968)
);

AOI211xp5_ASAP7_75t_L g19969 ( 
.A1(n_19888),
.A2(n_7605),
.B(n_7627),
.C(n_7560),
.Y(n_19969)
);

INVx2_ASAP7_75t_SL g19970 ( 
.A(n_19790),
.Y(n_19970)
);

AOI211x1_ASAP7_75t_L g19971 ( 
.A1(n_19701),
.A2(n_9492),
.B(n_9502),
.C(n_9481),
.Y(n_19971)
);

INVx1_ASAP7_75t_L g19972 ( 
.A(n_19677),
.Y(n_19972)
);

NOR3xp33_ASAP7_75t_L g19973 ( 
.A(n_19755),
.B(n_7217),
.C(n_7181),
.Y(n_19973)
);

O2A1O1Ixp33_ASAP7_75t_L g19974 ( 
.A1(n_19872),
.A2(n_9147),
.B(n_9331),
.C(n_9138),
.Y(n_19974)
);

NOR2x1_ASAP7_75t_L g19975 ( 
.A(n_19806),
.B(n_19868),
.Y(n_19975)
);

INVx1_ASAP7_75t_L g19976 ( 
.A(n_19751),
.Y(n_19976)
);

HB1xp67_ASAP7_75t_L g19977 ( 
.A(n_19863),
.Y(n_19977)
);

OAI21xp33_ASAP7_75t_L g19978 ( 
.A1(n_19759),
.A2(n_19768),
.B(n_19679),
.Y(n_19978)
);

AOI211x1_ASAP7_75t_L g19979 ( 
.A1(n_19738),
.A2(n_9492),
.B(n_9502),
.C(n_9481),
.Y(n_19979)
);

NAND2xp5_ASAP7_75t_SL g19980 ( 
.A(n_19828),
.B(n_9459),
.Y(n_19980)
);

NOR3xp33_ASAP7_75t_SL g19981 ( 
.A(n_19852),
.B(n_7749),
.C(n_7688),
.Y(n_19981)
);

INVxp67_ASAP7_75t_SL g19982 ( 
.A(n_19799),
.Y(n_19982)
);

OA22x2_ASAP7_75t_L g19983 ( 
.A1(n_19710),
.A2(n_7375),
.B1(n_7398),
.B2(n_7352),
.Y(n_19983)
);

OAI211xp5_ASAP7_75t_SL g19984 ( 
.A1(n_19879),
.A2(n_9502),
.B(n_9516),
.C(n_9492),
.Y(n_19984)
);

NAND2xp5_ASAP7_75t_L g19985 ( 
.A(n_19848),
.B(n_9459),
.Y(n_19985)
);

AOI21xp5_ASAP7_75t_L g19986 ( 
.A1(n_19703),
.A2(n_9571),
.B(n_9516),
.Y(n_19986)
);

INVx2_ASAP7_75t_L g19987 ( 
.A(n_19674),
.Y(n_19987)
);

NAND2xp5_ASAP7_75t_L g19988 ( 
.A(n_19776),
.B(n_19782),
.Y(n_19988)
);

CKINVDCx20_ASAP7_75t_R g19989 ( 
.A(n_19726),
.Y(n_19989)
);

NOR3x1_ASAP7_75t_L g19990 ( 
.A(n_19845),
.B(n_8648),
.C(n_8641),
.Y(n_19990)
);

NAND2xp5_ASAP7_75t_SL g19991 ( 
.A(n_19808),
.B(n_9493),
.Y(n_19991)
);

NOR3x1_ASAP7_75t_L g19992 ( 
.A(n_19884),
.B(n_9026),
.C(n_9557),
.Y(n_19992)
);

NOR2x1_ASAP7_75t_L g19993 ( 
.A(n_19732),
.B(n_9511),
.Y(n_19993)
);

INVx1_ASAP7_75t_L g19994 ( 
.A(n_19718),
.Y(n_19994)
);

AOI21xp5_ASAP7_75t_L g19995 ( 
.A1(n_19690),
.A2(n_9571),
.B(n_9516),
.Y(n_19995)
);

AOI211x1_ASAP7_75t_SL g19996 ( 
.A1(n_19861),
.A2(n_9499),
.B(n_9506),
.C(n_9493),
.Y(n_19996)
);

AOI22xp5_ASAP7_75t_L g19997 ( 
.A1(n_19892),
.A2(n_9506),
.B1(n_9532),
.B2(n_9499),
.Y(n_19997)
);

OAI21xp33_ASAP7_75t_L g19998 ( 
.A1(n_19697),
.A2(n_7963),
.B(n_7960),
.Y(n_19998)
);

NAND2xp5_ASAP7_75t_L g19999 ( 
.A(n_19804),
.B(n_9499),
.Y(n_19999)
);

NAND2xp5_ASAP7_75t_L g20000 ( 
.A(n_19804),
.B(n_9499),
.Y(n_20000)
);

OAI22xp5_ASAP7_75t_L g20001 ( 
.A1(n_19860),
.A2(n_9571),
.B1(n_7259),
.B2(n_7244),
.Y(n_20001)
);

INVx1_ASAP7_75t_L g20002 ( 
.A(n_19729),
.Y(n_20002)
);

NAND3xp33_ASAP7_75t_SL g20003 ( 
.A(n_19795),
.B(n_8893),
.C(n_8785),
.Y(n_20003)
);

INVx1_ASAP7_75t_L g20004 ( 
.A(n_19780),
.Y(n_20004)
);

AND2x2_ASAP7_75t_L g20005 ( 
.A(n_19752),
.B(n_19844),
.Y(n_20005)
);

AOI22xp5_ASAP7_75t_L g20006 ( 
.A1(n_19824),
.A2(n_9532),
.B1(n_9568),
.B2(n_9506),
.Y(n_20006)
);

NAND2xp5_ASAP7_75t_L g20007 ( 
.A(n_19766),
.B(n_9506),
.Y(n_20007)
);

AOI21xp5_ASAP7_75t_L g20008 ( 
.A1(n_19714),
.A2(n_7500),
.B(n_7463),
.Y(n_20008)
);

AOI21xp5_ASAP7_75t_SL g20009 ( 
.A1(n_19869),
.A2(n_7259),
.B(n_7244),
.Y(n_20009)
);

AOI211x1_ASAP7_75t_L g20010 ( 
.A1(n_19754),
.A2(n_7605),
.B(n_7627),
.C(n_7560),
.Y(n_20010)
);

AOI211x1_ASAP7_75t_L g20011 ( 
.A1(n_19689),
.A2(n_7627),
.B(n_7605),
.C(n_7963),
.Y(n_20011)
);

AOI211x1_ASAP7_75t_L g20012 ( 
.A1(n_19773),
.A2(n_19698),
.B(n_19842),
.C(n_19747),
.Y(n_20012)
);

NAND4xp75_ASAP7_75t_L g20013 ( 
.A(n_19853),
.B(n_7970),
.C(n_7985),
.D(n_7968),
.Y(n_20013)
);

OAI22xp5_ASAP7_75t_L g20014 ( 
.A1(n_19818),
.A2(n_7244),
.B1(n_8773),
.B2(n_8711),
.Y(n_20014)
);

NAND5xp2_ASAP7_75t_SL g20015 ( 
.A(n_19778),
.B(n_7048),
.C(n_7058),
.D(n_7014),
.E(n_7002),
.Y(n_20015)
);

AOI22xp5_ASAP7_75t_L g20016 ( 
.A1(n_19876),
.A2(n_9568),
.B1(n_9532),
.B2(n_8773),
.Y(n_20016)
);

OAI211xp5_ASAP7_75t_SL g20017 ( 
.A1(n_19885),
.A2(n_7970),
.B(n_7985),
.C(n_7968),
.Y(n_20017)
);

AOI211x1_ASAP7_75t_L g20018 ( 
.A1(n_19772),
.A2(n_7970),
.B(n_7985),
.C(n_7968),
.Y(n_20018)
);

NAND2xp5_ASAP7_75t_L g20019 ( 
.A(n_19825),
.B(n_9532),
.Y(n_20019)
);

INVx1_ASAP7_75t_L g20020 ( 
.A(n_19823),
.Y(n_20020)
);

AOI21xp5_ASAP7_75t_L g20021 ( 
.A1(n_19779),
.A2(n_7500),
.B(n_7463),
.Y(n_20021)
);

NAND2xp5_ASAP7_75t_SL g20022 ( 
.A(n_19815),
.B(n_9568),
.Y(n_20022)
);

INVx1_ASAP7_75t_L g20023 ( 
.A(n_19727),
.Y(n_20023)
);

INVx1_ASAP7_75t_L g20024 ( 
.A(n_19719),
.Y(n_20024)
);

AND2x2_ASAP7_75t_L g20025 ( 
.A(n_19834),
.B(n_9238),
.Y(n_20025)
);

INVx1_ASAP7_75t_L g20026 ( 
.A(n_19784),
.Y(n_20026)
);

INVx1_ASAP7_75t_L g20027 ( 
.A(n_19807),
.Y(n_20027)
);

HB1xp67_ASAP7_75t_L g20028 ( 
.A(n_19794),
.Y(n_20028)
);

INVx1_ASAP7_75t_L g20029 ( 
.A(n_19770),
.Y(n_20029)
);

INVx1_ASAP7_75t_L g20030 ( 
.A(n_19797),
.Y(n_20030)
);

NAND3xp33_ASAP7_75t_L g20031 ( 
.A(n_19847),
.B(n_9568),
.C(n_7299),
.Y(n_20031)
);

NAND2xp5_ASAP7_75t_L g20032 ( 
.A(n_19758),
.B(n_7299),
.Y(n_20032)
);

AOI21xp5_ASAP7_75t_L g20033 ( 
.A1(n_19800),
.A2(n_7524),
.B(n_7463),
.Y(n_20033)
);

OR2x2_ASAP7_75t_L g20034 ( 
.A(n_19846),
.B(n_7352),
.Y(n_20034)
);

NOR3xp33_ASAP7_75t_L g20035 ( 
.A(n_19821),
.B(n_7217),
.C(n_7181),
.Y(n_20035)
);

AOI211xp5_ASAP7_75t_L g20036 ( 
.A1(n_19889),
.A2(n_8713),
.B(n_8725),
.C(n_7524),
.Y(n_20036)
);

NAND2xp5_ASAP7_75t_L g20037 ( 
.A(n_19764),
.B(n_7299),
.Y(n_20037)
);

NOR2xp33_ASAP7_75t_L g20038 ( 
.A(n_19803),
.B(n_8711),
.Y(n_20038)
);

NOR3xp33_ASAP7_75t_L g20039 ( 
.A(n_19805),
.B(n_7217),
.C(n_7181),
.Y(n_20039)
);

AND2x2_ASAP7_75t_L g20040 ( 
.A(n_19809),
.B(n_9238),
.Y(n_20040)
);

NOR3xp33_ASAP7_75t_L g20041 ( 
.A(n_19878),
.B(n_7217),
.C(n_7181),
.Y(n_20041)
);

INVx1_ASAP7_75t_L g20042 ( 
.A(n_19781),
.Y(n_20042)
);

NAND2xp5_ASAP7_75t_L g20043 ( 
.A(n_19787),
.B(n_7299),
.Y(n_20043)
);

NAND2xp5_ASAP7_75t_L g20044 ( 
.A(n_19866),
.B(n_19864),
.Y(n_20044)
);

AOI21xp5_ASAP7_75t_L g20045 ( 
.A1(n_19891),
.A2(n_7996),
.B(n_7988),
.Y(n_20045)
);

AOI211xp5_ASAP7_75t_L g20046 ( 
.A1(n_19862),
.A2(n_8713),
.B(n_8725),
.C(n_9026),
.Y(n_20046)
);

OAI21xp5_ASAP7_75t_L g20047 ( 
.A1(n_19881),
.A2(n_8547),
.B(n_8543),
.Y(n_20047)
);

AO22x2_ASAP7_75t_L g20048 ( 
.A1(n_19783),
.A2(n_7983),
.B1(n_7996),
.B2(n_7988),
.Y(n_20048)
);

AOI21xp5_ASAP7_75t_L g20049 ( 
.A1(n_19887),
.A2(n_7996),
.B(n_7988),
.Y(n_20049)
);

INVx1_ASAP7_75t_L g20050 ( 
.A(n_19810),
.Y(n_20050)
);

INVxp67_ASAP7_75t_L g20051 ( 
.A(n_19720),
.Y(n_20051)
);

AOI21xp5_ASAP7_75t_L g20052 ( 
.A1(n_19855),
.A2(n_8000),
.B(n_7998),
.Y(n_20052)
);

AOI211xp5_ASAP7_75t_L g20053 ( 
.A1(n_19725),
.A2(n_8713),
.B(n_8725),
.C(n_9026),
.Y(n_20053)
);

INVx1_ASAP7_75t_L g20054 ( 
.A(n_19801),
.Y(n_20054)
);

INVx1_ASAP7_75t_L g20055 ( 
.A(n_19873),
.Y(n_20055)
);

NAND2xp33_ASAP7_75t_L g20056 ( 
.A(n_19874),
.B(n_7375),
.Y(n_20056)
);

INVx1_ASAP7_75t_L g20057 ( 
.A(n_19756),
.Y(n_20057)
);

OA22x2_ASAP7_75t_L g20058 ( 
.A1(n_19871),
.A2(n_7398),
.B1(n_7733),
.B2(n_7711),
.Y(n_20058)
);

INVx1_ASAP7_75t_L g20059 ( 
.A(n_19820),
.Y(n_20059)
);

AOI22x1_ASAP7_75t_L g20060 ( 
.A1(n_19822),
.A2(n_8101),
.B1(n_8107),
.B2(n_8078),
.Y(n_20060)
);

NAND2xp5_ASAP7_75t_SL g20061 ( 
.A(n_19771),
.B(n_9238),
.Y(n_20061)
);

INVx1_ASAP7_75t_L g20062 ( 
.A(n_19859),
.Y(n_20062)
);

AOI21xp5_ASAP7_75t_L g20063 ( 
.A1(n_19740),
.A2(n_8000),
.B(n_7998),
.Y(n_20063)
);

AOI22xp33_ASAP7_75t_SL g20064 ( 
.A1(n_19877),
.A2(n_9330),
.B1(n_9485),
.B2(n_8773),
.Y(n_20064)
);

AOI211x1_ASAP7_75t_SL g20065 ( 
.A1(n_19721),
.A2(n_8000),
.B(n_8026),
.C(n_7998),
.Y(n_20065)
);

INVx1_ASAP7_75t_L g20066 ( 
.A(n_19733),
.Y(n_20066)
);

AOI21xp5_ASAP7_75t_L g20067 ( 
.A1(n_19760),
.A2(n_8026),
.B(n_8127),
.Y(n_20067)
);

OAI21xp5_ASAP7_75t_L g20068 ( 
.A1(n_19735),
.A2(n_8547),
.B(n_8543),
.Y(n_20068)
);

NAND2xp5_ASAP7_75t_L g20069 ( 
.A(n_19814),
.B(n_7299),
.Y(n_20069)
);

NAND2xp5_ASAP7_75t_L g20070 ( 
.A(n_19707),
.B(n_7299),
.Y(n_20070)
);

INVx1_ASAP7_75t_L g20071 ( 
.A(n_19700),
.Y(n_20071)
);

AND2x2_ASAP7_75t_L g20072 ( 
.A(n_19858),
.B(n_9238),
.Y(n_20072)
);

NOR3xp33_ASAP7_75t_L g20073 ( 
.A(n_19839),
.B(n_7300),
.C(n_7217),
.Y(n_20073)
);

INVx2_ASAP7_75t_L g20074 ( 
.A(n_19792),
.Y(n_20074)
);

AOI22xp5_ASAP7_75t_L g20075 ( 
.A1(n_19748),
.A2(n_9330),
.B1(n_9485),
.B2(n_8773),
.Y(n_20075)
);

INVx1_ASAP7_75t_L g20076 ( 
.A(n_19890),
.Y(n_20076)
);

AOI21xp5_ASAP7_75t_L g20077 ( 
.A1(n_19762),
.A2(n_8026),
.B(n_8127),
.Y(n_20077)
);

AOI21xp33_ASAP7_75t_SL g20078 ( 
.A1(n_19742),
.A2(n_9331),
.B(n_9147),
.Y(n_20078)
);

NAND2xp5_ASAP7_75t_L g20079 ( 
.A(n_19883),
.B(n_7299),
.Y(n_20079)
);

AOI21xp5_ASAP7_75t_L g20080 ( 
.A1(n_19743),
.A2(n_8127),
.B(n_7073),
.Y(n_20080)
);

INVx1_ASAP7_75t_L g20081 ( 
.A(n_19761),
.Y(n_20081)
);

OAI211xp5_ASAP7_75t_L g20082 ( 
.A1(n_19811),
.A2(n_7752),
.B(n_7783),
.C(n_7733),
.Y(n_20082)
);

NOR2xp33_ASAP7_75t_L g20083 ( 
.A(n_19691),
.B(n_8773),
.Y(n_20083)
);

NAND2xp5_ASAP7_75t_L g20084 ( 
.A(n_19875),
.B(n_7496),
.Y(n_20084)
);

AND2x2_ASAP7_75t_L g20085 ( 
.A(n_19744),
.B(n_9240),
.Y(n_20085)
);

AOI21xp5_ASAP7_75t_L g20086 ( 
.A1(n_19882),
.A2(n_7073),
.B(n_8061),
.Y(n_20086)
);

NAND2xp5_ASAP7_75t_SL g20087 ( 
.A(n_19793),
.B(n_9240),
.Y(n_20087)
);

NAND2xp5_ASAP7_75t_L g20088 ( 
.A(n_19746),
.B(n_7496),
.Y(n_20088)
);

INVx1_ASAP7_75t_SL g20089 ( 
.A(n_19816),
.Y(n_20089)
);

INVx1_ASAP7_75t_SL g20090 ( 
.A(n_19789),
.Y(n_20090)
);

AOI32xp33_ASAP7_75t_L g20091 ( 
.A1(n_19896),
.A2(n_19840),
.A3(n_19870),
.B1(n_19867),
.B2(n_19802),
.Y(n_20091)
);

NAND2xp5_ASAP7_75t_L g20092 ( 
.A(n_19917),
.B(n_19832),
.Y(n_20092)
);

AOI21xp33_ASAP7_75t_L g20093 ( 
.A1(n_19894),
.A2(n_19734),
.B(n_7073),
.Y(n_20093)
);

INVx1_ASAP7_75t_L g20094 ( 
.A(n_19942),
.Y(n_20094)
);

INVxp67_ASAP7_75t_SL g20095 ( 
.A(n_19934),
.Y(n_20095)
);

OAI22xp5_ASAP7_75t_SL g20096 ( 
.A1(n_19897),
.A2(n_9485),
.B1(n_9330),
.B2(n_7694),
.Y(n_20096)
);

O2A1O1Ixp33_ASAP7_75t_L g20097 ( 
.A1(n_20057),
.A2(n_9331),
.B(n_9337),
.C(n_9147),
.Y(n_20097)
);

AOI221xp5_ASAP7_75t_L g20098 ( 
.A1(n_19902),
.A2(n_6943),
.B1(n_6957),
.B2(n_6937),
.C(n_6936),
.Y(n_20098)
);

AND2x2_ASAP7_75t_L g20099 ( 
.A(n_20072),
.B(n_9240),
.Y(n_20099)
);

INVx1_ASAP7_75t_L g20100 ( 
.A(n_19939),
.Y(n_20100)
);

BUFx2_ASAP7_75t_L g20101 ( 
.A(n_19939),
.Y(n_20101)
);

NAND2xp5_ASAP7_75t_L g20102 ( 
.A(n_19911),
.B(n_7496),
.Y(n_20102)
);

INVx1_ASAP7_75t_L g20103 ( 
.A(n_19945),
.Y(n_20103)
);

AOI22xp5_ASAP7_75t_L g20104 ( 
.A1(n_19982),
.A2(n_9330),
.B1(n_9485),
.B2(n_7073),
.Y(n_20104)
);

NAND2xp5_ASAP7_75t_SL g20105 ( 
.A(n_19929),
.B(n_9240),
.Y(n_20105)
);

INVx1_ASAP7_75t_L g20106 ( 
.A(n_20028),
.Y(n_20106)
);

OAI21xp5_ASAP7_75t_L g20107 ( 
.A1(n_19940),
.A2(n_19906),
.B(n_19975),
.Y(n_20107)
);

AOI221xp5_ASAP7_75t_L g20108 ( 
.A1(n_20054),
.A2(n_6943),
.B1(n_6957),
.B2(n_6937),
.C(n_6936),
.Y(n_20108)
);

NAND2xp33_ASAP7_75t_SL g20109 ( 
.A(n_19898),
.B(n_7931),
.Y(n_20109)
);

AOI221xp5_ASAP7_75t_L g20110 ( 
.A1(n_19967),
.A2(n_6943),
.B1(n_6957),
.B2(n_6937),
.C(n_6936),
.Y(n_20110)
);

NAND2xp5_ASAP7_75t_L g20111 ( 
.A(n_19941),
.B(n_7496),
.Y(n_20111)
);

OAI211xp5_ASAP7_75t_L g20112 ( 
.A1(n_19933),
.A2(n_7783),
.B(n_7752),
.C(n_7018),
.Y(n_20112)
);

O2A1O1Ixp33_ASAP7_75t_L g20113 ( 
.A1(n_19964),
.A2(n_9472),
.B(n_9331),
.C(n_9337),
.Y(n_20113)
);

NOR2x1_ASAP7_75t_L g20114 ( 
.A(n_19961),
.B(n_7725),
.Y(n_20114)
);

AOI221xp5_ASAP7_75t_L g20115 ( 
.A1(n_19904),
.A2(n_6966),
.B1(n_6970),
.B2(n_6964),
.C(n_6960),
.Y(n_20115)
);

A2O1A1Ixp33_ASAP7_75t_SL g20116 ( 
.A1(n_19919),
.A2(n_7150),
.B(n_7156),
.C(n_7141),
.Y(n_20116)
);

AOI21xp33_ASAP7_75t_L g20117 ( 
.A1(n_19977),
.A2(n_7073),
.B(n_7983),
.Y(n_20117)
);

INVx1_ASAP7_75t_L g20118 ( 
.A(n_20034),
.Y(n_20118)
);

NAND2xp5_ASAP7_75t_L g20119 ( 
.A(n_19931),
.B(n_7496),
.Y(n_20119)
);

INVx1_ASAP7_75t_L g20120 ( 
.A(n_19913),
.Y(n_20120)
);

OAI21xp33_ASAP7_75t_L g20121 ( 
.A1(n_20038),
.A2(n_7758),
.B(n_7725),
.Y(n_20121)
);

INVx1_ASAP7_75t_L g20122 ( 
.A(n_19989),
.Y(n_20122)
);

INVxp33_ASAP7_75t_SL g20123 ( 
.A(n_19899),
.Y(n_20123)
);

OAI311xp33_ASAP7_75t_L g20124 ( 
.A1(n_19895),
.A2(n_7410),
.A3(n_7983),
.B1(n_7425),
.C1(n_7414),
.Y(n_20124)
);

INVx1_ASAP7_75t_L g20125 ( 
.A(n_19993),
.Y(n_20125)
);

NOR2xp33_ASAP7_75t_L g20126 ( 
.A(n_20029),
.B(n_9330),
.Y(n_20126)
);

OAI22xp33_ASAP7_75t_L g20127 ( 
.A1(n_19970),
.A2(n_9485),
.B1(n_7725),
.B2(n_7773),
.Y(n_20127)
);

INVx1_ASAP7_75t_L g20128 ( 
.A(n_20005),
.Y(n_20128)
);

INVx1_ASAP7_75t_L g20129 ( 
.A(n_19956),
.Y(n_20129)
);

A2O1A1Ixp33_ASAP7_75t_L g20130 ( 
.A1(n_19978),
.A2(n_9128),
.B(n_9130),
.C(n_9124),
.Y(n_20130)
);

AND2x2_ASAP7_75t_L g20131 ( 
.A(n_20040),
.B(n_9240),
.Y(n_20131)
);

NAND2xp5_ASAP7_75t_L g20132 ( 
.A(n_19905),
.B(n_7496),
.Y(n_20132)
);

AOI22xp5_ASAP7_75t_L g20133 ( 
.A1(n_20089),
.A2(n_9485),
.B1(n_7073),
.B2(n_8027),
.Y(n_20133)
);

NAND5xp2_ASAP7_75t_L g20134 ( 
.A(n_20030),
.B(n_8893),
.C(n_8982),
.D(n_8785),
.E(n_9147),
.Y(n_20134)
);

INVx1_ASAP7_75t_L g20135 ( 
.A(n_19987),
.Y(n_20135)
);

AOI22xp33_ASAP7_75t_L g20136 ( 
.A1(n_20074),
.A2(n_9358),
.B1(n_7773),
.B2(n_7787),
.Y(n_20136)
);

OAI22xp5_ASAP7_75t_L g20137 ( 
.A1(n_19935),
.A2(n_7773),
.B1(n_7787),
.B2(n_7758),
.Y(n_20137)
);

INVx1_ASAP7_75t_L g20138 ( 
.A(n_19914),
.Y(n_20138)
);

INVx1_ASAP7_75t_L g20139 ( 
.A(n_19910),
.Y(n_20139)
);

XNOR2x2_ASAP7_75t_L g20140 ( 
.A(n_19901),
.B(n_9559),
.Y(n_20140)
);

AOI21xp33_ASAP7_75t_SL g20141 ( 
.A1(n_19988),
.A2(n_9337),
.B(n_9331),
.Y(n_20141)
);

OAI21xp33_ASAP7_75t_L g20142 ( 
.A1(n_19909),
.A2(n_7787),
.B(n_7758),
.Y(n_20142)
);

AOI21xp33_ASAP7_75t_L g20143 ( 
.A1(n_19946),
.A2(n_7983),
.B(n_8333),
.Y(n_20143)
);

INVx1_ASAP7_75t_L g20144 ( 
.A(n_19915),
.Y(n_20144)
);

OAI21xp5_ASAP7_75t_L g20145 ( 
.A1(n_19903),
.A2(n_8432),
.B(n_8543),
.Y(n_20145)
);

INVx1_ASAP7_75t_L g20146 ( 
.A(n_20056),
.Y(n_20146)
);

NAND5xp2_ASAP7_75t_L g20147 ( 
.A(n_19908),
.B(n_8893),
.C(n_8982),
.D(n_8785),
.E(n_9337),
.Y(n_20147)
);

CKINVDCx20_ASAP7_75t_R g20148 ( 
.A(n_19907),
.Y(n_20148)
);

INVx1_ASAP7_75t_L g20149 ( 
.A(n_20044),
.Y(n_20149)
);

AND2x2_ASAP7_75t_L g20150 ( 
.A(n_20025),
.B(n_9240),
.Y(n_20150)
);

HB1xp67_ASAP7_75t_L g20151 ( 
.A(n_19932),
.Y(n_20151)
);

AOI22xp5_ASAP7_75t_L g20152 ( 
.A1(n_20066),
.A2(n_7839),
.B1(n_8080),
.B2(n_7841),
.Y(n_20152)
);

AOI21xp33_ASAP7_75t_L g20153 ( 
.A1(n_20050),
.A2(n_8333),
.B(n_7425),
.Y(n_20153)
);

INVx2_ASAP7_75t_L g20154 ( 
.A(n_19893),
.Y(n_20154)
);

O2A1O1Ixp33_ASAP7_75t_L g20155 ( 
.A1(n_20051),
.A2(n_9448),
.B(n_9472),
.C(n_9337),
.Y(n_20155)
);

INVx1_ASAP7_75t_L g20156 ( 
.A(n_20012),
.Y(n_20156)
);

INVx1_ASAP7_75t_L g20157 ( 
.A(n_19949),
.Y(n_20157)
);

INVx1_ASAP7_75t_SL g20158 ( 
.A(n_20090),
.Y(n_20158)
);

OAI211xp5_ASAP7_75t_SL g20159 ( 
.A1(n_20055),
.A2(n_7911),
.B(n_7940),
.C(n_7933),
.Y(n_20159)
);

BUFx2_ASAP7_75t_L g20160 ( 
.A(n_19972),
.Y(n_20160)
);

AOI221xp5_ASAP7_75t_L g20161 ( 
.A1(n_19900),
.A2(n_6966),
.B1(n_6970),
.B2(n_6964),
.C(n_6960),
.Y(n_20161)
);

AOI211xp5_ASAP7_75t_L g20162 ( 
.A1(n_20081),
.A2(n_7688),
.B(n_8390),
.C(n_8388),
.Y(n_20162)
);

INVxp67_ASAP7_75t_SL g20163 ( 
.A(n_20004),
.Y(n_20163)
);

NOR3xp33_ASAP7_75t_L g20164 ( 
.A(n_20020),
.B(n_7300),
.C(n_8015),
.Y(n_20164)
);

INVx1_ASAP7_75t_L g20165 ( 
.A(n_20062),
.Y(n_20165)
);

AOI22xp5_ASAP7_75t_L g20166 ( 
.A1(n_20023),
.A2(n_7839),
.B1(n_8080),
.B2(n_7841),
.Y(n_20166)
);

OAI311xp33_ASAP7_75t_L g20167 ( 
.A1(n_20076),
.A2(n_7410),
.A3(n_7425),
.B1(n_7414),
.C1(n_7921),
.Y(n_20167)
);

INVx1_ASAP7_75t_L g20168 ( 
.A(n_20024),
.Y(n_20168)
);

AOI221xp5_ASAP7_75t_L g20169 ( 
.A1(n_20071),
.A2(n_6966),
.B1(n_6970),
.B2(n_6964),
.C(n_6960),
.Y(n_20169)
);

AOI322xp5_ASAP7_75t_L g20170 ( 
.A1(n_19960),
.A2(n_8015),
.A3(n_8001),
.B1(n_7378),
.B2(n_7278),
.C1(n_7284),
.C2(n_7273),
.Y(n_20170)
);

AOI22xp5_ASAP7_75t_L g20171 ( 
.A1(n_20083),
.A2(n_7787),
.B1(n_7841),
.B2(n_7839),
.Y(n_20171)
);

NOR2xp33_ASAP7_75t_L g20172 ( 
.A(n_19947),
.B(n_8893),
.Y(n_20172)
);

OAI211xp5_ASAP7_75t_SL g20173 ( 
.A1(n_19994),
.A2(n_7911),
.B(n_7940),
.C(n_7933),
.Y(n_20173)
);

AOI322xp5_ASAP7_75t_L g20174 ( 
.A1(n_20061),
.A2(n_8001),
.A3(n_7378),
.B1(n_7278),
.B2(n_7284),
.C1(n_7273),
.C2(n_7410),
.Y(n_20174)
);

AOI211xp5_ASAP7_75t_L g20175 ( 
.A1(n_19976),
.A2(n_7688),
.B(n_8388),
.C(n_7923),
.Y(n_20175)
);

AND2x2_ASAP7_75t_L g20176 ( 
.A(n_20085),
.B(n_7486),
.Y(n_20176)
);

AOI21xp5_ASAP7_75t_L g20177 ( 
.A1(n_20026),
.A2(n_8095),
.B(n_8061),
.Y(n_20177)
);

INVx1_ASAP7_75t_L g20178 ( 
.A(n_20027),
.Y(n_20178)
);

OA21x2_ASAP7_75t_L g20179 ( 
.A1(n_20042),
.A2(n_8762),
.B(n_8754),
.Y(n_20179)
);

INVxp67_ASAP7_75t_SL g20180 ( 
.A(n_20002),
.Y(n_20180)
);

NOR2x1_ASAP7_75t_L g20181 ( 
.A(n_20059),
.B(n_7839),
.Y(n_20181)
);

O2A1O1Ixp33_ASAP7_75t_L g20182 ( 
.A1(n_19928),
.A2(n_9448),
.B(n_9472),
.C(n_8982),
.Y(n_20182)
);

INVx1_ASAP7_75t_L g20183 ( 
.A(n_19962),
.Y(n_20183)
);

INVx1_ASAP7_75t_L g20184 ( 
.A(n_20022),
.Y(n_20184)
);

A2O1A1Ixp33_ASAP7_75t_L g20185 ( 
.A1(n_20016),
.A2(n_9128),
.B(n_9130),
.C(n_9124),
.Y(n_20185)
);

NOR3xp33_ASAP7_75t_L g20186 ( 
.A(n_19980),
.B(n_7300),
.C(n_8679),
.Y(n_20186)
);

INVx2_ASAP7_75t_SL g20187 ( 
.A(n_19991),
.Y(n_20187)
);

NAND2xp5_ASAP7_75t_L g20188 ( 
.A(n_20006),
.B(n_7496),
.Y(n_20188)
);

AOI31xp33_ASAP7_75t_SL g20189 ( 
.A1(n_19916),
.A2(n_7619),
.A3(n_7623),
.B(n_7599),
.Y(n_20189)
);

NOR3x1_ASAP7_75t_L g20190 ( 
.A(n_19952),
.B(n_9128),
.C(n_9124),
.Y(n_20190)
);

AOI211xp5_ASAP7_75t_SL g20191 ( 
.A1(n_19973),
.A2(n_7749),
.B(n_7923),
.C(n_7279),
.Y(n_20191)
);

OA22x2_ASAP7_75t_L g20192 ( 
.A1(n_19997),
.A2(n_9133),
.B1(n_9150),
.B2(n_9130),
.Y(n_20192)
);

AOI21xp5_ASAP7_75t_L g20193 ( 
.A1(n_20087),
.A2(n_8095),
.B(n_8061),
.Y(n_20193)
);

INVx2_ASAP7_75t_L g20194 ( 
.A(n_19944),
.Y(n_20194)
);

AOI21xp5_ASAP7_75t_L g20195 ( 
.A1(n_19953),
.A2(n_8097),
.B(n_8095),
.Y(n_20195)
);

INVx1_ASAP7_75t_SL g20196 ( 
.A(n_20007),
.Y(n_20196)
);

AOI22xp5_ASAP7_75t_L g20197 ( 
.A1(n_19948),
.A2(n_7841),
.B1(n_8027),
.B2(n_7950),
.Y(n_20197)
);

NAND2xp5_ASAP7_75t_L g20198 ( 
.A(n_19985),
.B(n_7496),
.Y(n_20198)
);

OR2x2_ASAP7_75t_L g20199 ( 
.A(n_20079),
.B(n_9579),
.Y(n_20199)
);

OAI221xp5_ASAP7_75t_L g20200 ( 
.A1(n_20060),
.A2(n_19943),
.B1(n_20064),
.B2(n_20039),
.C(n_20035),
.Y(n_20200)
);

AOI221x1_ASAP7_75t_L g20201 ( 
.A1(n_19957),
.A2(n_7749),
.B1(n_7923),
.B2(n_7150),
.C(n_7267),
.Y(n_20201)
);

O2A1O1Ixp33_ASAP7_75t_L g20202 ( 
.A1(n_19924),
.A2(n_9448),
.B(n_9472),
.C(n_8982),
.Y(n_20202)
);

AOI22xp33_ASAP7_75t_L g20203 ( 
.A1(n_20037),
.A2(n_9358),
.B1(n_8027),
.B2(n_8064),
.Y(n_20203)
);

NAND4xp75_ASAP7_75t_L g20204 ( 
.A(n_20018),
.B(n_7414),
.C(n_7494),
.D(n_7341),
.Y(n_20204)
);

INVx1_ASAP7_75t_L g20205 ( 
.A(n_19983),
.Y(n_20205)
);

INVx2_ASAP7_75t_SL g20206 ( 
.A(n_20019),
.Y(n_20206)
);

INVx1_ASAP7_75t_L g20207 ( 
.A(n_19996),
.Y(n_20207)
);

OA211x2_ASAP7_75t_L g20208 ( 
.A1(n_19959),
.A2(n_7541),
.B(n_7532),
.C(n_8097),
.Y(n_20208)
);

INVx1_ASAP7_75t_SL g20209 ( 
.A(n_19999),
.Y(n_20209)
);

OAI22xp5_ASAP7_75t_L g20210 ( 
.A1(n_20075),
.A2(n_8027),
.B1(n_8064),
.B2(n_7950),
.Y(n_20210)
);

AOI221xp5_ASAP7_75t_L g20211 ( 
.A1(n_20078),
.A2(n_6978),
.B1(n_6982),
.B2(n_6973),
.C(n_6971),
.Y(n_20211)
);

INVxp67_ASAP7_75t_SL g20212 ( 
.A(n_20000),
.Y(n_20212)
);

AOI22xp5_ASAP7_75t_L g20213 ( 
.A1(n_20043),
.A2(n_8064),
.B1(n_8080),
.B2(n_7950),
.Y(n_20213)
);

NOR2x1_ASAP7_75t_L g20214 ( 
.A(n_19966),
.B(n_7950),
.Y(n_20214)
);

AOI322xp5_ASAP7_75t_L g20215 ( 
.A1(n_19926),
.A2(n_7378),
.A3(n_7278),
.B1(n_7284),
.B2(n_7273),
.C1(n_8059),
.C2(n_7962),
.Y(n_20215)
);

INVxp67_ASAP7_75t_L g20216 ( 
.A(n_20084),
.Y(n_20216)
);

OAI211xp5_ASAP7_75t_L g20217 ( 
.A1(n_19955),
.A2(n_7018),
.B(n_7025),
.C(n_8078),
.Y(n_20217)
);

OAI22xp5_ASAP7_75t_SL g20218 ( 
.A1(n_19971),
.A2(n_8064),
.B1(n_8080),
.B2(n_9448),
.Y(n_20218)
);

AOI21xp5_ASAP7_75t_L g20219 ( 
.A1(n_20080),
.A2(n_8121),
.B(n_8097),
.Y(n_20219)
);

INVx2_ASAP7_75t_L g20220 ( 
.A(n_19944),
.Y(n_20220)
);

INVx2_ASAP7_75t_L g20221 ( 
.A(n_20058),
.Y(n_20221)
);

OAI22xp5_ASAP7_75t_SL g20222 ( 
.A1(n_20088),
.A2(n_9448),
.B1(n_9472),
.B2(n_7004),
.Y(n_20222)
);

INVx2_ASAP7_75t_L g20223 ( 
.A(n_19921),
.Y(n_20223)
);

OAI21xp33_ASAP7_75t_L g20224 ( 
.A1(n_19981),
.A2(n_8059),
.B(n_7962),
.Y(n_20224)
);

INVx2_ASAP7_75t_L g20225 ( 
.A(n_20048),
.Y(n_20225)
);

AOI22xp5_ASAP7_75t_L g20226 ( 
.A1(n_20032),
.A2(n_9358),
.B1(n_7278),
.B2(n_7284),
.Y(n_20226)
);

XOR2x2_ASAP7_75t_L g20227 ( 
.A(n_20041),
.B(n_7300),
.Y(n_20227)
);

OAI21xp33_ASAP7_75t_SL g20228 ( 
.A1(n_19950),
.A2(n_20009),
.B(n_19937),
.Y(n_20228)
);

XNOR2x1_ASAP7_75t_L g20229 ( 
.A(n_20014),
.B(n_8679),
.Y(n_20229)
);

OAI21xp5_ASAP7_75t_L g20230 ( 
.A1(n_20069),
.A2(n_8560),
.B(n_8547),
.Y(n_20230)
);

AOI22xp5_ASAP7_75t_L g20231 ( 
.A1(n_20070),
.A2(n_9358),
.B1(n_7378),
.B2(n_7273),
.Y(n_20231)
);

AOI22xp33_ASAP7_75t_L g20232 ( 
.A1(n_19963),
.A2(n_20031),
.B1(n_20073),
.B2(n_20047),
.Y(n_20232)
);

O2A1O1Ixp33_ASAP7_75t_L g20233 ( 
.A1(n_20045),
.A2(n_7931),
.B(n_8048),
.C(n_7939),
.Y(n_20233)
);

XNOR2xp5_ASAP7_75t_L g20234 ( 
.A(n_20065),
.B(n_9146),
.Y(n_20234)
);

INVxp67_ASAP7_75t_L g20235 ( 
.A(n_19958),
.Y(n_20235)
);

CKINVDCx20_ASAP7_75t_R g20236 ( 
.A(n_19938),
.Y(n_20236)
);

XNOR2xp5_ASAP7_75t_L g20237 ( 
.A(n_19979),
.B(n_9146),
.Y(n_20237)
);

NAND2xp33_ASAP7_75t_R g20238 ( 
.A(n_19912),
.B(n_8101),
.Y(n_20238)
);

INVx1_ASAP7_75t_L g20239 ( 
.A(n_20082),
.Y(n_20239)
);

NAND2xp5_ASAP7_75t_SL g20240 ( 
.A(n_19968),
.B(n_6976),
.Y(n_20240)
);

INVx1_ASAP7_75t_L g20241 ( 
.A(n_19918),
.Y(n_20241)
);

AOI222xp33_ASAP7_75t_L g20242 ( 
.A1(n_19927),
.A2(n_8720),
.B1(n_9144),
.B2(n_9387),
.C1(n_8388),
.C2(n_8369),
.Y(n_20242)
);

AOI22xp5_ASAP7_75t_L g20243 ( 
.A1(n_20086),
.A2(n_9358),
.B1(n_7300),
.B2(n_8954),
.Y(n_20243)
);

OA21x2_ASAP7_75t_L g20244 ( 
.A1(n_19995),
.A2(n_8762),
.B(n_8754),
.Y(n_20244)
);

OAI21xp5_ASAP7_75t_SL g20245 ( 
.A1(n_19922),
.A2(n_7040),
.B(n_6976),
.Y(n_20245)
);

INVx2_ASAP7_75t_L g20246 ( 
.A(n_20048),
.Y(n_20246)
);

AOI221xp5_ASAP7_75t_L g20247 ( 
.A1(n_20015),
.A2(n_6978),
.B1(n_6982),
.B2(n_6973),
.C(n_6971),
.Y(n_20247)
);

AOI211xp5_ASAP7_75t_SL g20248 ( 
.A1(n_20033),
.A2(n_7279),
.B(n_7852),
.C(n_7828),
.Y(n_20248)
);

NOR2xp33_ASAP7_75t_R g20249 ( 
.A(n_20094),
.B(n_20003),
.Y(n_20249)
);

NAND2xp5_ASAP7_75t_L g20250 ( 
.A(n_20101),
.B(n_20077),
.Y(n_20250)
);

XNOR2xp5_ASAP7_75t_L g20251 ( 
.A(n_20148),
.B(n_20010),
.Y(n_20251)
);

AOI221xp5_ASAP7_75t_L g20252 ( 
.A1(n_20095),
.A2(n_19984),
.B1(n_20001),
.B2(n_19986),
.C(n_20011),
.Y(n_20252)
);

NAND3xp33_ASAP7_75t_SL g20253 ( 
.A(n_20158),
.B(n_19920),
.C(n_20068),
.Y(n_20253)
);

NAND4xp25_ASAP7_75t_SL g20254 ( 
.A(n_20122),
.B(n_20021),
.C(n_20067),
.D(n_20052),
.Y(n_20254)
);

O2A1O1Ixp33_ASAP7_75t_L g20255 ( 
.A1(n_20107),
.A2(n_19930),
.B(n_19965),
.C(n_19925),
.Y(n_20255)
);

OAI211xp5_ASAP7_75t_L g20256 ( 
.A1(n_20106),
.A2(n_19936),
.B(n_19951),
.C(n_20063),
.Y(n_20256)
);

NAND4xp75_ASAP7_75t_L g20257 ( 
.A(n_20100),
.B(n_19992),
.C(n_19990),
.D(n_20008),
.Y(n_20257)
);

AOI21x1_ASAP7_75t_L g20258 ( 
.A1(n_20103),
.A2(n_20049),
.B(n_19923),
.Y(n_20258)
);

AOI21xp33_ASAP7_75t_L g20259 ( 
.A1(n_20151),
.A2(n_20180),
.B(n_20163),
.Y(n_20259)
);

AOI222xp33_ASAP7_75t_L g20260 ( 
.A1(n_20156),
.A2(n_19954),
.B1(n_19998),
.B2(n_20017),
.C1(n_20013),
.C2(n_20036),
.Y(n_20260)
);

HB1xp67_ASAP7_75t_L g20261 ( 
.A(n_20154),
.Y(n_20261)
);

NOR2x1_ASAP7_75t_L g20262 ( 
.A(n_20120),
.B(n_19974),
.Y(n_20262)
);

NAND4xp25_ASAP7_75t_L g20263 ( 
.A(n_20160),
.B(n_19969),
.C(n_20053),
.D(n_20046),
.Y(n_20263)
);

AND2x4_ASAP7_75t_L g20264 ( 
.A(n_20114),
.B(n_7486),
.Y(n_20264)
);

OAI32xp33_ASAP7_75t_L g20265 ( 
.A1(n_20123),
.A2(n_20092),
.A3(n_20118),
.B1(n_20149),
.B2(n_20128),
.Y(n_20265)
);

OAI21x1_ASAP7_75t_L g20266 ( 
.A1(n_20221),
.A2(n_9053),
.B(n_9050),
.Y(n_20266)
);

OAI211xp5_ASAP7_75t_L g20267 ( 
.A1(n_20129),
.A2(n_7300),
.B(n_8109),
.C(n_8107),
.Y(n_20267)
);

NOR3xp33_ASAP7_75t_L g20268 ( 
.A(n_20135),
.B(n_9150),
.C(n_9133),
.Y(n_20268)
);

NAND3xp33_ASAP7_75t_L g20269 ( 
.A(n_20165),
.B(n_7915),
.C(n_7568),
.Y(n_20269)
);

NOR3xp33_ASAP7_75t_L g20270 ( 
.A(n_20168),
.B(n_20178),
.C(n_20183),
.Y(n_20270)
);

AOI221xp5_ASAP7_75t_L g20271 ( 
.A1(n_20207),
.A2(n_20125),
.B1(n_20205),
.B2(n_20093),
.C(n_20132),
.Y(n_20271)
);

AOI22xp5_ASAP7_75t_L g20272 ( 
.A1(n_20126),
.A2(n_9358),
.B1(n_8954),
.B2(n_8997),
.Y(n_20272)
);

OAI221xp5_ASAP7_75t_L g20273 ( 
.A1(n_20091),
.A2(n_7939),
.B1(n_8079),
.B2(n_8048),
.C(n_7931),
.Y(n_20273)
);

OAI211xp5_ASAP7_75t_SL g20274 ( 
.A1(n_20216),
.A2(n_8059),
.B(n_8083),
.C(n_7962),
.Y(n_20274)
);

A2O1A1Ixp33_ASAP7_75t_L g20275 ( 
.A1(n_20223),
.A2(n_9150),
.B(n_9152),
.C(n_9133),
.Y(n_20275)
);

AOI21xp33_ASAP7_75t_SL g20276 ( 
.A1(n_20187),
.A2(n_8684),
.B(n_8679),
.Y(n_20276)
);

AOI21xp5_ASAP7_75t_L g20277 ( 
.A1(n_20212),
.A2(n_20220),
.B(n_20194),
.Y(n_20277)
);

OR2x2_ASAP7_75t_L g20278 ( 
.A(n_20105),
.B(n_9579),
.Y(n_20278)
);

AOI221x1_ASAP7_75t_L g20279 ( 
.A1(n_20138),
.A2(n_20146),
.B1(n_20157),
.B2(n_20184),
.C(n_20241),
.Y(n_20279)
);

AND2x2_ASAP7_75t_L g20280 ( 
.A(n_20099),
.B(n_9152),
.Y(n_20280)
);

NOR2xp33_ASAP7_75t_R g20281 ( 
.A(n_20139),
.B(n_7216),
.Y(n_20281)
);

NAND2xp5_ASAP7_75t_SL g20282 ( 
.A(n_20196),
.B(n_6976),
.Y(n_20282)
);

AOI22xp5_ASAP7_75t_L g20283 ( 
.A1(n_20181),
.A2(n_9358),
.B1(n_8954),
.B2(n_8997),
.Y(n_20283)
);

INVx1_ASAP7_75t_L g20284 ( 
.A(n_20225),
.Y(n_20284)
);

NOR2xp33_ASAP7_75t_L g20285 ( 
.A(n_20209),
.B(n_7372),
.Y(n_20285)
);

AOI22xp5_ASAP7_75t_L g20286 ( 
.A1(n_20236),
.A2(n_9358),
.B1(n_8954),
.B2(n_8997),
.Y(n_20286)
);

AOI22xp33_ASAP7_75t_L g20287 ( 
.A1(n_20206),
.A2(n_6973),
.B1(n_6978),
.B2(n_6971),
.Y(n_20287)
);

AOI211xp5_ASAP7_75t_SL g20288 ( 
.A1(n_20235),
.A2(n_7279),
.B(n_7852),
.C(n_7828),
.Y(n_20288)
);

NAND2xp5_ASAP7_75t_SL g20289 ( 
.A(n_20239),
.B(n_20246),
.Y(n_20289)
);

OAI211xp5_ASAP7_75t_L g20290 ( 
.A1(n_20144),
.A2(n_8109),
.B(n_8117),
.C(n_8107),
.Y(n_20290)
);

NOR2xp33_ASAP7_75t_L g20291 ( 
.A(n_20111),
.B(n_7380),
.Y(n_20291)
);

OAI221xp5_ASAP7_75t_L g20292 ( 
.A1(n_20232),
.A2(n_8048),
.B1(n_8079),
.B2(n_7939),
.C(n_7004),
.Y(n_20292)
);

OAI321xp33_ASAP7_75t_L g20293 ( 
.A1(n_20200),
.A2(n_9275),
.A3(n_9146),
.B1(n_8962),
.B2(n_8803),
.C(n_8876),
.Y(n_20293)
);

AOI211xp5_ASAP7_75t_L g20294 ( 
.A1(n_20228),
.A2(n_20115),
.B(n_20098),
.C(n_20245),
.Y(n_20294)
);

AOI211xp5_ASAP7_75t_L g20295 ( 
.A1(n_20222),
.A2(n_9050),
.B(n_9053),
.C(n_8560),
.Y(n_20295)
);

AOI221x1_ASAP7_75t_L g20296 ( 
.A1(n_20109),
.A2(n_7156),
.B1(n_7276),
.B2(n_7267),
.C(n_7173),
.Y(n_20296)
);

AND2x4_ASAP7_75t_L g20297 ( 
.A(n_20131),
.B(n_20150),
.Y(n_20297)
);

OAI21xp5_ASAP7_75t_L g20298 ( 
.A1(n_20119),
.A2(n_8560),
.B(n_8369),
.Y(n_20298)
);

AOI221xp5_ASAP7_75t_L g20299 ( 
.A1(n_20224),
.A2(n_6989),
.B1(n_6992),
.B2(n_6987),
.C(n_6982),
.Y(n_20299)
);

A2O1A1Ixp33_ASAP7_75t_L g20300 ( 
.A1(n_20108),
.A2(n_20142),
.B(n_20199),
.C(n_20172),
.Y(n_20300)
);

INVx2_ASAP7_75t_L g20301 ( 
.A(n_20140),
.Y(n_20301)
);

NAND2x1_ASAP7_75t_SL g20302 ( 
.A(n_20214),
.B(n_7939),
.Y(n_20302)
);

NAND4xp75_ASAP7_75t_L g20303 ( 
.A(n_20208),
.B(n_7494),
.C(n_7844),
.D(n_7341),
.Y(n_20303)
);

AOI22xp5_ASAP7_75t_L g20304 ( 
.A1(n_20176),
.A2(n_8954),
.B1(n_8997),
.B2(n_8672),
.Y(n_20304)
);

NOR2xp33_ASAP7_75t_R g20305 ( 
.A(n_20238),
.B(n_7216),
.Y(n_20305)
);

AOI221xp5_ASAP7_75t_L g20306 ( 
.A1(n_20102),
.A2(n_6992),
.B1(n_7016),
.B2(n_6989),
.C(n_6987),
.Y(n_20306)
);

NOR3x1_ASAP7_75t_L g20307 ( 
.A(n_20198),
.B(n_9156),
.C(n_9152),
.Y(n_20307)
);

AOI22xp5_ASAP7_75t_L g20308 ( 
.A1(n_20240),
.A2(n_8954),
.B1(n_8997),
.B2(n_8672),
.Y(n_20308)
);

NAND2xp5_ASAP7_75t_L g20309 ( 
.A(n_20227),
.B(n_7496),
.Y(n_20309)
);

A2O1A1Ixp33_ASAP7_75t_L g20310 ( 
.A1(n_20097),
.A2(n_9161),
.B(n_9162),
.C(n_9156),
.Y(n_20310)
);

AND2x2_ASAP7_75t_L g20311 ( 
.A(n_20234),
.B(n_9156),
.Y(n_20311)
);

OAI322xp33_ASAP7_75t_L g20312 ( 
.A1(n_20096),
.A2(n_7741),
.A3(n_7599),
.B1(n_7842),
.B2(n_7623),
.C1(n_7619),
.C2(n_8003),
.Y(n_20312)
);

OAI322xp33_ASAP7_75t_L g20313 ( 
.A1(n_20188),
.A2(n_7741),
.A3(n_7599),
.B1(n_7842),
.B2(n_7623),
.C1(n_7619),
.C2(n_8003),
.Y(n_20313)
);

O2A1O1Ixp5_ASAP7_75t_L g20314 ( 
.A1(n_20124),
.A2(n_7025),
.B(n_7018),
.C(n_7532),
.Y(n_20314)
);

OR2x2_ASAP7_75t_L g20315 ( 
.A(n_20229),
.B(n_9579),
.Y(n_20315)
);

AOI211xp5_ASAP7_75t_SL g20316 ( 
.A1(n_20217),
.A2(n_7852),
.B(n_7863),
.C(n_7828),
.Y(n_20316)
);

NOR2xp33_ASAP7_75t_L g20317 ( 
.A(n_20237),
.B(n_7380),
.Y(n_20317)
);

AO221x1_ASAP7_75t_L g20318 ( 
.A1(n_20127),
.A2(n_7918),
.B1(n_7957),
.B2(n_7889),
.C(n_7834),
.Y(n_20318)
);

O2A1O1Ixp33_ASAP7_75t_L g20319 ( 
.A1(n_20189),
.A2(n_7939),
.B(n_8079),
.C(n_8048),
.Y(n_20319)
);

AOI221xp5_ASAP7_75t_L g20320 ( 
.A1(n_20143),
.A2(n_6992),
.B1(n_7016),
.B2(n_6989),
.C(n_6987),
.Y(n_20320)
);

AND3x1_ASAP7_75t_L g20321 ( 
.A(n_20121),
.B(n_8124),
.C(n_8121),
.Y(n_20321)
);

OAI22xp5_ASAP7_75t_L g20322 ( 
.A1(n_20152),
.A2(n_20213),
.B1(n_20133),
.B2(n_20166),
.Y(n_20322)
);

NAND2xp5_ASAP7_75t_L g20323 ( 
.A(n_20112),
.B(n_7496),
.Y(n_20323)
);

OAI321xp33_ASAP7_75t_L g20324 ( 
.A1(n_20159),
.A2(n_9275),
.A3(n_9146),
.B1(n_8962),
.B2(n_8803),
.C(n_8876),
.Y(n_20324)
);

AOI322xp5_ASAP7_75t_L g20325 ( 
.A1(n_20153),
.A2(n_8121),
.A3(n_8124),
.B1(n_7632),
.B2(n_7645),
.C1(n_7577),
.C2(n_8115),
.Y(n_20325)
);

AOI21xp5_ASAP7_75t_SL g20326 ( 
.A1(n_20233),
.A2(n_7025),
.B(n_7018),
.Y(n_20326)
);

NOR2xp33_ASAP7_75t_L g20327 ( 
.A(n_20117),
.B(n_7380),
.Y(n_20327)
);

AOI222xp33_ASAP7_75t_L g20328 ( 
.A1(n_20145),
.A2(n_9144),
.B1(n_9387),
.B2(n_8720),
.C1(n_6976),
.C2(n_7071),
.Y(n_20328)
);

XNOR2xp5_ASAP7_75t_L g20329 ( 
.A(n_20137),
.B(n_9146),
.Y(n_20329)
);

AOI22xp5_ASAP7_75t_L g20330 ( 
.A1(n_20218),
.A2(n_8954),
.B1(n_8997),
.B2(n_8672),
.Y(n_20330)
);

NAND2xp5_ASAP7_75t_L g20331 ( 
.A(n_20161),
.B(n_7257),
.Y(n_20331)
);

BUFx2_ASAP7_75t_L g20332 ( 
.A(n_20230),
.Y(n_20332)
);

AOI211xp5_ASAP7_75t_L g20333 ( 
.A1(n_20173),
.A2(n_9053),
.B(n_9050),
.C(n_8583),
.Y(n_20333)
);

INVx1_ASAP7_75t_L g20334 ( 
.A(n_20195),
.Y(n_20334)
);

INVx1_ASAP7_75t_L g20335 ( 
.A(n_20243),
.Y(n_20335)
);

OAI211xp5_ASAP7_75t_L g20336 ( 
.A1(n_20201),
.A2(n_8117),
.B(n_8122),
.C(n_8109),
.Y(n_20336)
);

NOR4xp25_ASAP7_75t_L g20337 ( 
.A(n_20167),
.B(n_8115),
.C(n_8083),
.D(n_7811),
.Y(n_20337)
);

AOI211xp5_ASAP7_75t_L g20338 ( 
.A1(n_20141),
.A2(n_8583),
.B(n_8567),
.C(n_9063),
.Y(n_20338)
);

NAND4xp25_ASAP7_75t_L g20339 ( 
.A(n_20191),
.B(n_8122),
.C(n_8117),
.D(n_8115),
.Y(n_20339)
);

INVx1_ASAP7_75t_L g20340 ( 
.A(n_20177),
.Y(n_20340)
);

OA211x2_ASAP7_75t_L g20341 ( 
.A1(n_20211),
.A2(n_7541),
.B(n_7532),
.C(n_8124),
.Y(n_20341)
);

OAI221xp5_ASAP7_75t_SL g20342 ( 
.A1(n_20104),
.A2(n_8083),
.B1(n_7008),
.B2(n_7811),
.C(n_7833),
.Y(n_20342)
);

OAI221xp5_ASAP7_75t_L g20343 ( 
.A1(n_20116),
.A2(n_8048),
.B1(n_8079),
.B2(n_7004),
.C(n_7018),
.Y(n_20343)
);

XOR2xp5_ASAP7_75t_SL g20344 ( 
.A(n_20171),
.B(n_7599),
.Y(n_20344)
);

AOI222xp33_ASAP7_75t_L g20345 ( 
.A1(n_20169),
.A2(n_9387),
.B1(n_9144),
.B2(n_6976),
.C1(n_7071),
.C2(n_7098),
.Y(n_20345)
);

A2O1A1Ixp33_ASAP7_75t_L g20346 ( 
.A1(n_20248),
.A2(n_9162),
.B(n_9161),
.C(n_8762),
.Y(n_20346)
);

OR2x2_ASAP7_75t_L g20347 ( 
.A(n_20193),
.B(n_9579),
.Y(n_20347)
);

NAND4xp25_ASAP7_75t_SL g20348 ( 
.A(n_20175),
.B(n_20202),
.C(n_20226),
.D(n_20197),
.Y(n_20348)
);

OAI221xp5_ASAP7_75t_SL g20349 ( 
.A1(n_20203),
.A2(n_7008),
.B1(n_7811),
.B2(n_7833),
.C(n_7799),
.Y(n_20349)
);

OAI31xp33_ASAP7_75t_L g20350 ( 
.A1(n_20186),
.A2(n_8019),
.A3(n_6947),
.B(n_6994),
.Y(n_20350)
);

NAND2xp5_ASAP7_75t_L g20351 ( 
.A(n_20162),
.B(n_7257),
.Y(n_20351)
);

NOR3xp33_ASAP7_75t_L g20352 ( 
.A(n_20210),
.B(n_9162),
.C(n_9161),
.Y(n_20352)
);

NAND2xp5_ASAP7_75t_L g20353 ( 
.A(n_20231),
.B(n_20110),
.Y(n_20353)
);

OAI22xp5_ASAP7_75t_L g20354 ( 
.A1(n_20136),
.A2(n_7215),
.B1(n_7249),
.B2(n_7222),
.Y(n_20354)
);

AOI21xp33_ASAP7_75t_L g20355 ( 
.A1(n_20113),
.A2(n_9146),
.B(n_8803),
.Y(n_20355)
);

AOI221xp5_ASAP7_75t_L g20356 ( 
.A1(n_20164),
.A2(n_7024),
.B1(n_7021),
.B2(n_7016),
.C(n_7521),
.Y(n_20356)
);

NOR3xp33_ASAP7_75t_L g20357 ( 
.A(n_20147),
.B(n_8684),
.C(n_6411),
.Y(n_20357)
);

NAND3xp33_ASAP7_75t_L g20358 ( 
.A(n_20174),
.B(n_7915),
.C(n_7568),
.Y(n_20358)
);

NAND4xp25_ASAP7_75t_L g20359 ( 
.A(n_20242),
.B(n_20134),
.C(n_20155),
.D(n_20182),
.Y(n_20359)
);

NAND4xp25_ASAP7_75t_L g20360 ( 
.A(n_20215),
.B(n_8122),
.C(n_7025),
.D(n_7018),
.Y(n_20360)
);

OAI321xp33_ASAP7_75t_L g20361 ( 
.A1(n_20219),
.A2(n_9275),
.A3(n_9146),
.B1(n_8962),
.B2(n_8803),
.C(n_8876),
.Y(n_20361)
);

NOR3xp33_ASAP7_75t_SL g20362 ( 
.A(n_20130),
.B(n_7873),
.C(n_7863),
.Y(n_20362)
);

AOI211xp5_ASAP7_75t_L g20363 ( 
.A1(n_20247),
.A2(n_8567),
.B(n_8583),
.C(n_9063),
.Y(n_20363)
);

AOI211xp5_ASAP7_75t_L g20364 ( 
.A1(n_20185),
.A2(n_8567),
.B(n_9066),
.C(n_9063),
.Y(n_20364)
);

AOI222xp33_ASAP7_75t_L g20365 ( 
.A1(n_20190),
.A2(n_9387),
.B1(n_9144),
.B2(n_6976),
.C1(n_7071),
.C2(n_7098),
.Y(n_20365)
);

AOI21xp33_ASAP7_75t_L g20366 ( 
.A1(n_20192),
.A2(n_8803),
.B(n_8700),
.Y(n_20366)
);

NAND2xp33_ASAP7_75t_R g20367 ( 
.A(n_20244),
.B(n_7534),
.Y(n_20367)
);

AOI31xp33_ASAP7_75t_L g20368 ( 
.A1(n_20170),
.A2(n_7623),
.A3(n_7741),
.B(n_7619),
.Y(n_20368)
);

NAND3xp33_ASAP7_75t_L g20369 ( 
.A(n_20244),
.B(n_20179),
.C(n_20204),
.Y(n_20369)
);

AOI221xp5_ASAP7_75t_L g20370 ( 
.A1(n_20179),
.A2(n_7024),
.B1(n_7021),
.B2(n_7523),
.C(n_7521),
.Y(n_20370)
);

AOI22xp5_ASAP7_75t_L g20371 ( 
.A1(n_20095),
.A2(n_8954),
.B1(n_8997),
.B2(n_8672),
.Y(n_20371)
);

NOR3xp33_ASAP7_75t_SL g20372 ( 
.A(n_20107),
.B(n_7873),
.C(n_7863),
.Y(n_20372)
);

NOR2xp33_ASAP7_75t_R g20373 ( 
.A(n_20094),
.B(n_7216),
.Y(n_20373)
);

NAND4xp25_ASAP7_75t_SL g20374 ( 
.A(n_20094),
.B(n_7833),
.C(n_7888),
.D(n_7799),
.Y(n_20374)
);

OAI211xp5_ASAP7_75t_L g20375 ( 
.A1(n_20107),
.A2(n_7025),
.B(n_7771),
.C(n_7765),
.Y(n_20375)
);

OAI211xp5_ASAP7_75t_SL g20376 ( 
.A1(n_20107),
.A2(n_7581),
.B(n_7697),
.C(n_7565),
.Y(n_20376)
);

OAI221xp5_ASAP7_75t_L g20377 ( 
.A1(n_20107),
.A2(n_8079),
.B1(n_7004),
.B2(n_7025),
.C(n_7541),
.Y(n_20377)
);

NOR2xp33_ASAP7_75t_R g20378 ( 
.A(n_20094),
.B(n_7216),
.Y(n_20378)
);

AOI211xp5_ASAP7_75t_L g20379 ( 
.A1(n_20107),
.A2(n_9066),
.B(n_9068),
.C(n_9067),
.Y(n_20379)
);

BUFx2_ASAP7_75t_L g20380 ( 
.A(n_20101),
.Y(n_20380)
);

AOI221xp5_ASAP7_75t_L g20381 ( 
.A1(n_20095),
.A2(n_7024),
.B1(n_7021),
.B2(n_7523),
.C(n_7521),
.Y(n_20381)
);

AOI22xp33_ASAP7_75t_L g20382 ( 
.A1(n_20101),
.A2(n_7040),
.B1(n_7071),
.B2(n_6976),
.Y(n_20382)
);

O2A1O1Ixp33_ASAP7_75t_L g20383 ( 
.A1(n_20094),
.A2(n_7004),
.B(n_7873),
.C(n_6775),
.Y(n_20383)
);

INVx1_ASAP7_75t_L g20384 ( 
.A(n_20101),
.Y(n_20384)
);

AOI221xp5_ASAP7_75t_L g20385 ( 
.A1(n_20095),
.A2(n_7547),
.B1(n_7556),
.B2(n_7529),
.C(n_7523),
.Y(n_20385)
);

NAND2xp33_ASAP7_75t_R g20386 ( 
.A(n_20094),
.B(n_7535),
.Y(n_20386)
);

NAND4xp25_ASAP7_75t_L g20387 ( 
.A(n_20107),
.B(n_7844),
.C(n_7494),
.D(n_7581),
.Y(n_20387)
);

OAI211xp5_ASAP7_75t_SL g20388 ( 
.A1(n_20107),
.A2(n_7581),
.B(n_7697),
.C(n_7565),
.Y(n_20388)
);

OAI21xp5_ASAP7_75t_L g20389 ( 
.A1(n_20095),
.A2(n_8369),
.B(n_8595),
.Y(n_20389)
);

AOI222xp33_ASAP7_75t_L g20390 ( 
.A1(n_20101),
.A2(n_9387),
.B1(n_9144),
.B2(n_6976),
.C1(n_7071),
.C2(n_7098),
.Y(n_20390)
);

AOI211xp5_ASAP7_75t_L g20391 ( 
.A1(n_20107),
.A2(n_9067),
.B(n_9068),
.C(n_9066),
.Y(n_20391)
);

OAI21xp5_ASAP7_75t_L g20392 ( 
.A1(n_20095),
.A2(n_8595),
.B(n_8684),
.Y(n_20392)
);

OAI221xp5_ASAP7_75t_SL g20393 ( 
.A1(n_20094),
.A2(n_7008),
.B1(n_7888),
.B2(n_7901),
.C(n_7799),
.Y(n_20393)
);

OAI221xp5_ASAP7_75t_L g20394 ( 
.A1(n_20107),
.A2(n_7040),
.B1(n_7098),
.B2(n_7071),
.C(n_6976),
.Y(n_20394)
);

AOI221xp5_ASAP7_75t_L g20395 ( 
.A1(n_20095),
.A2(n_7556),
.B1(n_7557),
.B2(n_7547),
.C(n_7529),
.Y(n_20395)
);

INVx1_ASAP7_75t_L g20396 ( 
.A(n_20101),
.Y(n_20396)
);

NOR2xp33_ASAP7_75t_L g20397 ( 
.A(n_20380),
.B(n_7921),
.Y(n_20397)
);

NOR2x1_ASAP7_75t_L g20398 ( 
.A(n_20384),
.B(n_7104),
.Y(n_20398)
);

NOR4xp25_ASAP7_75t_L g20399 ( 
.A(n_20259),
.B(n_7901),
.C(n_7888),
.D(n_7697),
.Y(n_20399)
);

NOR2x1_ASAP7_75t_L g20400 ( 
.A(n_20396),
.B(n_7104),
.Y(n_20400)
);

NOR3xp33_ASAP7_75t_L g20401 ( 
.A(n_20265),
.B(n_6411),
.C(n_6405),
.Y(n_20401)
);

NAND2xp5_ASAP7_75t_L g20402 ( 
.A(n_20261),
.B(n_9292),
.Y(n_20402)
);

OAI21xp5_ASAP7_75t_L g20403 ( 
.A1(n_20277),
.A2(n_8368),
.B(n_8595),
.Y(n_20403)
);

NAND2xp5_ASAP7_75t_L g20404 ( 
.A(n_20297),
.B(n_9292),
.Y(n_20404)
);

NAND4xp75_ASAP7_75t_L g20405 ( 
.A(n_20279),
.B(n_7844),
.C(n_8016),
.D(n_5869),
.Y(n_20405)
);

INVx1_ASAP7_75t_L g20406 ( 
.A(n_20251),
.Y(n_20406)
);

AOI22xp33_ASAP7_75t_L g20407 ( 
.A1(n_20270),
.A2(n_8954),
.B1(n_8997),
.B2(n_8672),
.Y(n_20407)
);

NOR2x1_ASAP7_75t_L g20408 ( 
.A(n_20289),
.B(n_7104),
.Y(n_20408)
);

NOR3xp33_ASAP7_75t_SL g20409 ( 
.A(n_20271),
.B(n_7547),
.C(n_7529),
.Y(n_20409)
);

INVx2_ASAP7_75t_SL g20410 ( 
.A(n_20297),
.Y(n_20410)
);

NAND2xp5_ASAP7_75t_L g20411 ( 
.A(n_20284),
.B(n_7257),
.Y(n_20411)
);

INVx1_ASAP7_75t_L g20412 ( 
.A(n_20257),
.Y(n_20412)
);

INVx1_ASAP7_75t_L g20413 ( 
.A(n_20301),
.Y(n_20413)
);

INVx1_ASAP7_75t_L g20414 ( 
.A(n_20369),
.Y(n_20414)
);

NAND4xp75_ASAP7_75t_L g20415 ( 
.A(n_20262),
.B(n_8016),
.C(n_5869),
.D(n_5878),
.Y(n_20415)
);

NOR2x1_ASAP7_75t_L g20416 ( 
.A(n_20250),
.B(n_7104),
.Y(n_20416)
);

NOR3x2_ASAP7_75t_L g20417 ( 
.A(n_20249),
.B(n_7205),
.C(n_7180),
.Y(n_20417)
);

NAND3xp33_ASAP7_75t_SL g20418 ( 
.A(n_20255),
.B(n_8019),
.C(n_7938),
.Y(n_20418)
);

NOR2x1_ASAP7_75t_L g20419 ( 
.A(n_20253),
.B(n_7180),
.Y(n_20419)
);

INVx2_ASAP7_75t_L g20420 ( 
.A(n_20302),
.Y(n_20420)
);

NOR2x1_ASAP7_75t_L g20421 ( 
.A(n_20263),
.B(n_7180),
.Y(n_20421)
);

OA22x2_ASAP7_75t_L g20422 ( 
.A1(n_20256),
.A2(n_7698),
.B1(n_7714),
.B2(n_7565),
.Y(n_20422)
);

NAND4xp75_ASAP7_75t_L g20423 ( 
.A(n_20334),
.B(n_8016),
.C(n_5869),
.D(n_5878),
.Y(n_20423)
);

OR2x2_ASAP7_75t_L g20424 ( 
.A(n_20315),
.B(n_9579),
.Y(n_20424)
);

INVx1_ASAP7_75t_L g20425 ( 
.A(n_20332),
.Y(n_20425)
);

OR2x2_ASAP7_75t_L g20426 ( 
.A(n_20264),
.B(n_9579),
.Y(n_20426)
);

INVx1_ASAP7_75t_L g20427 ( 
.A(n_20258),
.Y(n_20427)
);

NOR2xp33_ASAP7_75t_L g20428 ( 
.A(n_20254),
.B(n_20300),
.Y(n_20428)
);

NOR3xp33_ASAP7_75t_L g20429 ( 
.A(n_20340),
.B(n_20322),
.C(n_20335),
.Y(n_20429)
);

INVx1_ASAP7_75t_L g20430 ( 
.A(n_20305),
.Y(n_20430)
);

INVx2_ASAP7_75t_L g20431 ( 
.A(n_20264),
.Y(n_20431)
);

INVx1_ASAP7_75t_L g20432 ( 
.A(n_20285),
.Y(n_20432)
);

INVx1_ASAP7_75t_L g20433 ( 
.A(n_20260),
.Y(n_20433)
);

NAND3xp33_ASAP7_75t_SL g20434 ( 
.A(n_20294),
.B(n_8019),
.C(n_7938),
.Y(n_20434)
);

NAND4xp75_ASAP7_75t_L g20435 ( 
.A(n_20252),
.B(n_8016),
.C(n_5878),
.D(n_5887),
.Y(n_20435)
);

NAND2xp5_ASAP7_75t_L g20436 ( 
.A(n_20317),
.B(n_7257),
.Y(n_20436)
);

OAI21xp5_ASAP7_75t_L g20437 ( 
.A1(n_20282),
.A2(n_8368),
.B(n_9074),
.Y(n_20437)
);

NAND3xp33_ASAP7_75t_L g20438 ( 
.A(n_20386),
.B(n_8091),
.C(n_7915),
.Y(n_20438)
);

NAND2xp5_ASAP7_75t_L g20439 ( 
.A(n_20311),
.B(n_7257),
.Y(n_20439)
);

NAND3xp33_ASAP7_75t_L g20440 ( 
.A(n_20359),
.B(n_8091),
.C(n_7915),
.Y(n_20440)
);

NOR4xp75_ASAP7_75t_L g20441 ( 
.A(n_20273),
.B(n_7173),
.C(n_7267),
.D(n_7156),
.Y(n_20441)
);

NAND4xp75_ASAP7_75t_L g20442 ( 
.A(n_20353),
.B(n_8016),
.C(n_5887),
.D(n_5935),
.Y(n_20442)
);

NAND2xp33_ASAP7_75t_L g20443 ( 
.A(n_20373),
.B(n_8672),
.Y(n_20443)
);

NOR2xp33_ASAP7_75t_SL g20444 ( 
.A(n_20269),
.B(n_7674),
.Y(n_20444)
);

NOR2x1_ASAP7_75t_L g20445 ( 
.A(n_20348),
.B(n_7180),
.Y(n_20445)
);

INVx1_ASAP7_75t_L g20446 ( 
.A(n_20309),
.Y(n_20446)
);

NOR3xp33_ASAP7_75t_L g20447 ( 
.A(n_20291),
.B(n_6411),
.C(n_7340),
.Y(n_20447)
);

INVx2_ASAP7_75t_L g20448 ( 
.A(n_20347),
.Y(n_20448)
);

NOR3x1_ASAP7_75t_L g20449 ( 
.A(n_20339),
.B(n_9068),
.C(n_9067),
.Y(n_20449)
);

NOR2x1_ASAP7_75t_L g20450 ( 
.A(n_20336),
.B(n_20313),
.Y(n_20450)
);

INVx2_ASAP7_75t_SL g20451 ( 
.A(n_20378),
.Y(n_20451)
);

NAND4xp25_ASAP7_75t_L g20452 ( 
.A(n_20367),
.B(n_7714),
.C(n_7724),
.D(n_7698),
.Y(n_20452)
);

NAND3xp33_ASAP7_75t_L g20453 ( 
.A(n_20306),
.B(n_8091),
.C(n_7915),
.Y(n_20453)
);

INVx1_ASAP7_75t_L g20454 ( 
.A(n_20323),
.Y(n_20454)
);

NAND2xp5_ASAP7_75t_SL g20455 ( 
.A(n_20337),
.B(n_20281),
.Y(n_20455)
);

NAND2xp5_ASAP7_75t_L g20456 ( 
.A(n_20351),
.B(n_20280),
.Y(n_20456)
);

NOR3xp33_ASAP7_75t_SL g20457 ( 
.A(n_20376),
.B(n_7557),
.C(n_7556),
.Y(n_20457)
);

OR2x2_ASAP7_75t_L g20458 ( 
.A(n_20344),
.B(n_7535),
.Y(n_20458)
);

XNOR2x1_ASAP7_75t_L g20459 ( 
.A(n_20329),
.B(n_8336),
.Y(n_20459)
);

AND2x2_ASAP7_75t_L g20460 ( 
.A(n_20362),
.B(n_9387),
.Y(n_20460)
);

INVx1_ASAP7_75t_L g20461 ( 
.A(n_20331),
.Y(n_20461)
);

NOR2xp67_ASAP7_75t_L g20462 ( 
.A(n_20360),
.B(n_20374),
.Y(n_20462)
);

INVxp33_ASAP7_75t_L g20463 ( 
.A(n_20327),
.Y(n_20463)
);

NAND3xp33_ASAP7_75t_SL g20464 ( 
.A(n_20278),
.B(n_8019),
.C(n_7938),
.Y(n_20464)
);

NOR3xp33_ASAP7_75t_L g20465 ( 
.A(n_20388),
.B(n_7392),
.C(n_7340),
.Y(n_20465)
);

AND2x4_ASAP7_75t_L g20466 ( 
.A(n_20321),
.B(n_7486),
.Y(n_20466)
);

CKINVDCx16_ASAP7_75t_R g20467 ( 
.A(n_20389),
.Y(n_20467)
);

NAND3xp33_ASAP7_75t_L g20468 ( 
.A(n_20299),
.B(n_8091),
.C(n_7915),
.Y(n_20468)
);

NOR2xp33_ASAP7_75t_SL g20469 ( 
.A(n_20350),
.B(n_4532),
.Y(n_20469)
);

INVx1_ASAP7_75t_L g20470 ( 
.A(n_20372),
.Y(n_20470)
);

AOI22xp5_ASAP7_75t_L g20471 ( 
.A1(n_20358),
.A2(n_8954),
.B1(n_9191),
.B2(n_8997),
.Y(n_20471)
);

NOR2x1_ASAP7_75t_L g20472 ( 
.A(n_20326),
.B(n_7205),
.Y(n_20472)
);

AOI22xp5_ASAP7_75t_L g20473 ( 
.A1(n_20274),
.A2(n_8954),
.B1(n_9191),
.B2(n_8997),
.Y(n_20473)
);

NAND2xp5_ASAP7_75t_L g20474 ( 
.A(n_20320),
.B(n_7257),
.Y(n_20474)
);

INVx1_ASAP7_75t_L g20475 ( 
.A(n_20298),
.Y(n_20475)
);

NAND4xp75_ASAP7_75t_L g20476 ( 
.A(n_20341),
.B(n_8016),
.C(n_5887),
.D(n_5935),
.Y(n_20476)
);

NAND2xp5_ASAP7_75t_L g20477 ( 
.A(n_20356),
.B(n_7257),
.Y(n_20477)
);

INVx1_ASAP7_75t_L g20478 ( 
.A(n_20314),
.Y(n_20478)
);

INVxp67_ASAP7_75t_L g20479 ( 
.A(n_20368),
.Y(n_20479)
);

INVxp67_ASAP7_75t_SL g20480 ( 
.A(n_20307),
.Y(n_20480)
);

NAND4xp75_ASAP7_75t_L g20481 ( 
.A(n_20392),
.B(n_5935),
.C(n_5957),
.D(n_5805),
.Y(n_20481)
);

NOR2x1_ASAP7_75t_L g20482 ( 
.A(n_20312),
.B(n_20375),
.Y(n_20482)
);

AND2x2_ASAP7_75t_L g20483 ( 
.A(n_20316),
.B(n_9387),
.Y(n_20483)
);

NOR2xp67_ASAP7_75t_L g20484 ( 
.A(n_20267),
.B(n_7340),
.Y(n_20484)
);

AND2x2_ASAP7_75t_L g20485 ( 
.A(n_20357),
.B(n_9559),
.Y(n_20485)
);

INVxp67_ASAP7_75t_SL g20486 ( 
.A(n_20342),
.Y(n_20486)
);

OA22x2_ASAP7_75t_L g20487 ( 
.A1(n_20318),
.A2(n_7714),
.B1(n_7724),
.B2(n_7698),
.Y(n_20487)
);

NOR2x1_ASAP7_75t_L g20488 ( 
.A(n_20346),
.B(n_7205),
.Y(n_20488)
);

NAND4xp75_ASAP7_75t_L g20489 ( 
.A(n_20296),
.B(n_5957),
.C(n_5805),
.D(n_7557),
.Y(n_20489)
);

AOI21xp5_ASAP7_75t_L g20490 ( 
.A1(n_20370),
.A2(n_20349),
.B(n_20354),
.Y(n_20490)
);

OAI22xp5_ASAP7_75t_L g20491 ( 
.A1(n_20382),
.A2(n_7215),
.B1(n_7249),
.B2(n_7222),
.Y(n_20491)
);

NOR3x2_ASAP7_75t_L g20492 ( 
.A(n_20303),
.B(n_7205),
.C(n_7741),
.Y(n_20492)
);

OA21x2_ASAP7_75t_L g20493 ( 
.A1(n_20290),
.A2(n_8768),
.B(n_8754),
.Y(n_20493)
);

NAND3x1_ASAP7_75t_SL g20494 ( 
.A(n_20381),
.B(n_7014),
.C(n_7002),
.Y(n_20494)
);

INVx1_ASAP7_75t_L g20495 ( 
.A(n_20319),
.Y(n_20495)
);

OR2x2_ASAP7_75t_L g20496 ( 
.A(n_20393),
.B(n_20366),
.Y(n_20496)
);

BUFx8_ASAP7_75t_SL g20497 ( 
.A(n_20288),
.Y(n_20497)
);

BUFx12f_ASAP7_75t_L g20498 ( 
.A(n_20394),
.Y(n_20498)
);

NAND3xp33_ASAP7_75t_SL g20499 ( 
.A(n_20364),
.B(n_7938),
.C(n_7842),
.Y(n_20499)
);

AND2x2_ASAP7_75t_L g20500 ( 
.A(n_20365),
.B(n_9559),
.Y(n_20500)
);

INVx1_ASAP7_75t_SL g20501 ( 
.A(n_20308),
.Y(n_20501)
);

NOR3xp33_ASAP7_75t_L g20502 ( 
.A(n_20363),
.B(n_7392),
.C(n_7340),
.Y(n_20502)
);

NAND3xp33_ASAP7_75t_L g20503 ( 
.A(n_20325),
.B(n_8091),
.C(n_7915),
.Y(n_20503)
);

AOI22xp33_ASAP7_75t_SL g20504 ( 
.A1(n_20377),
.A2(n_8997),
.B1(n_9191),
.B2(n_8672),
.Y(n_20504)
);

OAI22xp5_ASAP7_75t_L g20505 ( 
.A1(n_20330),
.A2(n_7215),
.B1(n_7249),
.B2(n_7222),
.Y(n_20505)
);

NAND4xp75_ASAP7_75t_L g20506 ( 
.A(n_20355),
.B(n_5957),
.C(n_5805),
.D(n_7558),
.Y(n_20506)
);

NAND2xp33_ASAP7_75t_L g20507 ( 
.A(n_20352),
.B(n_8672),
.Y(n_20507)
);

NOR2x1_ASAP7_75t_L g20508 ( 
.A(n_20387),
.B(n_6947),
.Y(n_20508)
);

NAND3xp33_ASAP7_75t_L g20509 ( 
.A(n_20338),
.B(n_8091),
.C(n_7040),
.Y(n_20509)
);

NOR2x1_ASAP7_75t_L g20510 ( 
.A(n_20383),
.B(n_6947),
.Y(n_20510)
);

NOR4xp25_ASAP7_75t_L g20511 ( 
.A(n_20324),
.B(n_7901),
.C(n_7724),
.D(n_7842),
.Y(n_20511)
);

AOI22xp5_ASAP7_75t_L g20512 ( 
.A1(n_20333),
.A2(n_8672),
.B1(n_9191),
.B2(n_7561),
.Y(n_20512)
);

NOR2x1_ASAP7_75t_L g20513 ( 
.A(n_20310),
.B(n_6947),
.Y(n_20513)
);

NOR2x1_ASAP7_75t_L g20514 ( 
.A(n_20292),
.B(n_6947),
.Y(n_20514)
);

NAND4xp75_ASAP7_75t_L g20515 ( 
.A(n_20283),
.B(n_7561),
.C(n_7566),
.D(n_7558),
.Y(n_20515)
);

NOR3xp33_ASAP7_75t_L g20516 ( 
.A(n_20295),
.B(n_20361),
.C(n_20293),
.Y(n_20516)
);

XNOR2xp5_ASAP7_75t_L g20517 ( 
.A(n_20410),
.B(n_20304),
.Y(n_20517)
);

NOR3xp33_ASAP7_75t_L g20518 ( 
.A(n_20414),
.B(n_20343),
.C(n_20385),
.Y(n_20518)
);

AOI211xp5_ASAP7_75t_L g20519 ( 
.A1(n_20425),
.A2(n_20395),
.B(n_20268),
.C(n_20391),
.Y(n_20519)
);

NOR3x1_ASAP7_75t_L g20520 ( 
.A(n_20480),
.B(n_20266),
.C(n_20328),
.Y(n_20520)
);

NOR3xp33_ASAP7_75t_L g20521 ( 
.A(n_20406),
.B(n_20276),
.C(n_20379),
.Y(n_20521)
);

OA22x2_ASAP7_75t_L g20522 ( 
.A1(n_20427),
.A2(n_20272),
.B1(n_20371),
.B2(n_20286),
.Y(n_20522)
);

INVx2_ASAP7_75t_SL g20523 ( 
.A(n_20431),
.Y(n_20523)
);

OAI211xp5_ASAP7_75t_SL g20524 ( 
.A1(n_20413),
.A2(n_20345),
.B(n_20287),
.C(n_20390),
.Y(n_20524)
);

OR3x1_ASAP7_75t_L g20525 ( 
.A(n_20428),
.B(n_20275),
.C(n_7561),
.Y(n_20525)
);

NOR3xp33_ASAP7_75t_L g20526 ( 
.A(n_20412),
.B(n_20433),
.C(n_20446),
.Y(n_20526)
);

NAND3xp33_ASAP7_75t_SL g20527 ( 
.A(n_20429),
.B(n_7392),
.C(n_7340),
.Y(n_20527)
);

NAND5xp2_ASAP7_75t_L g20528 ( 
.A(n_20516),
.B(n_7161),
.C(n_7587),
.D(n_7555),
.E(n_7554),
.Y(n_20528)
);

NAND5xp2_ASAP7_75t_L g20529 ( 
.A(n_20479),
.B(n_7161),
.C(n_7587),
.D(n_7555),
.E(n_7554),
.Y(n_20529)
);

NAND5xp2_ASAP7_75t_L g20530 ( 
.A(n_20470),
.B(n_7161),
.C(n_7587),
.D(n_7555),
.E(n_7554),
.Y(n_20530)
);

AND2x4_ASAP7_75t_L g20531 ( 
.A(n_20398),
.B(n_7486),
.Y(n_20531)
);

NAND3xp33_ASAP7_75t_SL g20532 ( 
.A(n_20420),
.B(n_7392),
.C(n_7340),
.Y(n_20532)
);

NOR4xp25_ASAP7_75t_L g20533 ( 
.A(n_20454),
.B(n_8006),
.C(n_8051),
.D(n_8003),
.Y(n_20533)
);

NOR2xp33_ASAP7_75t_SL g20534 ( 
.A(n_20486),
.B(n_4532),
.Y(n_20534)
);

NOR4xp25_ASAP7_75t_L g20535 ( 
.A(n_20461),
.B(n_8006),
.C(n_8051),
.D(n_8003),
.Y(n_20535)
);

INVx1_ASAP7_75t_L g20536 ( 
.A(n_20400),
.Y(n_20536)
);

OAI21xp5_ASAP7_75t_L g20537 ( 
.A1(n_20408),
.A2(n_8368),
.B(n_8585),
.Y(n_20537)
);

NOR4xp25_ASAP7_75t_L g20538 ( 
.A(n_20448),
.B(n_8051),
.C(n_8006),
.D(n_7222),
.Y(n_20538)
);

AND4x2_ASAP7_75t_L g20539 ( 
.A(n_20450),
.B(n_7301),
.C(n_7424),
.D(n_7216),
.Y(n_20539)
);

NOR2xp33_ASAP7_75t_L g20540 ( 
.A(n_20463),
.B(n_6976),
.Y(n_20540)
);

AOI21xp5_ASAP7_75t_L g20541 ( 
.A1(n_20456),
.A2(n_9074),
.B(n_6837),
.Y(n_20541)
);

NOR4xp25_ASAP7_75t_L g20542 ( 
.A(n_20430),
.B(n_20451),
.C(n_20495),
.D(n_20475),
.Y(n_20542)
);

AND4x1_ASAP7_75t_L g20543 ( 
.A(n_20478),
.B(n_7161),
.C(n_7014),
.D(n_7048),
.Y(n_20543)
);

NOR2x1_ASAP7_75t_L g20544 ( 
.A(n_20432),
.B(n_20455),
.Y(n_20544)
);

OAI211xp5_ASAP7_75t_SL g20545 ( 
.A1(n_20496),
.A2(n_8051),
.B(n_8006),
.C(n_7249),
.Y(n_20545)
);

OR3x1_ASAP7_75t_L g20546 ( 
.A(n_20499),
.B(n_7566),
.C(n_7558),
.Y(n_20546)
);

NAND3xp33_ASAP7_75t_SL g20547 ( 
.A(n_20501),
.B(n_7468),
.C(n_7392),
.Y(n_20547)
);

NAND3x1_ASAP7_75t_L g20548 ( 
.A(n_20445),
.B(n_5680),
.C(n_5673),
.Y(n_20548)
);

AOI21xp5_ASAP7_75t_L g20549 ( 
.A1(n_20462),
.A2(n_9074),
.B(n_6837),
.Y(n_20549)
);

NOR4xp25_ASAP7_75t_L g20550 ( 
.A(n_20411),
.B(n_7401),
.C(n_7446),
.D(n_7215),
.Y(n_20550)
);

NAND5xp2_ASAP7_75t_L g20551 ( 
.A(n_20397),
.B(n_7161),
.C(n_7626),
.D(n_7607),
.E(n_7591),
.Y(n_20551)
);

NAND4xp25_ASAP7_75t_L g20552 ( 
.A(n_20419),
.B(n_20421),
.C(n_20482),
.D(n_20416),
.Y(n_20552)
);

NAND4xp25_ASAP7_75t_L g20553 ( 
.A(n_20401),
.B(n_20444),
.C(n_20490),
.D(n_20440),
.Y(n_20553)
);

OA211x2_ASAP7_75t_L g20554 ( 
.A1(n_20469),
.A2(n_9573),
.B(n_9572),
.C(n_8772),
.Y(n_20554)
);

OAI211xp5_ASAP7_75t_L g20555 ( 
.A1(n_20409),
.A2(n_7607),
.B(n_7626),
.C(n_7591),
.Y(n_20555)
);

AOI211xp5_ASAP7_75t_L g20556 ( 
.A1(n_20452),
.A2(n_7889),
.B(n_7918),
.C(n_7834),
.Y(n_20556)
);

OAI211xp5_ASAP7_75t_L g20557 ( 
.A1(n_20511),
.A2(n_7607),
.B(n_7626),
.C(n_7591),
.Y(n_20557)
);

OAI211xp5_ASAP7_75t_SL g20558 ( 
.A1(n_20439),
.A2(n_7446),
.B(n_7450),
.C(n_7401),
.Y(n_20558)
);

NAND2xp5_ASAP7_75t_L g20559 ( 
.A(n_20467),
.B(n_7257),
.Y(n_20559)
);

AOI221xp5_ASAP7_75t_L g20560 ( 
.A1(n_20509),
.A2(n_7098),
.B1(n_7071),
.B2(n_7040),
.C(n_7889),
.Y(n_20560)
);

NAND2x1p5_ASAP7_75t_L g20561 ( 
.A(n_20514),
.B(n_5545),
.Y(n_20561)
);

AOI322xp5_ASAP7_75t_L g20562 ( 
.A1(n_20502),
.A2(n_7632),
.A3(n_7645),
.B1(n_7577),
.B2(n_7771),
.C1(n_7817),
.C2(n_7765),
.Y(n_20562)
);

NAND2xp5_ASAP7_75t_L g20563 ( 
.A(n_20436),
.B(n_7257),
.Y(n_20563)
);

NAND3xp33_ASAP7_75t_L g20564 ( 
.A(n_20507),
.B(n_7161),
.C(n_8091),
.Y(n_20564)
);

AOI211xp5_ASAP7_75t_L g20565 ( 
.A1(n_20484),
.A2(n_7918),
.B(n_7957),
.C(n_7889),
.Y(n_20565)
);

OAI221xp5_ASAP7_75t_SL g20566 ( 
.A1(n_20424),
.A2(n_7661),
.B1(n_7690),
.B2(n_7686),
.C(n_7642),
.Y(n_20566)
);

OAI221xp5_ASAP7_75t_SL g20567 ( 
.A1(n_20458),
.A2(n_7661),
.B1(n_7690),
.B2(n_7686),
.C(n_7642),
.Y(n_20567)
);

NAND4xp25_ASAP7_75t_SL g20568 ( 
.A(n_20472),
.B(n_7446),
.C(n_7450),
.D(n_7401),
.Y(n_20568)
);

OR2x2_ASAP7_75t_L g20569 ( 
.A(n_20404),
.B(n_7642),
.Y(n_20569)
);

OAI221xp5_ASAP7_75t_L g20570 ( 
.A1(n_20402),
.A2(n_7817),
.B1(n_7823),
.B2(n_7771),
.C(n_7765),
.Y(n_20570)
);

NAND3xp33_ASAP7_75t_L g20571 ( 
.A(n_20488),
.B(n_7161),
.C(n_7071),
.Y(n_20571)
);

AND4x1_ASAP7_75t_L g20572 ( 
.A(n_20438),
.B(n_20510),
.C(n_20513),
.D(n_20512),
.Y(n_20572)
);

A2O1A1Ixp33_ASAP7_75t_L g20573 ( 
.A1(n_20457),
.A2(n_8772),
.B(n_8776),
.C(n_8774),
.Y(n_20573)
);

NOR2x1p5_ASAP7_75t_L g20574 ( 
.A(n_20498),
.B(n_7040),
.Y(n_20574)
);

NOR3xp33_ASAP7_75t_L g20575 ( 
.A(n_20464),
.B(n_7468),
.C(n_7392),
.Y(n_20575)
);

AOI22xp5_ASAP7_75t_L g20576 ( 
.A1(n_20418),
.A2(n_9191),
.B1(n_8672),
.B2(n_7040),
.Y(n_20576)
);

AOI211xp5_ASAP7_75t_L g20577 ( 
.A1(n_20443),
.A2(n_7918),
.B(n_7957),
.C(n_7889),
.Y(n_20577)
);

A2O1A1Ixp33_ASAP7_75t_L g20578 ( 
.A1(n_20483),
.A2(n_8772),
.B(n_8776),
.C(n_8774),
.Y(n_20578)
);

O2A1O1Ixp33_ASAP7_75t_L g20579 ( 
.A1(n_20474),
.A2(n_20477),
.B(n_20403),
.C(n_20434),
.Y(n_20579)
);

NAND4xp75_ASAP7_75t_L g20580 ( 
.A(n_20508),
.B(n_7014),
.C(n_7048),
.D(n_7002),
.Y(n_20580)
);

NAND3xp33_ASAP7_75t_L g20581 ( 
.A(n_20459),
.B(n_7071),
.C(n_7040),
.Y(n_20581)
);

NOR2x1_ASAP7_75t_L g20582 ( 
.A(n_20476),
.B(n_6983),
.Y(n_20582)
);

OR3x1_ASAP7_75t_L g20583 ( 
.A(n_20497),
.B(n_7575),
.C(n_7566),
.Y(n_20583)
);

OAI221xp5_ASAP7_75t_L g20584 ( 
.A1(n_20399),
.A2(n_7829),
.B1(n_7836),
.B2(n_7823),
.C(n_7817),
.Y(n_20584)
);

NOR3xp33_ASAP7_75t_L g20585 ( 
.A(n_20494),
.B(n_7478),
.C(n_7468),
.Y(n_20585)
);

AND2x2_ASAP7_75t_L g20586 ( 
.A(n_20466),
.B(n_9275),
.Y(n_20586)
);

AOI221xp5_ASAP7_75t_SL g20587 ( 
.A1(n_20460),
.A2(n_7686),
.B1(n_7700),
.B2(n_7690),
.C(n_7661),
.Y(n_20587)
);

NOR4xp25_ASAP7_75t_L g20588 ( 
.A(n_20485),
.B(n_7446),
.C(n_7450),
.D(n_7401),
.Y(n_20588)
);

AOI221xp5_ASAP7_75t_L g20589 ( 
.A1(n_20500),
.A2(n_7098),
.B1(n_7071),
.B2(n_7040),
.C(n_7889),
.Y(n_20589)
);

NAND5xp2_ASAP7_75t_L g20590 ( 
.A(n_20447),
.B(n_7737),
.C(n_7740),
.D(n_7731),
.E(n_7700),
.Y(n_20590)
);

OR3x1_ASAP7_75t_L g20591 ( 
.A(n_20417),
.B(n_7582),
.C(n_7575),
.Y(n_20591)
);

NOR3xp33_ASAP7_75t_L g20592 ( 
.A(n_20506),
.B(n_7478),
.C(n_7468),
.Y(n_20592)
);

NAND5xp2_ASAP7_75t_L g20593 ( 
.A(n_20465),
.B(n_7737),
.C(n_7740),
.D(n_7731),
.E(n_7700),
.Y(n_20593)
);

NAND2xp5_ASAP7_75t_SL g20594 ( 
.A(n_20422),
.B(n_7040),
.Y(n_20594)
);

AND2x2_ASAP7_75t_L g20595 ( 
.A(n_20466),
.B(n_9275),
.Y(n_20595)
);

AOI221xp5_ASAP7_75t_L g20596 ( 
.A1(n_20453),
.A2(n_7098),
.B1(n_7918),
.B2(n_7957),
.C(n_7889),
.Y(n_20596)
);

AOI221xp5_ASAP7_75t_L g20597 ( 
.A1(n_20505),
.A2(n_7098),
.B1(n_7918),
.B2(n_7957),
.C(n_7889),
.Y(n_20597)
);

OAI211xp5_ASAP7_75t_L g20598 ( 
.A1(n_20468),
.A2(n_7731),
.B(n_7740),
.C(n_7737),
.Y(n_20598)
);

NAND4xp75_ASAP7_75t_L g20599 ( 
.A(n_20449),
.B(n_7048),
.C(n_7058),
.D(n_7002),
.Y(n_20599)
);

OAI221xp5_ASAP7_75t_L g20600 ( 
.A1(n_20487),
.A2(n_7829),
.B1(n_7855),
.B2(n_7836),
.C(n_7823),
.Y(n_20600)
);

AND2x2_ASAP7_75t_L g20601 ( 
.A(n_20473),
.B(n_9275),
.Y(n_20601)
);

NAND5xp2_ASAP7_75t_L g20602 ( 
.A(n_20471),
.B(n_7750),
.C(n_7836),
.D(n_7855),
.E(n_7829),
.Y(n_20602)
);

INVxp67_ASAP7_75t_SL g20603 ( 
.A(n_20426),
.Y(n_20603)
);

AND5x1_ASAP7_75t_L g20604 ( 
.A(n_20441),
.B(n_7257),
.C(n_7750),
.D(n_8478),
.E(n_8472),
.Y(n_20604)
);

HB1xp67_ASAP7_75t_L g20605 ( 
.A(n_20481),
.Y(n_20605)
);

OR5x1_ASAP7_75t_L g20606 ( 
.A(n_20515),
.B(n_8748),
.C(n_8768),
.D(n_9573),
.E(n_9572),
.Y(n_20606)
);

AOI22xp5_ASAP7_75t_L g20607 ( 
.A1(n_20503),
.A2(n_9191),
.B1(n_8672),
.B2(n_7098),
.Y(n_20607)
);

INVxp33_ASAP7_75t_L g20608 ( 
.A(n_20435),
.Y(n_20608)
);

NOR3xp33_ASAP7_75t_SL g20609 ( 
.A(n_20489),
.B(n_7582),
.C(n_7575),
.Y(n_20609)
);

NOR3xp33_ASAP7_75t_L g20610 ( 
.A(n_20405),
.B(n_7478),
.C(n_7468),
.Y(n_20610)
);

NAND4xp25_ASAP7_75t_L g20611 ( 
.A(n_20504),
.B(n_7750),
.C(n_7862),
.D(n_7855),
.Y(n_20611)
);

NOR2x1_ASAP7_75t_L g20612 ( 
.A(n_20415),
.B(n_6983),
.Y(n_20612)
);

INVx1_ASAP7_75t_L g20613 ( 
.A(n_20492),
.Y(n_20613)
);

OAI211xp5_ASAP7_75t_SL g20614 ( 
.A1(n_20491),
.A2(n_7450),
.B(n_7583),
.C(n_7582),
.Y(n_20614)
);

NOR3xp33_ASAP7_75t_L g20615 ( 
.A(n_20442),
.B(n_7478),
.C(n_7468),
.Y(n_20615)
);

AOI322xp5_ASAP7_75t_L g20616 ( 
.A1(n_20407),
.A2(n_7632),
.A3(n_7645),
.B1(n_7577),
.B2(n_7904),
.C1(n_7886),
.C2(n_7862),
.Y(n_20616)
);

OAI211xp5_ASAP7_75t_SL g20617 ( 
.A1(n_20437),
.A2(n_7584),
.B(n_7585),
.C(n_7583),
.Y(n_20617)
);

OAI221xp5_ASAP7_75t_SL g20618 ( 
.A1(n_20423),
.A2(n_7886),
.B1(n_7904),
.B2(n_7862),
.C(n_7008),
.Y(n_20618)
);

OAI221xp5_ASAP7_75t_L g20619 ( 
.A1(n_20493),
.A2(n_7904),
.B1(n_7886),
.B2(n_7831),
.C(n_7798),
.Y(n_20619)
);

NAND3xp33_ASAP7_75t_L g20620 ( 
.A(n_20493),
.B(n_7098),
.C(n_6267),
.Y(n_20620)
);

AOI211x1_ASAP7_75t_L g20621 ( 
.A1(n_20427),
.A2(n_7584),
.B(n_7585),
.C(n_7583),
.Y(n_20621)
);

INVx2_ASAP7_75t_L g20622 ( 
.A(n_20410),
.Y(n_20622)
);

NAND4xp75_ASAP7_75t_L g20623 ( 
.A(n_20410),
.B(n_7176),
.C(n_7188),
.D(n_7058),
.Y(n_20623)
);

NOR5xp2_ASAP7_75t_L g20624 ( 
.A(n_20427),
.B(n_7588),
.C(n_7589),
.D(n_7585),
.E(n_7584),
.Y(n_20624)
);

OAI221xp5_ASAP7_75t_L g20625 ( 
.A1(n_20410),
.A2(n_7798),
.B1(n_7831),
.B2(n_7005),
.C(n_7889),
.Y(n_20625)
);

NAND2xp5_ASAP7_75t_L g20626 ( 
.A(n_20410),
.B(n_7380),
.Y(n_20626)
);

NOR2x1_ASAP7_75t_L g20627 ( 
.A(n_20622),
.B(n_6983),
.Y(n_20627)
);

NAND2xp5_ASAP7_75t_SL g20628 ( 
.A(n_20526),
.B(n_7976),
.Y(n_20628)
);

INVx1_ASAP7_75t_L g20629 ( 
.A(n_20536),
.Y(n_20629)
);

INVx2_ASAP7_75t_SL g20630 ( 
.A(n_20544),
.Y(n_20630)
);

INVx1_ASAP7_75t_L g20631 ( 
.A(n_20552),
.Y(n_20631)
);

NAND4xp75_ASAP7_75t_L g20632 ( 
.A(n_20523),
.B(n_6338),
.C(n_6492),
.D(n_6477),
.Y(n_20632)
);

INVx1_ASAP7_75t_L g20633 ( 
.A(n_20613),
.Y(n_20633)
);

INVx1_ASAP7_75t_L g20634 ( 
.A(n_20520),
.Y(n_20634)
);

NOR3xp33_ASAP7_75t_L g20635 ( 
.A(n_20603),
.B(n_7525),
.C(n_7478),
.Y(n_20635)
);

INVx1_ASAP7_75t_L g20636 ( 
.A(n_20521),
.Y(n_20636)
);

INVx1_ASAP7_75t_L g20637 ( 
.A(n_20517),
.Y(n_20637)
);

OR2x2_ASAP7_75t_L g20638 ( 
.A(n_20542),
.B(n_20626),
.Y(n_20638)
);

NOR3xp33_ASAP7_75t_L g20639 ( 
.A(n_20553),
.B(n_7525),
.C(n_7478),
.Y(n_20639)
);

NAND4xp75_ASAP7_75t_L g20640 ( 
.A(n_20540),
.B(n_6477),
.C(n_6562),
.D(n_6492),
.Y(n_20640)
);

NOR2x1_ASAP7_75t_L g20641 ( 
.A(n_20524),
.B(n_6983),
.Y(n_20641)
);

AO22x2_ASAP7_75t_L g20642 ( 
.A1(n_20518),
.A2(n_7798),
.B1(n_7831),
.B2(n_7005),
.Y(n_20642)
);

INVx1_ASAP7_75t_L g20643 ( 
.A(n_20579),
.Y(n_20643)
);

XOR2x2_ASAP7_75t_L g20644 ( 
.A(n_20519),
.B(n_5705),
.Y(n_20644)
);

BUFx6f_ASAP7_75t_L g20645 ( 
.A(n_20569),
.Y(n_20645)
);

NOR2x1_ASAP7_75t_L g20646 ( 
.A(n_20525),
.B(n_6983),
.Y(n_20646)
);

INVx2_ASAP7_75t_L g20647 ( 
.A(n_20561),
.Y(n_20647)
);

NOR2x1p5_ASAP7_75t_L g20648 ( 
.A(n_20559),
.B(n_5705),
.Y(n_20648)
);

OR2x2_ASAP7_75t_L g20649 ( 
.A(n_20550),
.B(n_8666),
.Y(n_20649)
);

NAND4xp75_ASAP7_75t_L g20650 ( 
.A(n_20563),
.B(n_6477),
.C(n_6562),
.D(n_6492),
.Y(n_20650)
);

AO22x1_ASAP7_75t_L g20651 ( 
.A1(n_20608),
.A2(n_9191),
.B1(n_6267),
.B2(n_6812),
.Y(n_20651)
);

NAND4xp75_ASAP7_75t_L g20652 ( 
.A(n_20582),
.B(n_6562),
.C(n_6633),
.D(n_6610),
.Y(n_20652)
);

AND2x2_ASAP7_75t_L g20653 ( 
.A(n_20531),
.B(n_8666),
.Y(n_20653)
);

INVx2_ASAP7_75t_SL g20654 ( 
.A(n_20572),
.Y(n_20654)
);

NOR2x1_ASAP7_75t_L g20655 ( 
.A(n_20599),
.B(n_6994),
.Y(n_20655)
);

INVxp33_ASAP7_75t_SL g20656 ( 
.A(n_20522),
.Y(n_20656)
);

NAND4xp75_ASAP7_75t_L g20657 ( 
.A(n_20594),
.B(n_6610),
.C(n_6637),
.D(n_6633),
.Y(n_20657)
);

AND2x2_ASAP7_75t_SL g20658 ( 
.A(n_20605),
.B(n_6837),
.Y(n_20658)
);

NOR2xp33_ASAP7_75t_L g20659 ( 
.A(n_20534),
.B(n_7380),
.Y(n_20659)
);

AOI22xp5_ASAP7_75t_L g20660 ( 
.A1(n_20574),
.A2(n_9191),
.B1(n_7301),
.B2(n_7424),
.Y(n_20660)
);

AND2x4_ASAP7_75t_L g20661 ( 
.A(n_20586),
.B(n_7486),
.Y(n_20661)
);

AO22x1_ASAP7_75t_L g20662 ( 
.A1(n_20531),
.A2(n_20612),
.B1(n_20575),
.B2(n_20595),
.Y(n_20662)
);

INVx2_ASAP7_75t_L g20663 ( 
.A(n_20583),
.Y(n_20663)
);

INVx1_ASAP7_75t_L g20664 ( 
.A(n_20546),
.Y(n_20664)
);

OR3x2_ASAP7_75t_L g20665 ( 
.A(n_20528),
.B(n_8125),
.C(n_8082),
.Y(n_20665)
);

INVx1_ASAP7_75t_SL g20666 ( 
.A(n_20591),
.Y(n_20666)
);

INVx1_ASAP7_75t_L g20667 ( 
.A(n_20548),
.Y(n_20667)
);

INVx1_ASAP7_75t_L g20668 ( 
.A(n_20557),
.Y(n_20668)
);

NAND4xp75_ASAP7_75t_L g20669 ( 
.A(n_20587),
.B(n_6610),
.C(n_6637),
.D(n_6633),
.Y(n_20669)
);

INVx1_ASAP7_75t_L g20670 ( 
.A(n_20581),
.Y(n_20670)
);

OAI22xp33_ASAP7_75t_L g20671 ( 
.A1(n_20571),
.A2(n_7918),
.B1(n_7957),
.B2(n_7889),
.Y(n_20671)
);

AND2x4_ASAP7_75t_L g20672 ( 
.A(n_20564),
.B(n_7486),
.Y(n_20672)
);

AND2x4_ASAP7_75t_L g20673 ( 
.A(n_20601),
.B(n_7486),
.Y(n_20673)
);

INVx1_ASAP7_75t_L g20674 ( 
.A(n_20558),
.Y(n_20674)
);

NOR2x1_ASAP7_75t_L g20675 ( 
.A(n_20611),
.B(n_6994),
.Y(n_20675)
);

OR2x2_ASAP7_75t_L g20676 ( 
.A(n_20566),
.B(n_8666),
.Y(n_20676)
);

INVx2_ASAP7_75t_L g20677 ( 
.A(n_20620),
.Y(n_20677)
);

INVxp33_ASAP7_75t_SL g20678 ( 
.A(n_20533),
.Y(n_20678)
);

HB1xp67_ASAP7_75t_L g20679 ( 
.A(n_20570),
.Y(n_20679)
);

INVx1_ASAP7_75t_L g20680 ( 
.A(n_20545),
.Y(n_20680)
);

OA22x2_ASAP7_75t_L g20681 ( 
.A1(n_20555),
.A2(n_8478),
.B1(n_8491),
.B2(n_8472),
.Y(n_20681)
);

AND2x2_ASAP7_75t_L g20682 ( 
.A(n_20535),
.B(n_8666),
.Y(n_20682)
);

NOR4xp25_ASAP7_75t_L g20683 ( 
.A(n_20598),
.B(n_7589),
.C(n_7590),
.D(n_7588),
.Y(n_20683)
);

INVx1_ASAP7_75t_L g20684 ( 
.A(n_20609),
.Y(n_20684)
);

NAND4xp75_ASAP7_75t_L g20685 ( 
.A(n_20589),
.B(n_6637),
.C(n_6657),
.D(n_6656),
.Y(n_20685)
);

OAI221xp5_ASAP7_75t_L g20686 ( 
.A1(n_20604),
.A2(n_7005),
.B1(n_7918),
.B2(n_7957),
.C(n_6837),
.Y(n_20686)
);

NOR2xp33_ASAP7_75t_L g20687 ( 
.A(n_20602),
.B(n_7380),
.Y(n_20687)
);

HB1xp67_ASAP7_75t_L g20688 ( 
.A(n_20580),
.Y(n_20688)
);

AOI221xp5_ASAP7_75t_L g20689 ( 
.A1(n_20588),
.A2(n_7957),
.B1(n_7918),
.B2(n_7995),
.C(n_7976),
.Y(n_20689)
);

NAND4xp25_ASAP7_75t_L g20690 ( 
.A(n_20593),
.B(n_5717),
.C(n_5705),
.D(n_6942),
.Y(n_20690)
);

INVx1_ASAP7_75t_L g20691 ( 
.A(n_20539),
.Y(n_20691)
);

NAND4xp75_ASAP7_75t_L g20692 ( 
.A(n_20560),
.B(n_6656),
.C(n_6678),
.D(n_6657),
.Y(n_20692)
);

NAND4xp75_ASAP7_75t_L g20693 ( 
.A(n_20621),
.B(n_6656),
.C(n_6678),
.D(n_6657),
.Y(n_20693)
);

NOR2x1_ASAP7_75t_L g20694 ( 
.A(n_20527),
.B(n_6994),
.Y(n_20694)
);

AND2x4_ASAP7_75t_L g20695 ( 
.A(n_20592),
.B(n_5705),
.Y(n_20695)
);

INVx1_ASAP7_75t_L g20696 ( 
.A(n_20617),
.Y(n_20696)
);

INVxp33_ASAP7_75t_L g20697 ( 
.A(n_20538),
.Y(n_20697)
);

NAND3x1_ASAP7_75t_SL g20698 ( 
.A(n_20596),
.B(n_7301),
.C(n_7216),
.Y(n_20698)
);

NOR2xp33_ASAP7_75t_L g20699 ( 
.A(n_20590),
.B(n_7380),
.Y(n_20699)
);

XOR2xp5_ASAP7_75t_L g20700 ( 
.A(n_20547),
.B(n_4532),
.Y(n_20700)
);

NOR3xp33_ASAP7_75t_SL g20701 ( 
.A(n_20618),
.B(n_20600),
.C(n_20532),
.Y(n_20701)
);

NAND2xp5_ASAP7_75t_L g20702 ( 
.A(n_20556),
.B(n_7380),
.Y(n_20702)
);

NAND3xp33_ASAP7_75t_L g20703 ( 
.A(n_20567),
.B(n_6267),
.C(n_6225),
.Y(n_20703)
);

INVx1_ASAP7_75t_L g20704 ( 
.A(n_20619),
.Y(n_20704)
);

INVx1_ASAP7_75t_L g20705 ( 
.A(n_20543),
.Y(n_20705)
);

BUFx2_ASAP7_75t_L g20706 ( 
.A(n_20576),
.Y(n_20706)
);

INVx1_ASAP7_75t_L g20707 ( 
.A(n_20584),
.Y(n_20707)
);

INVx1_ASAP7_75t_L g20708 ( 
.A(n_20529),
.Y(n_20708)
);

NOR2xp33_ASAP7_75t_L g20709 ( 
.A(n_20551),
.B(n_7380),
.Y(n_20709)
);

NOR2x1_ASAP7_75t_L g20710 ( 
.A(n_20568),
.B(n_20530),
.Y(n_20710)
);

NOR2x1_ASAP7_75t_L g20711 ( 
.A(n_20614),
.B(n_6994),
.Y(n_20711)
);

INVx1_ASAP7_75t_L g20712 ( 
.A(n_20585),
.Y(n_20712)
);

INVx1_ASAP7_75t_L g20713 ( 
.A(n_20577),
.Y(n_20713)
);

AOI22xp5_ASAP7_75t_L g20714 ( 
.A1(n_20610),
.A2(n_9191),
.B1(n_7301),
.B2(n_7424),
.Y(n_20714)
);

OR3x2_ASAP7_75t_L g20715 ( 
.A(n_20615),
.B(n_20565),
.C(n_20624),
.Y(n_20715)
);

INVx1_ASAP7_75t_L g20716 ( 
.A(n_20607),
.Y(n_20716)
);

AOI221xp5_ASAP7_75t_SL g20717 ( 
.A1(n_20549),
.A2(n_7957),
.B1(n_7918),
.B2(n_7590),
.C(n_7593),
.Y(n_20717)
);

INVx2_ASAP7_75t_L g20718 ( 
.A(n_20606),
.Y(n_20718)
);

INVx2_ASAP7_75t_L g20719 ( 
.A(n_20623),
.Y(n_20719)
);

AO22x2_ASAP7_75t_L g20720 ( 
.A1(n_20537),
.A2(n_8070),
.B1(n_8094),
.B2(n_8125),
.Y(n_20720)
);

XNOR2xp5_ASAP7_75t_L g20721 ( 
.A(n_20597),
.B(n_8336),
.Y(n_20721)
);

XOR2xp5_ASAP7_75t_L g20722 ( 
.A(n_20554),
.B(n_4532),
.Y(n_20722)
);

INVx1_ASAP7_75t_L g20723 ( 
.A(n_20541),
.Y(n_20723)
);

INVx2_ASAP7_75t_L g20724 ( 
.A(n_20625),
.Y(n_20724)
);

CKINVDCx16_ASAP7_75t_R g20725 ( 
.A(n_20630),
.Y(n_20725)
);

NAND2x1_ASAP7_75t_L g20726 ( 
.A(n_20634),
.B(n_20616),
.Y(n_20726)
);

NAND4xp25_ASAP7_75t_L g20727 ( 
.A(n_20656),
.B(n_20562),
.C(n_20573),
.D(n_20578),
.Y(n_20727)
);

NOR4xp25_ASAP7_75t_L g20728 ( 
.A(n_20643),
.B(n_7589),
.C(n_7590),
.D(n_7588),
.Y(n_20728)
);

NAND4xp25_ASAP7_75t_L g20729 ( 
.A(n_20629),
.B(n_5717),
.C(n_7061),
.D(n_6942),
.Y(n_20729)
);

NAND2xp5_ASAP7_75t_L g20730 ( 
.A(n_20637),
.B(n_8666),
.Y(n_20730)
);

NOR4xp25_ASAP7_75t_L g20731 ( 
.A(n_20654),
.B(n_7594),
.C(n_7596),
.D(n_7593),
.Y(n_20731)
);

NAND2xp5_ASAP7_75t_L g20732 ( 
.A(n_20631),
.B(n_20645),
.Y(n_20732)
);

NOR3xp33_ASAP7_75t_SL g20733 ( 
.A(n_20636),
.B(n_7594),
.C(n_7593),
.Y(n_20733)
);

OAI211xp5_ASAP7_75t_SL g20734 ( 
.A1(n_20638),
.A2(n_5673),
.B(n_5685),
.C(n_5680),
.Y(n_20734)
);

AND2x4_ASAP7_75t_L g20735 ( 
.A(n_20663),
.B(n_7553),
.Y(n_20735)
);

NAND4xp75_ASAP7_75t_L g20736 ( 
.A(n_20633),
.B(n_6709),
.C(n_6711),
.D(n_6678),
.Y(n_20736)
);

NOR5xp2_ASAP7_75t_L g20737 ( 
.A(n_20679),
.B(n_7601),
.C(n_7610),
.D(n_7596),
.E(n_7594),
.Y(n_20737)
);

XNOR2xp5_ASAP7_75t_L g20738 ( 
.A(n_20708),
.B(n_8666),
.Y(n_20738)
);

NOR3xp33_ASAP7_75t_L g20739 ( 
.A(n_20704),
.B(n_7542),
.C(n_7525),
.Y(n_20739)
);

NOR5xp2_ASAP7_75t_L g20740 ( 
.A(n_20688),
.B(n_7610),
.C(n_7612),
.D(n_7601),
.E(n_7596),
.Y(n_20740)
);

AO211x2_ASAP7_75t_L g20741 ( 
.A1(n_20664),
.A2(n_7610),
.B(n_7612),
.C(n_7601),
.Y(n_20741)
);

NOR3xp33_ASAP7_75t_L g20742 ( 
.A(n_20666),
.B(n_7542),
.C(n_7525),
.Y(n_20742)
);

NAND4xp75_ASAP7_75t_L g20743 ( 
.A(n_20712),
.B(n_6711),
.C(n_6774),
.D(n_6709),
.Y(n_20743)
);

OAI222xp33_ASAP7_75t_L g20744 ( 
.A1(n_20718),
.A2(n_8700),
.B1(n_8876),
.B2(n_8962),
.C1(n_8803),
.C2(n_9275),
.Y(n_20744)
);

NOR2xp67_ASAP7_75t_SL g20745 ( 
.A(n_20645),
.B(n_5545),
.Y(n_20745)
);

NAND5xp2_ASAP7_75t_L g20746 ( 
.A(n_20678),
.B(n_4622),
.C(n_7216),
.D(n_7424),
.E(n_7301),
.Y(n_20746)
);

AND2x4_ASAP7_75t_L g20747 ( 
.A(n_20647),
.B(n_7553),
.Y(n_20747)
);

NAND3xp33_ASAP7_75t_L g20748 ( 
.A(n_20707),
.B(n_6267),
.C(n_6225),
.Y(n_20748)
);

NAND3xp33_ASAP7_75t_L g20749 ( 
.A(n_20668),
.B(n_6267),
.C(n_6225),
.Y(n_20749)
);

NOR4xp75_ASAP7_75t_L g20750 ( 
.A(n_20628),
.B(n_7173),
.C(n_7267),
.D(n_7156),
.Y(n_20750)
);

NOR2x1p5_ASAP7_75t_L g20751 ( 
.A(n_20691),
.B(n_5717),
.Y(n_20751)
);

AOI21xp5_ASAP7_75t_L g20752 ( 
.A1(n_20662),
.A2(n_9421),
.B(n_8592),
.Y(n_20752)
);

INVx3_ASAP7_75t_L g20753 ( 
.A(n_20644),
.Y(n_20753)
);

NOR3xp33_ASAP7_75t_L g20754 ( 
.A(n_20684),
.B(n_7542),
.C(n_7525),
.Y(n_20754)
);

NAND3xp33_ASAP7_75t_L g20755 ( 
.A(n_20724),
.B(n_6812),
.C(n_6225),
.Y(n_20755)
);

INVx1_ASAP7_75t_L g20756 ( 
.A(n_20710),
.Y(n_20756)
);

NOR4xp25_ASAP7_75t_L g20757 ( 
.A(n_20723),
.B(n_7617),
.C(n_7618),
.D(n_7612),
.Y(n_20757)
);

NOR3xp33_ASAP7_75t_L g20758 ( 
.A(n_20670),
.B(n_7542),
.C(n_7525),
.Y(n_20758)
);

AO21x1_ASAP7_75t_L g20759 ( 
.A1(n_20697),
.A2(n_9573),
.B(n_9572),
.Y(n_20759)
);

BUFx6f_ASAP7_75t_L g20760 ( 
.A(n_20677),
.Y(n_20760)
);

NOR3xp33_ASAP7_75t_SL g20761 ( 
.A(n_20713),
.B(n_7618),
.C(n_7617),
.Y(n_20761)
);

AND4x1_ASAP7_75t_L g20762 ( 
.A(n_20701),
.B(n_20641),
.C(n_20705),
.D(n_20716),
.Y(n_20762)
);

HB1xp67_ASAP7_75t_L g20763 ( 
.A(n_20674),
.Y(n_20763)
);

OR5x1_ASAP7_75t_L g20764 ( 
.A(n_20690),
.B(n_7512),
.C(n_7424),
.D(n_7301),
.E(n_9191),
.Y(n_20764)
);

NAND5xp2_ASAP7_75t_L g20765 ( 
.A(n_20680),
.B(n_4622),
.C(n_7301),
.D(n_7512),
.E(n_7424),
.Y(n_20765)
);

NAND4xp25_ASAP7_75t_L g20766 ( 
.A(n_20706),
.B(n_5717),
.C(n_7061),
.D(n_6942),
.Y(n_20766)
);

OAI211xp5_ASAP7_75t_L g20767 ( 
.A1(n_20667),
.A2(n_7957),
.B(n_5605),
.C(n_5608),
.Y(n_20767)
);

NAND3xp33_ASAP7_75t_L g20768 ( 
.A(n_20696),
.B(n_6812),
.C(n_6225),
.Y(n_20768)
);

OR2x2_ASAP7_75t_L g20769 ( 
.A(n_20687),
.B(n_8673),
.Y(n_20769)
);

NOR4xp25_ASAP7_75t_L g20770 ( 
.A(n_20719),
.B(n_7618),
.C(n_7628),
.D(n_7617),
.Y(n_20770)
);

NAND2x1_ASAP7_75t_SL g20771 ( 
.A(n_20646),
.B(n_8070),
.Y(n_20771)
);

OR5x1_ASAP7_75t_L g20772 ( 
.A(n_20715),
.B(n_20648),
.C(n_20699),
.D(n_20722),
.E(n_20709),
.Y(n_20772)
);

HB1xp67_ASAP7_75t_L g20773 ( 
.A(n_20695),
.Y(n_20773)
);

NAND4xp25_ASAP7_75t_SL g20774 ( 
.A(n_20694),
.B(n_8125),
.C(n_7638),
.D(n_7643),
.Y(n_20774)
);

NAND5xp2_ASAP7_75t_L g20775 ( 
.A(n_20639),
.B(n_7512),
.C(n_7424),
.D(n_6033),
.E(n_7553),
.Y(n_20775)
);

NAND4xp25_ASAP7_75t_L g20776 ( 
.A(n_20627),
.B(n_7061),
.C(n_7085),
.D(n_6942),
.Y(n_20776)
);

OAI22xp5_ASAP7_75t_L g20777 ( 
.A1(n_20675),
.A2(n_8094),
.B1(n_8070),
.B2(n_8125),
.Y(n_20777)
);

NOR4xp75_ASAP7_75t_L g20778 ( 
.A(n_20650),
.B(n_7173),
.C(n_7267),
.D(n_7156),
.Y(n_20778)
);

OR2x2_ASAP7_75t_L g20779 ( 
.A(n_20676),
.B(n_8673),
.Y(n_20779)
);

NAND4xp75_ASAP7_75t_L g20780 ( 
.A(n_20655),
.B(n_6711),
.C(n_6774),
.D(n_6709),
.Y(n_20780)
);

NOR4xp75_ASAP7_75t_L g20781 ( 
.A(n_20702),
.B(n_7173),
.C(n_7267),
.D(n_7156),
.Y(n_20781)
);

INVx2_ASAP7_75t_L g20782 ( 
.A(n_20665),
.Y(n_20782)
);

AOI31xp33_ASAP7_75t_L g20783 ( 
.A1(n_20700),
.A2(n_5773),
.A3(n_5775),
.B(n_5746),
.Y(n_20783)
);

NOR4xp25_ASAP7_75t_L g20784 ( 
.A(n_20649),
.B(n_7638),
.C(n_7643),
.D(n_7628),
.Y(n_20784)
);

NOR3xp33_ASAP7_75t_L g20785 ( 
.A(n_20698),
.B(n_7552),
.C(n_7542),
.Y(n_20785)
);

NAND3x1_ASAP7_75t_L g20786 ( 
.A(n_20711),
.B(n_5680),
.C(n_5673),
.Y(n_20786)
);

OAI211xp5_ASAP7_75t_SL g20787 ( 
.A1(n_20659),
.A2(n_5673),
.B(n_5685),
.C(n_5680),
.Y(n_20787)
);

OR3x2_ASAP7_75t_L g20788 ( 
.A(n_20721),
.B(n_8082),
.C(n_7638),
.Y(n_20788)
);

NOR3xp33_ASAP7_75t_SL g20789 ( 
.A(n_20669),
.B(n_20703),
.C(n_20686),
.Y(n_20789)
);

HB1xp67_ASAP7_75t_L g20790 ( 
.A(n_20673),
.Y(n_20790)
);

NAND4xp25_ASAP7_75t_L g20791 ( 
.A(n_20682),
.B(n_7061),
.C(n_7264),
.D(n_7085),
.Y(n_20791)
);

AOI22xp33_ASAP7_75t_L g20792 ( 
.A1(n_20661),
.A2(n_20653),
.B1(n_20635),
.B2(n_20672),
.Y(n_20792)
);

NOR3xp33_ASAP7_75t_SL g20793 ( 
.A(n_20693),
.B(n_7643),
.C(n_7628),
.Y(n_20793)
);

OR2x2_ASAP7_75t_L g20794 ( 
.A(n_20683),
.B(n_8673),
.Y(n_20794)
);

NAND5xp2_ASAP7_75t_L g20795 ( 
.A(n_20717),
.B(n_7512),
.C(n_6033),
.D(n_7553),
.E(n_5622),
.Y(n_20795)
);

NOR3xp33_ASAP7_75t_L g20796 ( 
.A(n_20689),
.B(n_7552),
.C(n_7542),
.Y(n_20796)
);

NAND4xp75_ASAP7_75t_L g20797 ( 
.A(n_20658),
.B(n_6863),
.C(n_6891),
.D(n_6774),
.Y(n_20797)
);

OAI211xp5_ASAP7_75t_SL g20798 ( 
.A1(n_20714),
.A2(n_20671),
.B(n_20660),
.C(n_20720),
.Y(n_20798)
);

NOR2x1_ASAP7_75t_L g20799 ( 
.A(n_20652),
.B(n_7085),
.Y(n_20799)
);

NOR2x1_ASAP7_75t_L g20800 ( 
.A(n_20657),
.B(n_7085),
.Y(n_20800)
);

NAND4xp75_ASAP7_75t_L g20801 ( 
.A(n_20720),
.B(n_6891),
.C(n_6911),
.D(n_6863),
.Y(n_20801)
);

NAND3x1_ASAP7_75t_L g20802 ( 
.A(n_20692),
.B(n_5704),
.C(n_5685),
.Y(n_20802)
);

NOR5xp2_ASAP7_75t_L g20803 ( 
.A(n_20685),
.B(n_7656),
.C(n_7668),
.D(n_7651),
.E(n_7648),
.Y(n_20803)
);

INVxp33_ASAP7_75t_SL g20804 ( 
.A(n_20640),
.Y(n_20804)
);

OR2x2_ASAP7_75t_L g20805 ( 
.A(n_20632),
.B(n_8673),
.Y(n_20805)
);

NOR3xp33_ASAP7_75t_SL g20806 ( 
.A(n_20681),
.B(n_20642),
.C(n_20651),
.Y(n_20806)
);

NOR3xp33_ASAP7_75t_L g20807 ( 
.A(n_20642),
.B(n_7604),
.C(n_7552),
.Y(n_20807)
);

NAND4xp25_ASAP7_75t_SL g20808 ( 
.A(n_20634),
.B(n_7651),
.C(n_7656),
.D(n_7648),
.Y(n_20808)
);

HB1xp67_ASAP7_75t_L g20809 ( 
.A(n_20630),
.Y(n_20809)
);

NOR3xp33_ASAP7_75t_L g20810 ( 
.A(n_20630),
.B(n_7604),
.C(n_7552),
.Y(n_20810)
);

INVx1_ASAP7_75t_L g20811 ( 
.A(n_20630),
.Y(n_20811)
);

OAI211xp5_ASAP7_75t_SL g20812 ( 
.A1(n_20630),
.A2(n_5685),
.B(n_5704),
.C(n_7648),
.Y(n_20812)
);

AND4x1_ASAP7_75t_L g20813 ( 
.A(n_20634),
.B(n_7176),
.C(n_7188),
.D(n_7058),
.Y(n_20813)
);

AND3x2_ASAP7_75t_L g20814 ( 
.A(n_20634),
.B(n_5773),
.C(n_5746),
.Y(n_20814)
);

INVxp67_ASAP7_75t_L g20815 ( 
.A(n_20630),
.Y(n_20815)
);

OR2x2_ASAP7_75t_L g20816 ( 
.A(n_20630),
.B(n_8673),
.Y(n_20816)
);

OR3x2_ASAP7_75t_L g20817 ( 
.A(n_20634),
.B(n_8082),
.C(n_7656),
.Y(n_20817)
);

NOR3xp33_ASAP7_75t_L g20818 ( 
.A(n_20630),
.B(n_7604),
.C(n_7552),
.Y(n_20818)
);

AND2x4_ASAP7_75t_L g20819 ( 
.A(n_20630),
.B(n_7553),
.Y(n_20819)
);

NAND4xp75_ASAP7_75t_L g20820 ( 
.A(n_20630),
.B(n_6891),
.C(n_6911),
.D(n_6863),
.Y(n_20820)
);

NAND3xp33_ASAP7_75t_SL g20821 ( 
.A(n_20634),
.B(n_7604),
.C(n_7552),
.Y(n_20821)
);

NAND5xp2_ASAP7_75t_L g20822 ( 
.A(n_20756),
.B(n_7512),
.C(n_6033),
.D(n_5634),
.E(n_5652),
.Y(n_20822)
);

NAND4xp25_ASAP7_75t_SL g20823 ( 
.A(n_20811),
.B(n_7668),
.C(n_7689),
.D(n_7651),
.Y(n_20823)
);

AOI222xp33_ASAP7_75t_L g20824 ( 
.A1(n_20815),
.A2(n_20809),
.B1(n_20760),
.B2(n_20763),
.C1(n_20732),
.C2(n_20790),
.Y(n_20824)
);

INVx2_ASAP7_75t_SL g20825 ( 
.A(n_20725),
.Y(n_20825)
);

NOR3xp33_ASAP7_75t_L g20826 ( 
.A(n_20753),
.B(n_7639),
.C(n_7604),
.Y(n_20826)
);

NOR3xp33_ASAP7_75t_L g20827 ( 
.A(n_20726),
.B(n_7639),
.C(n_7604),
.Y(n_20827)
);

NAND3xp33_ASAP7_75t_L g20828 ( 
.A(n_20760),
.B(n_6812),
.C(n_4540),
.Y(n_20828)
);

OAI211xp5_ASAP7_75t_L g20829 ( 
.A1(n_20760),
.A2(n_7704),
.B(n_7728),
.C(n_7639),
.Y(n_20829)
);

NAND2xp5_ASAP7_75t_L g20830 ( 
.A(n_20773),
.B(n_9191),
.Y(n_20830)
);

NOR2x1_ASAP7_75t_L g20831 ( 
.A(n_20782),
.B(n_20727),
.Y(n_20831)
);

AOI222xp33_ASAP7_75t_L g20832 ( 
.A1(n_20745),
.A2(n_7553),
.B1(n_7871),
.B2(n_7909),
.C1(n_7866),
.C2(n_7739),
.Y(n_20832)
);

AND2x4_ASAP7_75t_L g20833 ( 
.A(n_20762),
.B(n_7553),
.Y(n_20833)
);

INVx2_ASAP7_75t_L g20834 ( 
.A(n_20772),
.Y(n_20834)
);

NOR3xp33_ASAP7_75t_L g20835 ( 
.A(n_20798),
.B(n_7704),
.C(n_7639),
.Y(n_20835)
);

AND2x4_ASAP7_75t_L g20836 ( 
.A(n_20806),
.B(n_7553),
.Y(n_20836)
);

NAND4xp25_ASAP7_75t_L g20837 ( 
.A(n_20792),
.B(n_7361),
.C(n_7383),
.D(n_7264),
.Y(n_20837)
);

NAND2x1p5_ASAP7_75t_L g20838 ( 
.A(n_20751),
.B(n_5545),
.Y(n_20838)
);

NOR4xp25_ASAP7_75t_L g20839 ( 
.A(n_20769),
.B(n_7689),
.C(n_7691),
.D(n_7668),
.Y(n_20839)
);

NOR2x1p5_ASAP7_75t_L g20840 ( 
.A(n_20730),
.B(n_7264),
.Y(n_20840)
);

NAND4xp25_ASAP7_75t_L g20841 ( 
.A(n_20804),
.B(n_7361),
.C(n_7383),
.D(n_7264),
.Y(n_20841)
);

AOI22xp33_ASAP7_75t_L g20842 ( 
.A1(n_20738),
.A2(n_20788),
.B1(n_20807),
.B2(n_20779),
.Y(n_20842)
);

NOR2x1_ASAP7_75t_L g20843 ( 
.A(n_20794),
.B(n_8700),
.Y(n_20843)
);

AOI22xp5_ASAP7_75t_L g20844 ( 
.A1(n_20789),
.A2(n_7512),
.B1(n_5605),
.B2(n_5608),
.Y(n_20844)
);

OAI22xp33_ASAP7_75t_L g20845 ( 
.A1(n_20805),
.A2(n_5545),
.B1(n_5608),
.B2(n_5605),
.Y(n_20845)
);

INVx1_ASAP7_75t_L g20846 ( 
.A(n_20771),
.Y(n_20846)
);

NOR2x1_ASAP7_75t_L g20847 ( 
.A(n_20799),
.B(n_8700),
.Y(n_20847)
);

NOR4xp25_ASAP7_75t_L g20848 ( 
.A(n_20786),
.B(n_7691),
.C(n_7693),
.D(n_7689),
.Y(n_20848)
);

AND4x1_ASAP7_75t_L g20849 ( 
.A(n_20784),
.B(n_7512),
.C(n_7188),
.D(n_7189),
.Y(n_20849)
);

NAND5xp2_ASAP7_75t_L g20850 ( 
.A(n_20796),
.B(n_6033),
.C(n_5634),
.D(n_5652),
.E(n_5495),
.Y(n_20850)
);

INVx3_ASAP7_75t_L g20851 ( 
.A(n_20802),
.Y(n_20851)
);

AOI32xp33_ASAP7_75t_L g20852 ( 
.A1(n_20800),
.A2(n_9421),
.A3(n_8693),
.B1(n_7728),
.B2(n_7764),
.Y(n_20852)
);

INVx1_ASAP7_75t_L g20853 ( 
.A(n_20781),
.Y(n_20853)
);

AND3x4_ASAP7_75t_L g20854 ( 
.A(n_20785),
.B(n_7383),
.C(n_7361),
.Y(n_20854)
);

NAND4xp25_ASAP7_75t_L g20855 ( 
.A(n_20795),
.B(n_7383),
.C(n_7514),
.D(n_7361),
.Y(n_20855)
);

NAND3xp33_ASAP7_75t_L g20856 ( 
.A(n_20787),
.B(n_20793),
.C(n_20761),
.Y(n_20856)
);

OAI211xp5_ASAP7_75t_SL g20857 ( 
.A1(n_20733),
.A2(n_5704),
.B(n_7693),
.C(n_7691),
.Y(n_20857)
);

AND2x2_ASAP7_75t_L g20858 ( 
.A(n_20816),
.B(n_8673),
.Y(n_20858)
);

OAI211xp5_ASAP7_75t_L g20859 ( 
.A1(n_20752),
.A2(n_7704),
.B(n_7728),
.C(n_7639),
.Y(n_20859)
);

A2O1A1Ixp33_ASAP7_75t_L g20860 ( 
.A1(n_20737),
.A2(n_8478),
.B(n_8491),
.C(n_8472),
.Y(n_20860)
);

AND2x4_ASAP7_75t_L g20861 ( 
.A(n_20778),
.B(n_8202),
.Y(n_20861)
);

AND2x4_ASAP7_75t_L g20862 ( 
.A(n_20750),
.B(n_20755),
.Y(n_20862)
);

OAI221xp5_ASAP7_75t_L g20863 ( 
.A1(n_20742),
.A2(n_5608),
.B1(n_5621),
.B2(n_5605),
.C(n_5545),
.Y(n_20863)
);

AND4x1_ASAP7_75t_L g20864 ( 
.A(n_20748),
.B(n_7176),
.C(n_7189),
.D(n_7188),
.Y(n_20864)
);

NOR3xp33_ASAP7_75t_L g20865 ( 
.A(n_20734),
.B(n_7704),
.C(n_7639),
.Y(n_20865)
);

OAI211xp5_ASAP7_75t_L g20866 ( 
.A1(n_20791),
.A2(n_7728),
.B(n_7764),
.C(n_7704),
.Y(n_20866)
);

XOR2xp5_ASAP7_75t_L g20867 ( 
.A(n_20817),
.B(n_4532),
.Y(n_20867)
);

INVx1_ASAP7_75t_L g20868 ( 
.A(n_20741),
.Y(n_20868)
);

OAI22xp5_ASAP7_75t_L g20869 ( 
.A1(n_20749),
.A2(n_8094),
.B1(n_8070),
.B2(n_8069),
.Y(n_20869)
);

OAI221xp5_ASAP7_75t_L g20870 ( 
.A1(n_20739),
.A2(n_5608),
.B1(n_5621),
.B2(n_5605),
.C(n_5545),
.Y(n_20870)
);

AOI211xp5_ASAP7_75t_L g20871 ( 
.A1(n_20774),
.A2(n_4532),
.B(n_4581),
.C(n_4540),
.Y(n_20871)
);

AOI22xp5_ASAP7_75t_L g20872 ( 
.A1(n_20821),
.A2(n_5605),
.B1(n_5608),
.B2(n_5545),
.Y(n_20872)
);

NAND2xp5_ASAP7_75t_L g20873 ( 
.A(n_20801),
.B(n_8336),
.Y(n_20873)
);

NAND4xp25_ASAP7_75t_SL g20874 ( 
.A(n_20754),
.B(n_7695),
.C(n_7696),
.D(n_7693),
.Y(n_20874)
);

NOR2xp33_ASAP7_75t_L g20875 ( 
.A(n_20783),
.B(n_7380),
.Y(n_20875)
);

INVxp33_ASAP7_75t_L g20876 ( 
.A(n_20780),
.Y(n_20876)
);

AOI22xp5_ASAP7_75t_L g20877 ( 
.A1(n_20768),
.A2(n_5605),
.B1(n_5608),
.B2(n_5545),
.Y(n_20877)
);

INVx1_ASAP7_75t_L g20878 ( 
.A(n_20814),
.Y(n_20878)
);

NOR3xp33_ASAP7_75t_L g20879 ( 
.A(n_20775),
.B(n_7728),
.C(n_7704),
.Y(n_20879)
);

AND2x2_ASAP7_75t_SL g20880 ( 
.A(n_20803),
.B(n_5605),
.Y(n_20880)
);

OAI22xp5_ASAP7_75t_L g20881 ( 
.A1(n_20797),
.A2(n_8094),
.B1(n_8070),
.B2(n_8069),
.Y(n_20881)
);

NAND3xp33_ASAP7_75t_L g20882 ( 
.A(n_20777),
.B(n_6812),
.C(n_4540),
.Y(n_20882)
);

NAND4xp25_ASAP7_75t_L g20883 ( 
.A(n_20758),
.B(n_7559),
.C(n_7576),
.D(n_7514),
.Y(n_20883)
);

AND2x2_ASAP7_75t_L g20884 ( 
.A(n_20813),
.B(n_8336),
.Y(n_20884)
);

INVx1_ASAP7_75t_L g20885 ( 
.A(n_20812),
.Y(n_20885)
);

INVx1_ASAP7_75t_L g20886 ( 
.A(n_20759),
.Y(n_20886)
);

AOI22xp5_ASAP7_75t_L g20887 ( 
.A1(n_20767),
.A2(n_5621),
.B1(n_5629),
.B2(n_5608),
.Y(n_20887)
);

NAND4xp25_ASAP7_75t_L g20888 ( 
.A(n_20746),
.B(n_7559),
.C(n_7576),
.D(n_7514),
.Y(n_20888)
);

NAND2xp5_ASAP7_75t_L g20889 ( 
.A(n_20731),
.B(n_8336),
.Y(n_20889)
);

INVx1_ASAP7_75t_L g20890 ( 
.A(n_20770),
.Y(n_20890)
);

NAND3x1_ASAP7_75t_L g20891 ( 
.A(n_20764),
.B(n_5704),
.C(n_7173),
.Y(n_20891)
);

AOI311xp33_ASAP7_75t_L g20892 ( 
.A1(n_20744),
.A2(n_7699),
.A3(n_7701),
.B(n_7696),
.C(n_7695),
.Y(n_20892)
);

AOI22xp33_ASAP7_75t_L g20893 ( 
.A1(n_20810),
.A2(n_7074),
.B1(n_7240),
.B2(n_7053),
.Y(n_20893)
);

INVxp67_ASAP7_75t_L g20894 ( 
.A(n_20765),
.Y(n_20894)
);

OAI22xp5_ASAP7_75t_L g20895 ( 
.A1(n_20736),
.A2(n_8094),
.B1(n_8070),
.B2(n_8069),
.Y(n_20895)
);

AO22x1_ASAP7_75t_L g20896 ( 
.A1(n_20818),
.A2(n_4779),
.B1(n_4863),
.B2(n_4713),
.Y(n_20896)
);

XNOR2xp5_ASAP7_75t_L g20897 ( 
.A(n_20776),
.B(n_8336),
.Y(n_20897)
);

AOI221xp5_ASAP7_75t_L g20898 ( 
.A1(n_20728),
.A2(n_8002),
.B1(n_8021),
.B2(n_7995),
.C(n_7976),
.Y(n_20898)
);

NAND4xp25_ASAP7_75t_L g20899 ( 
.A(n_20740),
.B(n_7559),
.C(n_7576),
.D(n_7514),
.Y(n_20899)
);

AOI22xp5_ASAP7_75t_L g20900 ( 
.A1(n_20825),
.A2(n_20766),
.B1(n_20808),
.B2(n_20735),
.Y(n_20900)
);

HB1xp67_ASAP7_75t_L g20901 ( 
.A(n_20834),
.Y(n_20901)
);

AOI22xp33_ASAP7_75t_L g20902 ( 
.A1(n_20824),
.A2(n_20735),
.B1(n_20729),
.B2(n_20747),
.Y(n_20902)
);

INVx3_ASAP7_75t_L g20903 ( 
.A(n_20846),
.Y(n_20903)
);

NAND2xp5_ASAP7_75t_L g20904 ( 
.A(n_20831),
.B(n_20757),
.Y(n_20904)
);

AND2x4_ASAP7_75t_L g20905 ( 
.A(n_20894),
.B(n_20747),
.Y(n_20905)
);

AND3x4_ASAP7_75t_L g20906 ( 
.A(n_20862),
.B(n_20879),
.C(n_20835),
.Y(n_20906)
);

NAND2xp5_ASAP7_75t_L g20907 ( 
.A(n_20842),
.B(n_20743),
.Y(n_20907)
);

INVx1_ASAP7_75t_L g20908 ( 
.A(n_20890),
.Y(n_20908)
);

INVx1_ASAP7_75t_L g20909 ( 
.A(n_20886),
.Y(n_20909)
);

NOR2xp67_ASAP7_75t_SL g20910 ( 
.A(n_20878),
.B(n_20820),
.Y(n_20910)
);

AOI22xp33_ASAP7_75t_L g20911 ( 
.A1(n_20853),
.A2(n_20819),
.B1(n_7074),
.B2(n_7240),
.Y(n_20911)
);

OAI22x1_ASAP7_75t_L g20912 ( 
.A1(n_20868),
.A2(n_20851),
.B1(n_20856),
.B2(n_20885),
.Y(n_20912)
);

AND2x4_ASAP7_75t_L g20913 ( 
.A(n_20862),
.B(n_20819),
.Y(n_20913)
);

NOR4xp25_ASAP7_75t_SL g20914 ( 
.A(n_20857),
.B(n_7696),
.C(n_7699),
.D(n_7695),
.Y(n_20914)
);

NAND2x1p5_ASAP7_75t_L g20915 ( 
.A(n_20840),
.B(n_5621),
.Y(n_20915)
);

AOI22xp5_ASAP7_75t_L g20916 ( 
.A1(n_20876),
.A2(n_5629),
.B1(n_5661),
.B2(n_5621),
.Y(n_20916)
);

AO22x2_ASAP7_75t_L g20917 ( 
.A1(n_20867),
.A2(n_8094),
.B1(n_7764),
.B2(n_7766),
.Y(n_20917)
);

AOI21xp33_ASAP7_75t_SL g20918 ( 
.A1(n_20838),
.A2(n_8365),
.B(n_8336),
.Y(n_20918)
);

INVx2_ASAP7_75t_L g20919 ( 
.A(n_20880),
.Y(n_20919)
);

NOR2x1_ASAP7_75t_L g20920 ( 
.A(n_20889),
.B(n_20897),
.Y(n_20920)
);

INVx1_ASAP7_75t_L g20921 ( 
.A(n_20891),
.Y(n_20921)
);

OAI22x1_ASAP7_75t_L g20922 ( 
.A1(n_20849),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_20922)
);

NOR2x1_ASAP7_75t_L g20923 ( 
.A(n_20845),
.B(n_8700),
.Y(n_20923)
);

INVx1_ASAP7_75t_L g20924 ( 
.A(n_20884),
.Y(n_20924)
);

NOR3xp33_ASAP7_75t_L g20925 ( 
.A(n_20875),
.B(n_7764),
.C(n_7728),
.Y(n_20925)
);

OAI21xp5_ASAP7_75t_L g20926 ( 
.A1(n_20843),
.A2(n_9421),
.B(n_8592),
.Y(n_20926)
);

INVx1_ASAP7_75t_L g20927 ( 
.A(n_20861),
.Y(n_20927)
);

NAND3xp33_ASAP7_75t_L g20928 ( 
.A(n_20827),
.B(n_4540),
.C(n_4532),
.Y(n_20928)
);

NOR2xp67_ASAP7_75t_SL g20929 ( 
.A(n_20882),
.B(n_5621),
.Y(n_20929)
);

INVx1_ASAP7_75t_SL g20930 ( 
.A(n_20836),
.Y(n_20930)
);

INVx1_ASAP7_75t_L g20931 ( 
.A(n_20873),
.Y(n_20931)
);

NOR2xp33_ASAP7_75t_L g20932 ( 
.A(n_20836),
.B(n_7387),
.Y(n_20932)
);

NAND2xp5_ASAP7_75t_L g20933 ( 
.A(n_20839),
.B(n_8365),
.Y(n_20933)
);

INVx2_ASAP7_75t_L g20934 ( 
.A(n_20858),
.Y(n_20934)
);

NOR2xp67_ASAP7_75t_L g20935 ( 
.A(n_20899),
.B(n_20855),
.Y(n_20935)
);

OAI21xp5_ASAP7_75t_L g20936 ( 
.A1(n_20859),
.A2(n_8592),
.B(n_8585),
.Y(n_20936)
);

NAND3x1_ASAP7_75t_L g20937 ( 
.A(n_20847),
.B(n_5704),
.C(n_7276),
.Y(n_20937)
);

INVx3_ASAP7_75t_SL g20938 ( 
.A(n_20833),
.Y(n_20938)
);

AND3x4_ASAP7_75t_L g20939 ( 
.A(n_20864),
.B(n_7576),
.C(n_7559),
.Y(n_20939)
);

XNOR2x1_ASAP7_75t_L g20940 ( 
.A(n_20854),
.B(n_8365),
.Y(n_20940)
);

INVx1_ASAP7_75t_L g20941 ( 
.A(n_20848),
.Y(n_20941)
);

AOI22xp33_ASAP7_75t_L g20942 ( 
.A1(n_20833),
.A2(n_7074),
.B1(n_7240),
.B2(n_7053),
.Y(n_20942)
);

NAND2xp5_ASAP7_75t_L g20943 ( 
.A(n_20871),
.B(n_8365),
.Y(n_20943)
);

AOI211xp5_ASAP7_75t_L g20944 ( 
.A1(n_20866),
.A2(n_20888),
.B(n_20850),
.C(n_20870),
.Y(n_20944)
);

NOR4xp75_ASAP7_75t_L g20945 ( 
.A(n_20863),
.B(n_7276),
.C(n_7303),
.D(n_7302),
.Y(n_20945)
);

AOI222xp33_ASAP7_75t_L g20946 ( 
.A1(n_20869),
.A2(n_20830),
.B1(n_20896),
.B2(n_20828),
.C1(n_20881),
.C2(n_20895),
.Y(n_20946)
);

NAND4xp25_ASAP7_75t_L g20947 ( 
.A(n_20892),
.B(n_7665),
.C(n_7687),
.D(n_7600),
.Y(n_20947)
);

OAI32xp33_ASAP7_75t_L g20948 ( 
.A1(n_20865),
.A2(n_8082),
.A3(n_7303),
.B1(n_7315),
.B2(n_7302),
.Y(n_20948)
);

HB1xp67_ASAP7_75t_L g20949 ( 
.A(n_20874),
.Y(n_20949)
);

NAND4xp75_ASAP7_75t_L g20950 ( 
.A(n_20844),
.B(n_6911),
.C(n_7189),
.D(n_7176),
.Y(n_20950)
);

INVx1_ASAP7_75t_L g20951 ( 
.A(n_20822),
.Y(n_20951)
);

OAI221xp5_ASAP7_75t_L g20952 ( 
.A1(n_20826),
.A2(n_4540),
.B1(n_4618),
.B2(n_4614),
.C(n_4581),
.Y(n_20952)
);

OAI221xp5_ASAP7_75t_L g20953 ( 
.A1(n_20872),
.A2(n_4540),
.B1(n_4618),
.B2(n_4614),
.C(n_4581),
.Y(n_20953)
);

INVx4_ASAP7_75t_L g20954 ( 
.A(n_20883),
.Y(n_20954)
);

NOR2xp33_ASAP7_75t_R g20955 ( 
.A(n_20893),
.B(n_5621),
.Y(n_20955)
);

INVx2_ASAP7_75t_L g20956 ( 
.A(n_20877),
.Y(n_20956)
);

XNOR2xp5_ASAP7_75t_L g20957 ( 
.A(n_20829),
.B(n_8365),
.Y(n_20957)
);

INVx1_ASAP7_75t_L g20958 ( 
.A(n_20887),
.Y(n_20958)
);

BUFx2_ASAP7_75t_L g20959 ( 
.A(n_20898),
.Y(n_20959)
);

INVx1_ASAP7_75t_L g20960 ( 
.A(n_20823),
.Y(n_20960)
);

AO22x2_ASAP7_75t_L g20961 ( 
.A1(n_20852),
.A2(n_7766),
.B1(n_7801),
.B2(n_7764),
.Y(n_20961)
);

INVx1_ASAP7_75t_SL g20962 ( 
.A(n_20832),
.Y(n_20962)
);

INVx1_ASAP7_75t_L g20963 ( 
.A(n_20901),
.Y(n_20963)
);

AO22x2_ASAP7_75t_L g20964 ( 
.A1(n_20908),
.A2(n_20837),
.B1(n_20841),
.B2(n_20860),
.Y(n_20964)
);

OAI22xp5_ASAP7_75t_L g20965 ( 
.A1(n_20903),
.A2(n_8803),
.B1(n_8876),
.B2(n_8700),
.Y(n_20965)
);

INVxp67_ASAP7_75t_L g20966 ( 
.A(n_20912),
.Y(n_20966)
);

NAND2xp5_ASAP7_75t_L g20967 ( 
.A(n_20909),
.B(n_7739),
.Y(n_20967)
);

INVx1_ASAP7_75t_L g20968 ( 
.A(n_20904),
.Y(n_20968)
);

AO22x2_ASAP7_75t_L g20969 ( 
.A1(n_20906),
.A2(n_20927),
.B1(n_20919),
.B2(n_20941),
.Y(n_20969)
);

XNOR2x1_ASAP7_75t_L g20970 ( 
.A(n_20920),
.B(n_8585),
.Y(n_20970)
);

INVx1_ASAP7_75t_L g20971 ( 
.A(n_20905),
.Y(n_20971)
);

HB1xp67_ASAP7_75t_L g20972 ( 
.A(n_20934),
.Y(n_20972)
);

INVx1_ASAP7_75t_L g20973 ( 
.A(n_20913),
.Y(n_20973)
);

INVxp67_ASAP7_75t_L g20974 ( 
.A(n_20924),
.Y(n_20974)
);

INVx2_ASAP7_75t_L g20975 ( 
.A(n_20951),
.Y(n_20975)
);

INVx2_ASAP7_75t_L g20976 ( 
.A(n_20921),
.Y(n_20976)
);

INVx1_ASAP7_75t_L g20977 ( 
.A(n_20935),
.Y(n_20977)
);

INVx1_ASAP7_75t_L g20978 ( 
.A(n_20900),
.Y(n_20978)
);

OAI22xp5_ASAP7_75t_L g20979 ( 
.A1(n_20902),
.A2(n_8876),
.B1(n_8962),
.B2(n_8700),
.Y(n_20979)
);

NOR2xp33_ASAP7_75t_L g20980 ( 
.A(n_20938),
.B(n_5621),
.Y(n_20980)
);

NOR2xp33_ASAP7_75t_L g20981 ( 
.A(n_20930),
.B(n_5629),
.Y(n_20981)
);

INVx1_ASAP7_75t_L g20982 ( 
.A(n_20907),
.Y(n_20982)
);

INVx2_ASAP7_75t_L g20983 ( 
.A(n_20954),
.Y(n_20983)
);

INVx1_ASAP7_75t_L g20984 ( 
.A(n_20959),
.Y(n_20984)
);

INVx5_ASAP7_75t_L g20985 ( 
.A(n_20931),
.Y(n_20985)
);

XNOR2x1_ASAP7_75t_L g20986 ( 
.A(n_20962),
.B(n_8365),
.Y(n_20986)
);

INVx1_ASAP7_75t_L g20987 ( 
.A(n_20949),
.Y(n_20987)
);

OA22x2_ASAP7_75t_L g20988 ( 
.A1(n_20960),
.A2(n_8496),
.B1(n_8491),
.B2(n_8748),
.Y(n_20988)
);

OAI211xp5_ASAP7_75t_L g20989 ( 
.A1(n_20958),
.A2(n_4540),
.B(n_4614),
.C(n_4581),
.Y(n_20989)
);

INVx2_ASAP7_75t_L g20990 ( 
.A(n_20956),
.Y(n_20990)
);

AO22x2_ASAP7_75t_L g20991 ( 
.A1(n_20910),
.A2(n_7766),
.B1(n_7801),
.B2(n_7764),
.Y(n_20991)
);

AOI22xp33_ASAP7_75t_L g20992 ( 
.A1(n_20915),
.A2(n_7388),
.B1(n_7396),
.B2(n_7387),
.Y(n_20992)
);

AO22x2_ASAP7_75t_L g20993 ( 
.A1(n_20940),
.A2(n_7801),
.B1(n_7927),
.B2(n_7766),
.Y(n_20993)
);

INVx1_ASAP7_75t_L g20994 ( 
.A(n_20944),
.Y(n_20994)
);

AND3x4_ASAP7_75t_L g20995 ( 
.A(n_20925),
.B(n_5773),
.C(n_5746),
.Y(n_20995)
);

INVx1_ASAP7_75t_L g20996 ( 
.A(n_20946),
.Y(n_20996)
);

AOI22xp5_ASAP7_75t_L g20997 ( 
.A1(n_20932),
.A2(n_4540),
.B1(n_4614),
.B2(n_4581),
.Y(n_20997)
);

INVx1_ASAP7_75t_L g20998 ( 
.A(n_20957),
.Y(n_20998)
);

INVx2_ASAP7_75t_L g20999 ( 
.A(n_20937),
.Y(n_20999)
);

XOR2xp5_ASAP7_75t_L g21000 ( 
.A(n_20933),
.B(n_20961),
.Y(n_21000)
);

INVx1_ASAP7_75t_L g21001 ( 
.A(n_20929),
.Y(n_21001)
);

INVx1_ASAP7_75t_L g21002 ( 
.A(n_20955),
.Y(n_21002)
);

INVx1_ASAP7_75t_L g21003 ( 
.A(n_20943),
.Y(n_21003)
);

INVx1_ASAP7_75t_L g21004 ( 
.A(n_20961),
.Y(n_21004)
);

OAI22xp5_ASAP7_75t_L g21005 ( 
.A1(n_20939),
.A2(n_8962),
.B1(n_8876),
.B2(n_7616),
.Y(n_21005)
);

INVx1_ASAP7_75t_L g21006 ( 
.A(n_20947),
.Y(n_21006)
);

BUFx2_ASAP7_75t_L g21007 ( 
.A(n_20966),
.Y(n_21007)
);

BUFx2_ASAP7_75t_L g21008 ( 
.A(n_20975),
.Y(n_21008)
);

AOI21xp5_ASAP7_75t_L g21009 ( 
.A1(n_20963),
.A2(n_20914),
.B(n_20922),
.Y(n_21009)
);

INVx1_ASAP7_75t_L g21010 ( 
.A(n_20972),
.Y(n_21010)
);

INVx2_ASAP7_75t_SL g21011 ( 
.A(n_20985),
.Y(n_21011)
);

CKINVDCx20_ASAP7_75t_R g21012 ( 
.A(n_20973),
.Y(n_21012)
);

OAI22x1_ASAP7_75t_L g21013 ( 
.A1(n_20990),
.A2(n_20928),
.B1(n_20923),
.B2(n_20916),
.Y(n_21013)
);

INVx1_ASAP7_75t_SL g21014 ( 
.A(n_20996),
.Y(n_21014)
);

AOI222xp33_ASAP7_75t_L g21015 ( 
.A1(n_20984),
.A2(n_20974),
.B1(n_20971),
.B2(n_20987),
.C1(n_20985),
.C2(n_20968),
.Y(n_21015)
);

INVxp67_ASAP7_75t_L g21016 ( 
.A(n_20969),
.Y(n_21016)
);

NOR2xp67_ASAP7_75t_L g21017 ( 
.A(n_20983),
.B(n_20926),
.Y(n_21017)
);

INVx1_ASAP7_75t_L g21018 ( 
.A(n_20982),
.Y(n_21018)
);

NAND4xp25_ASAP7_75t_L g21019 ( 
.A(n_20978),
.B(n_20911),
.C(n_20952),
.D(n_20936),
.Y(n_21019)
);

INVx1_ASAP7_75t_L g21020 ( 
.A(n_20976),
.Y(n_21020)
);

BUFx2_ASAP7_75t_L g21021 ( 
.A(n_20977),
.Y(n_21021)
);

OAI22xp5_ASAP7_75t_SL g21022 ( 
.A1(n_20994),
.A2(n_21000),
.B1(n_21006),
.B2(n_21004),
.Y(n_21022)
);

INVx1_ASAP7_75t_L g21023 ( 
.A(n_20964),
.Y(n_21023)
);

AOI22xp5_ASAP7_75t_L g21024 ( 
.A1(n_20998),
.A2(n_21002),
.B1(n_21001),
.B2(n_21003),
.Y(n_21024)
);

INVx2_ASAP7_75t_L g21025 ( 
.A(n_20999),
.Y(n_21025)
);

CKINVDCx20_ASAP7_75t_R g21026 ( 
.A(n_20981),
.Y(n_21026)
);

OAI22xp5_ASAP7_75t_L g21027 ( 
.A1(n_20980),
.A2(n_20950),
.B1(n_20917),
.B2(n_20953),
.Y(n_21027)
);

NOR2xp33_ASAP7_75t_L g21028 ( 
.A(n_20986),
.B(n_20948),
.Y(n_21028)
);

OAI22xp5_ASAP7_75t_SL g21029 ( 
.A1(n_20995),
.A2(n_20942),
.B1(n_20945),
.B2(n_20917),
.Y(n_21029)
);

AOI221x1_ASAP7_75t_L g21030 ( 
.A1(n_20967),
.A2(n_20918),
.B1(n_5702),
.B2(n_5724),
.C(n_5661),
.Y(n_21030)
);

BUFx2_ASAP7_75t_L g21031 ( 
.A(n_20970),
.Y(n_21031)
);

HB1xp67_ASAP7_75t_L g21032 ( 
.A(n_20993),
.Y(n_21032)
);

INVx1_ASAP7_75t_L g21033 ( 
.A(n_20997),
.Y(n_21033)
);

INVxp67_ASAP7_75t_L g21034 ( 
.A(n_20991),
.Y(n_21034)
);

AOI21xp5_ASAP7_75t_L g21035 ( 
.A1(n_21005),
.A2(n_20992),
.B(n_20989),
.Y(n_21035)
);

AND4x1_ASAP7_75t_L g21036 ( 
.A(n_20979),
.B(n_5652),
.C(n_5495),
.D(n_5490),
.Y(n_21036)
);

AO21x2_ASAP7_75t_L g21037 ( 
.A1(n_20965),
.A2(n_8496),
.B(n_8748),
.Y(n_21037)
);

INVx2_ASAP7_75t_L g21038 ( 
.A(n_20988),
.Y(n_21038)
);

NAND3xp33_ASAP7_75t_L g21039 ( 
.A(n_21015),
.B(n_4614),
.C(n_4581),
.Y(n_21039)
);

AOI21xp5_ASAP7_75t_L g21040 ( 
.A1(n_21014),
.A2(n_7979),
.B(n_7975),
.Y(n_21040)
);

AND3x4_ASAP7_75t_L g21041 ( 
.A(n_21017),
.B(n_5773),
.C(n_5746),
.Y(n_21041)
);

AOI22xp5_ASAP7_75t_L g21042 ( 
.A1(n_21012),
.A2(n_8962),
.B1(n_6030),
.B2(n_6007),
.Y(n_21042)
);

XNOR2xp5_ASAP7_75t_L g21043 ( 
.A(n_21007),
.B(n_21010),
.Y(n_21043)
);

OAI221xp5_ASAP7_75t_L g21044 ( 
.A1(n_21011),
.A2(n_4618),
.B1(n_4614),
.B2(n_4581),
.C(n_5629),
.Y(n_21044)
);

NAND3xp33_ASAP7_75t_SL g21045 ( 
.A(n_21021),
.B(n_21008),
.C(n_21016),
.Y(n_21045)
);

OAI22xp5_ASAP7_75t_SL g21046 ( 
.A1(n_21018),
.A2(n_7616),
.B1(n_7890),
.B2(n_7606),
.Y(n_21046)
);

XNOR2xp5_ASAP7_75t_L g21047 ( 
.A(n_21022),
.B(n_5746),
.Y(n_21047)
);

INVx2_ASAP7_75t_SL g21048 ( 
.A(n_21020),
.Y(n_21048)
);

AOI22xp33_ASAP7_75t_L g21049 ( 
.A1(n_21023),
.A2(n_7388),
.B1(n_7396),
.B2(n_7387),
.Y(n_21049)
);

INVx4_ASAP7_75t_L g21050 ( 
.A(n_21025),
.Y(n_21050)
);

INVx1_ASAP7_75t_L g21051 ( 
.A(n_21024),
.Y(n_21051)
);

AOI22xp5_ASAP7_75t_L g21052 ( 
.A1(n_21026),
.A2(n_4614),
.B1(n_4618),
.B2(n_4581),
.Y(n_21052)
);

INVx1_ASAP7_75t_L g21053 ( 
.A(n_21032),
.Y(n_21053)
);

XNOR2x1_ASAP7_75t_L g21054 ( 
.A(n_21038),
.B(n_5773),
.Y(n_21054)
);

INVxp67_ASAP7_75t_SL g21055 ( 
.A(n_21034),
.Y(n_21055)
);

NAND2x1_ASAP7_75t_L g21056 ( 
.A(n_21031),
.B(n_21009),
.Y(n_21056)
);

AND2x2_ASAP7_75t_SL g21057 ( 
.A(n_21028),
.B(n_5629),
.Y(n_21057)
);

OA21x2_ASAP7_75t_L g21058 ( 
.A1(n_21019),
.A2(n_8496),
.B(n_8726),
.Y(n_21058)
);

INVx1_ASAP7_75t_L g21059 ( 
.A(n_21013),
.Y(n_21059)
);

INVx1_ASAP7_75t_L g21060 ( 
.A(n_21033),
.Y(n_21060)
);

XNOR2x1_ASAP7_75t_L g21061 ( 
.A(n_21027),
.B(n_5775),
.Y(n_21061)
);

XNOR2xp5_ASAP7_75t_L g21062 ( 
.A(n_21029),
.B(n_5775),
.Y(n_21062)
);

INVx1_ASAP7_75t_L g21063 ( 
.A(n_21035),
.Y(n_21063)
);

OR2x2_ASAP7_75t_L g21064 ( 
.A(n_21030),
.B(n_8206),
.Y(n_21064)
);

INVx2_ASAP7_75t_L g21065 ( 
.A(n_21050),
.Y(n_21065)
);

OR2x2_ASAP7_75t_SL g21066 ( 
.A(n_21045),
.B(n_21036),
.Y(n_21066)
);

NAND2xp5_ASAP7_75t_L g21067 ( 
.A(n_21043),
.B(n_21037),
.Y(n_21067)
);

INVx3_ASAP7_75t_SL g21068 ( 
.A(n_21048),
.Y(n_21068)
);

INVx2_ASAP7_75t_L g21069 ( 
.A(n_21051),
.Y(n_21069)
);

HB1xp67_ASAP7_75t_L g21070 ( 
.A(n_21060),
.Y(n_21070)
);

OAI21xp5_ASAP7_75t_L g21071 ( 
.A1(n_21059),
.A2(n_9464),
.B(n_9450),
.Y(n_21071)
);

XNOR2xp5_ASAP7_75t_L g21072 ( 
.A(n_21056),
.B(n_5775),
.Y(n_21072)
);

INVx1_ASAP7_75t_L g21073 ( 
.A(n_21055),
.Y(n_21073)
);

AND3x2_ASAP7_75t_L g21074 ( 
.A(n_21053),
.B(n_5775),
.C(n_5879),
.Y(n_21074)
);

OAI22xp5_ASAP7_75t_L g21075 ( 
.A1(n_21063),
.A2(n_8383),
.B1(n_8502),
.B2(n_8365),
.Y(n_21075)
);

XNOR2xp5_ASAP7_75t_L g21076 ( 
.A(n_21047),
.B(n_5879),
.Y(n_21076)
);

AND2x2_ASAP7_75t_L g21077 ( 
.A(n_21062),
.B(n_8202),
.Y(n_21077)
);

INVx4_ASAP7_75t_L g21078 ( 
.A(n_21057),
.Y(n_21078)
);

OAI22x1_ASAP7_75t_L g21079 ( 
.A1(n_21064),
.A2(n_7866),
.B1(n_7871),
.B2(n_7739),
.Y(n_21079)
);

OAI221xp5_ASAP7_75t_L g21080 ( 
.A1(n_21054),
.A2(n_4618),
.B1(n_4614),
.B2(n_5661),
.C(n_5629),
.Y(n_21080)
);

INVx1_ASAP7_75t_L g21081 ( 
.A(n_21061),
.Y(n_21081)
);

AOI22xp5_ASAP7_75t_L g21082 ( 
.A1(n_21041),
.A2(n_8502),
.B1(n_8383),
.B2(n_5629),
.Y(n_21082)
);

INVx1_ASAP7_75t_L g21083 ( 
.A(n_21070),
.Y(n_21083)
);

INVxp33_ASAP7_75t_SL g21084 ( 
.A(n_21073),
.Y(n_21084)
);

OAI221xp5_ASAP7_75t_L g21085 ( 
.A1(n_21068),
.A2(n_21039),
.B1(n_21040),
.B2(n_21052),
.C(n_21049),
.Y(n_21085)
);

OAI221xp5_ASAP7_75t_L g21086 ( 
.A1(n_21069),
.A2(n_21065),
.B1(n_21067),
.B2(n_21078),
.C(n_21081),
.Y(n_21086)
);

AOI322xp5_ASAP7_75t_L g21087 ( 
.A1(n_21066),
.A2(n_21042),
.A3(n_21044),
.B1(n_21058),
.B2(n_21046),
.C1(n_7645),
.C2(n_7632),
.Y(n_21087)
);

OR2x2_ASAP7_75t_L g21088 ( 
.A(n_21072),
.B(n_5629),
.Y(n_21088)
);

OR2x2_ASAP7_75t_L g21089 ( 
.A(n_21076),
.B(n_5661),
.Y(n_21089)
);

XNOR2xp5_ASAP7_75t_L g21090 ( 
.A(n_21077),
.B(n_5879),
.Y(n_21090)
);

NAND5xp2_ASAP7_75t_L g21091 ( 
.A(n_21080),
.B(n_5495),
.C(n_5490),
.D(n_6033),
.E(n_6893),
.Y(n_21091)
);

INVx1_ASAP7_75t_L g21092 ( 
.A(n_21079),
.Y(n_21092)
);

XOR2xp5_ASAP7_75t_L g21093 ( 
.A(n_21082),
.B(n_4618),
.Y(n_21093)
);

INVx1_ASAP7_75t_L g21094 ( 
.A(n_21083),
.Y(n_21094)
);

INVx1_ASAP7_75t_L g21095 ( 
.A(n_21084),
.Y(n_21095)
);

OAI21xp5_ASAP7_75t_L g21096 ( 
.A1(n_21086),
.A2(n_21071),
.B(n_21075),
.Y(n_21096)
);

OAI21xp5_ASAP7_75t_L g21097 ( 
.A1(n_21092),
.A2(n_21074),
.B(n_9464),
.Y(n_21097)
);

OAI21x1_ASAP7_75t_L g21098 ( 
.A1(n_21089),
.A2(n_9464),
.B(n_9450),
.Y(n_21098)
);

AO21x1_ASAP7_75t_L g21099 ( 
.A1(n_21088),
.A2(n_7801),
.B(n_7766),
.Y(n_21099)
);

OR2x2_ASAP7_75t_L g21100 ( 
.A(n_21085),
.B(n_5661),
.Y(n_21100)
);

AOI21xp33_ASAP7_75t_SL g21101 ( 
.A1(n_21090),
.A2(n_8726),
.B(n_9047),
.Y(n_21101)
);

AOI22x1_ASAP7_75t_L g21102 ( 
.A1(n_21093),
.A2(n_4618),
.B1(n_5702),
.B2(n_5661),
.Y(n_21102)
);

OAI21xp5_ASAP7_75t_L g21103 ( 
.A1(n_21087),
.A2(n_9468),
.B(n_9450),
.Y(n_21103)
);

INVx1_ASAP7_75t_L g21104 ( 
.A(n_21094),
.Y(n_21104)
);

AOI22xp5_ASAP7_75t_L g21105 ( 
.A1(n_21095),
.A2(n_21091),
.B1(n_4618),
.B2(n_8502),
.Y(n_21105)
);

AOI22xp33_ASAP7_75t_L g21106 ( 
.A1(n_21096),
.A2(n_8502),
.B1(n_8383),
.B2(n_7388),
.Y(n_21106)
);

NAND3xp33_ASAP7_75t_L g21107 ( 
.A(n_21100),
.B(n_5702),
.C(n_5661),
.Y(n_21107)
);

AOI21xp33_ASAP7_75t_SL g21108 ( 
.A1(n_21097),
.A2(n_21102),
.B(n_21103),
.Y(n_21108)
);

NAND2xp5_ASAP7_75t_L g21109 ( 
.A(n_21099),
.B(n_5661),
.Y(n_21109)
);

OAI21xp5_ASAP7_75t_SL g21110 ( 
.A1(n_21101),
.A2(n_21098),
.B(n_5724),
.Y(n_21110)
);

AOI22xp5_ASAP7_75t_L g21111 ( 
.A1(n_21094),
.A2(n_8502),
.B1(n_8383),
.B2(n_7616),
.Y(n_21111)
);

AOI21xp5_ASAP7_75t_L g21112 ( 
.A1(n_21104),
.A2(n_7979),
.B(n_7975),
.Y(n_21112)
);

NAND2xp5_ASAP7_75t_L g21113 ( 
.A(n_21108),
.B(n_5702),
.Y(n_21113)
);

AOI22xp5_ASAP7_75t_L g21114 ( 
.A1(n_21110),
.A2(n_8502),
.B1(n_8383),
.B2(n_7616),
.Y(n_21114)
);

AOI22xp33_ASAP7_75t_L g21115 ( 
.A1(n_21107),
.A2(n_8502),
.B1(n_8383),
.B2(n_7388),
.Y(n_21115)
);

NAND2xp5_ASAP7_75t_L g21116 ( 
.A(n_21109),
.B(n_5702),
.Y(n_21116)
);

NAND2xp5_ASAP7_75t_L g21117 ( 
.A(n_21105),
.B(n_5702),
.Y(n_21117)
);

OAI21xp5_ASAP7_75t_L g21118 ( 
.A1(n_21106),
.A2(n_8693),
.B(n_8615),
.Y(n_21118)
);

AOI21xp5_ASAP7_75t_L g21119 ( 
.A1(n_21111),
.A2(n_7979),
.B(n_7975),
.Y(n_21119)
);

NAND2xp5_ASAP7_75t_SL g21120 ( 
.A(n_21117),
.B(n_7976),
.Y(n_21120)
);

OAI21xp5_ASAP7_75t_SL g21121 ( 
.A1(n_21113),
.A2(n_7631),
.B(n_5879),
.Y(n_21121)
);

INVx1_ASAP7_75t_L g21122 ( 
.A(n_21116),
.Y(n_21122)
);

OR2x6_ASAP7_75t_L g21123 ( 
.A(n_21122),
.B(n_21119),
.Y(n_21123)
);

INVxp67_ASAP7_75t_SL g21124 ( 
.A(n_21120),
.Y(n_21124)
);

NAND2xp5_ASAP7_75t_L g21125 ( 
.A(n_21121),
.B(n_21115),
.Y(n_21125)
);

NAND2xp5_ASAP7_75t_L g21126 ( 
.A(n_21124),
.B(n_21114),
.Y(n_21126)
);

OAI221xp5_ASAP7_75t_R g21127 ( 
.A1(n_21126),
.A2(n_21123),
.B1(n_21125),
.B2(n_21112),
.C(n_21118),
.Y(n_21127)
);

AOI22xp5_ASAP7_75t_SL g21128 ( 
.A1(n_21127),
.A2(n_5702),
.B1(n_5724),
.B2(n_5879),
.Y(n_21128)
);

AOI211xp5_ASAP7_75t_L g21129 ( 
.A1(n_21128),
.A2(n_5702),
.B(n_5724),
.C(n_5431),
.Y(n_21129)
);


endmodule