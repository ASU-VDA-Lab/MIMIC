module fake_jpeg_22764_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_28),
.B1(n_30),
.B2(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_26),
.B1(n_35),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_53),
.B1(n_62),
.B2(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_7),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_22),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_39),
.B1(n_32),
.B2(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_61),
.B1(n_55),
.B2(n_65),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_81),
.B1(n_28),
.B2(n_21),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_28),
.B1(n_47),
.B2(n_27),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_39),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_41),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_38),
.B1(n_20),
.B2(n_19),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_32),
.C(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_87),
.C(n_17),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_43),
.B1(n_22),
.B2(n_23),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_42),
.A2(n_40),
.B(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_38),
.B1(n_28),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_47),
.B1(n_49),
.B2(n_41),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_64),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_103),
.C(n_106),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_88),
.A3(n_72),
.B1(n_78),
.B2(n_66),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_110),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_60),
.B1(n_53),
.B2(n_51),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_60),
.Y(n_106)
);

NOR2x1p5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_43),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_43),
.B1(n_22),
.B2(n_23),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_24),
.B(n_15),
.C(n_16),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_27),
.B1(n_15),
.B2(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_87),
.B(n_82),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_135),
.B(n_137),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_66),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_69),
.B1(n_74),
.B2(n_73),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_133),
.B1(n_139),
.B2(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_72),
.C(n_78),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_24),
.C(n_98),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_115),
.B(n_60),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_75),
.B(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_83),
.B(n_17),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_69),
.B1(n_27),
.B2(n_15),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_54),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_91),
.B1(n_103),
.B2(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_148),
.B1(n_153),
.B2(n_127),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_108),
.B(n_54),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_132),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_150),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_111),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_152),
.C(n_165),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_109),
.B1(n_96),
.B2(n_23),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_130),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_25),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_164),
.Y(n_168)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_25),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_175),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_124),
.A3(n_122),
.B1(n_132),
.B2(n_121),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_185),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_131),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_187),
.C(n_31),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_184),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_147),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_25),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_132),
.A3(n_133),
.B1(n_127),
.B2(n_120),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_120),
.B1(n_137),
.B2(n_126),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_147),
.B1(n_158),
.B2(n_143),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_131),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_125),
.B1(n_119),
.B2(n_118),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_139),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_161),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_166),
.B1(n_173),
.B2(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_159),
.B1(n_148),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_200),
.B1(n_212),
.B2(n_168),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_109),
.B1(n_84),
.B2(n_23),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_10),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_8),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_172),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_109),
.B1(n_84),
.B2(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_207),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_84),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_170),
.B(n_171),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_31),
.B1(n_18),
.B2(n_25),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_31),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_167),
.B1(n_181),
.B2(n_185),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_173),
.C(n_174),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_231),
.C(n_208),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_230),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_223),
.B1(n_208),
.B2(n_205),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_192),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_31),
.B(n_18),
.C(n_7),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_197),
.B1(n_196),
.B2(n_191),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_18),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_18),
.C(n_1),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_204),
.B1(n_203),
.B2(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_218),
.B1(n_224),
.B2(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_199),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_216),
.C(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_14),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_208),
.B1(n_198),
.B2(n_194),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_202),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_202),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_210),
.B1(n_195),
.B2(n_2),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_6),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_14),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_7),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_260),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_263),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_262),
.C(n_0),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_229),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_259),
.B(n_238),
.Y(n_264)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_14),
.B(n_13),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_0),
.C(n_1),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_239),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_273),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_242),
.B(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_275),
.C(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_272),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_235),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_261),
.B1(n_12),
.B2(n_9),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_253),
.B1(n_262),
.B2(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_4),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_0),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_275),
.B(n_269),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_4),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_1),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_290),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_271),
.B(n_265),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_289),
.B(n_291),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_2),
.B(n_4),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_281),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_296),
.B(n_277),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.C(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_277),
.C(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_4),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_5),
.Y(n_303)
);


endmodule