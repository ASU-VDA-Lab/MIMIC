module real_jpeg_11260_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_17),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_9),
.B1(n_17),
.B2(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_18),
.B1(n_19),
.B2(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_8),
.B(n_18),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_5),
.A2(n_25),
.B(n_64),
.C(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_25),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_5),
.A2(n_8),
.B(n_45),
.Y(n_112)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_19),
.B(n_22),
.C(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_9),
.B1(n_32),
.B2(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_33),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_9),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_39),
.B(n_40),
.C(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_9),
.B(n_40),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_32),
.B(n_40),
.C(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_100),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_98),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_69),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_13),
.B(n_69),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_55),
.C(n_62),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_14),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_37),
.C(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_30),
.B2(n_33),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_16),
.A2(n_33),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_31),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_25),
.A2(n_29),
.B(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_26),
.A2(n_32),
.B(n_66),
.C(n_112),
.Y(n_111)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_32),
.B(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_32),
.B(n_65),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_53),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_38),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_41),
.B(n_105),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B(n_49),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_44),
.B(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_53),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_129),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_59),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_62),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_62),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_94),
.C(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_68),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_88),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_76),
.A2(n_77),
.B1(n_106),
.B2(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_106),
.C(n_137),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_94),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_119),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_139),
.B(n_143),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_131),
.B(n_138),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_122),
.B(n_130),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_114),
.B(n_121),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_111),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B(n_120),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_133),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_141),
.Y(n_143)
);


endmodule