module fake_jpeg_17469_n_179 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_36),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_16),
.B1(n_27),
.B2(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_43),
.B1(n_24),
.B2(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_16),
.B1(n_13),
.B2(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_13),
.B1(n_25),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_48),
.B1(n_21),
.B2(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_36),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_3),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_30),
.C(n_26),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_69),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_26),
.B1(n_36),
.B2(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_11),
.B(n_2),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_33),
.B(n_36),
.C(n_17),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_47),
.B(n_44),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_19),
.C(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_17),
.B1(n_1),
.B2(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_68),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_33),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_47),
.C(n_39),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_49),
.B(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_68),
.B1(n_84),
.B2(n_87),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_65),
.B(n_55),
.C(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_97),
.B1(n_108),
.B2(n_74),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_109),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_106),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_102),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_50),
.B1(n_59),
.B2(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_70),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_59),
.C(n_66),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_75),
.B1(n_88),
.B2(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_117),
.C(n_93),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_85),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_80),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_121),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_93),
.B1(n_106),
.B2(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_77),
.C(n_95),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_72),
.C(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_120),
.A3(n_125),
.B1(n_123),
.B2(n_121),
.C(n_73),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_137),
.A3(n_94),
.B1(n_71),
.B2(n_113),
.C(n_110),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_73),
.B(n_94),
.C(n_119),
.D(n_122),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_71),
.C(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_74),
.B1(n_113),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_150),
.B1(n_139),
.B2(n_140),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_94),
.B(n_56),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_94),
.B(n_58),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_17),
.B(n_1),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_133),
.B1(n_132),
.B2(n_135),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_146),
.C(n_150),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_158),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_130),
.B1(n_138),
.B2(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_147),
.B1(n_142),
.B2(n_10),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_58),
.B1(n_46),
.B2(n_5),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_157),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_9),
.B1(n_4),
.B2(n_6),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_7),
.B(n_9),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_142),
.C(n_154),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_12),
.B(n_29),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_12),
.Y(n_172)
);

NAND4xp25_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_7),
.C(n_9),
.D(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_168),
.C(n_170),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_162),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_174),
.B(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_29),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_29),
.Y(n_179)
);


endmodule