module fake_jpeg_32093_n_52 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_17;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

AND2x6_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_11),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_1),
.B(n_3),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_17),
.B(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_14),
.B1(n_20),
.B2(n_24),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_32),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_30),
.B1(n_16),
.B2(n_20),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_41),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx24_ASAP7_75t_SL g43 ( 
.A(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_42),
.B1(n_14),
.B2(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_25),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_48),
.C2(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.Y(n_52)
);


endmodule