module fake_jpeg_31809_n_445 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_445);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_18),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_12),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_12),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_66),
.B(n_74),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_34),
.B1(n_45),
.B2(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_39),
.B1(n_27),
.B2(n_36),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_125),
.Y(n_144)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_86),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_129),
.Y(n_166)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_140),
.Y(n_200)
);

CKINVDCx12_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_146),
.B(n_157),
.Y(n_189)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_114),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_171),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_175),
.B1(n_39),
.B2(n_27),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_88),
.B1(n_55),
.B2(n_67),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_29),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_31),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_166),
.Y(n_194)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_167),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_44),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_94),
.B(n_26),
.C(n_72),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_106),
.C(n_27),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_37),
.B1(n_30),
.B2(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_39),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_176),
.Y(n_204)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_174),
.Y(n_201)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_123),
.A2(n_82),
.B1(n_79),
.B2(n_84),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_134),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_100),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_176),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_156),
.B1(n_28),
.B2(n_112),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_109),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_150),
.C(n_36),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_150),
.B(n_28),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_164),
.Y(n_217)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_81),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_226),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_151),
.B(n_161),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_204),
.B1(n_187),
.B2(n_184),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_213),
.B1(n_224),
.B2(n_227),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_216),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_153),
.B1(n_168),
.B2(n_162),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_225),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_186),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_143),
.C(n_141),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_159),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_186),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_158),
.B(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_183),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_110),
.B1(n_118),
.B2(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_192),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_202),
.B1(n_189),
.B2(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_243),
.B1(n_227),
.B2(n_216),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_252),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_189),
.B1(n_119),
.B2(n_131),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_246),
.B1(n_221),
.B2(n_207),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_115),
.B1(n_136),
.B2(n_118),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_192),
.B1(n_200),
.B2(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_210),
.B(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_197),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_226),
.C(n_197),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_253),
.B1(n_247),
.B2(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_208),
.B(n_207),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_278),
.B(n_235),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_263),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_212),
.C(n_220),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_269),
.C(n_281),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_272),
.B1(n_274),
.B2(n_239),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_254),
.A2(n_216),
.B(n_206),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_283),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_222),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_275),
.B(n_20),
.C(n_76),
.D(n_49),
.Y(n_311)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_271),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_218),
.B1(n_200),
.B2(n_205),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_180),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_218),
.B1(n_200),
.B2(n_177),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_234),
.B(n_180),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_199),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_279),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_191),
.B(n_95),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_179),
.C(n_199),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_179),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_95),
.B1(n_45),
.B2(n_127),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_284),
.A2(n_288),
.B1(n_290),
.B2(n_295),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_286),
.A2(n_287),
.B1(n_297),
.B2(n_283),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_231),
.B1(n_246),
.B2(n_251),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_270),
.B1(n_261),
.B2(n_264),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_231),
.B1(n_253),
.B2(n_243),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_236),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_301),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_236),
.B1(n_245),
.B2(n_177),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_174),
.B1(n_173),
.B2(n_148),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_300),
.A2(n_267),
.B(n_276),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_122),
.B(n_127),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_195),
.C(n_121),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_274),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_195),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_259),
.A2(n_147),
.B1(n_175),
.B2(n_140),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_136),
.B1(n_110),
.B2(n_92),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_139),
.C(n_105),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.C(n_289),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_89),
.C(n_87),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_73),
.C(n_99),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_286),
.B1(n_299),
.B2(n_297),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_276),
.C(n_267),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_335),
.C(n_328),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_324),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_325),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_266),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_273),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_334),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_277),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_329),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_282),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_337),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_336),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_272),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_280),
.C(n_257),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_256),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_338),
.A2(n_290),
.B1(n_292),
.B2(n_295),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_356),
.B1(n_14),
.B2(n_1),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_300),
.B1(n_296),
.B2(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_307),
.B1(n_287),
.B2(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_348),
.Y(n_363)
);

FAx1_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_310),
.CI(n_303),
.CON(n_346),
.SN(n_346)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_355),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_320),
.A2(n_315),
.B(n_337),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_306),
.B1(n_309),
.B2(n_285),
.Y(n_352)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_16),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_83),
.B1(n_80),
.B2(n_78),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_331),
.A2(n_15),
.B(n_17),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_16),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_361),
.C(n_324),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_375),
.C(n_339),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_330),
.B1(n_335),
.B2(n_314),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_367),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_336),
.B1(n_321),
.B2(n_34),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_371),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_14),
.C(n_17),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_369),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_13),
.Y(n_371)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_380),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_34),
.B1(n_69),
.B2(n_99),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_380),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_353),
.A2(n_16),
.B(n_14),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_374),
.A2(n_370),
.B(n_377),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_34),
.C(n_51),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_355),
.B1(n_350),
.B2(n_360),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_0),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_384),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_347),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_388),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_347),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_390),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_378),
.B(n_370),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_361),
.C(n_339),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_396),
.C(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_346),
.C(n_342),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_399),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_394),
.A2(n_381),
.B1(n_364),
.B2(n_376),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_396),
.A2(n_344),
.B1(n_372),
.B2(n_341),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_404),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_375),
.B(n_341),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_403),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_362),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_385),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_408),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_358),
.B(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_393),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_401),
.A2(n_383),
.B(n_388),
.C(n_387),
.Y(n_411)
);

OAI21x1_ASAP7_75t_SL g422 ( 
.A1(n_411),
.A2(n_414),
.B(n_419),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_382),
.C(n_383),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_416),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_407),
.A2(n_406),
.B(n_398),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_393),
.C(n_356),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_420),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_399),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_410),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_424),
.Y(n_431)
);

BUFx24_ASAP7_75t_SL g424 ( 
.A(n_415),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_412),
.B(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_426),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_411),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_427),
.A2(n_3),
.B(n_4),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_24),
.C(n_1),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_428),
.B(n_0),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_2),
.B(n_3),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_423),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_429),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_3),
.B(n_4),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_436),
.A2(n_438),
.B(n_430),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_5),
.C(n_6),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_24),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_441),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_442),
.B(n_439),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_5),
.C(n_24),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_5),
.B(n_24),
.Y(n_445)
);


endmodule