module fake_jpeg_29939_n_414 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_414);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_71),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_76),
.Y(n_93)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_14),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_74),
.Y(n_117)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_81),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_1),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_85),
.Y(n_124)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_45),
.B(n_1),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_116),
.C(n_47),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_70),
.B1(n_32),
.B2(n_28),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_95),
.A2(n_107),
.B1(n_111),
.B2(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_17),
.B1(n_41),
.B2(n_37),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_20),
.B(n_18),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_84),
.B1(n_60),
.B2(n_61),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_31),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_51),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_119),
.B(n_35),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_25),
.B1(n_29),
.B2(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_29),
.B1(n_25),
.B2(n_36),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_46),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_50),
.B1(n_64),
.B2(n_48),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_134),
.A2(n_152),
.B1(n_103),
.B2(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_145),
.B1(n_103),
.B2(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_68),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_23),
.Y(n_140)
);

OR2x2_ASAP7_75t_SL g141 ( 
.A(n_93),
.B(n_67),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_149),
.Y(n_182)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_144),
.B(n_159),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_78),
.B1(n_63),
.B2(n_59),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_16),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_158),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_65),
.B1(n_56),
.B2(n_18),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_133),
.B1(n_102),
.B2(n_114),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_58),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g155 ( 
.A(n_100),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_101),
.Y(n_157)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_36),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_83),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_13),
.B(n_24),
.C(n_5),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_165),
.Y(n_200)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_35),
.B(n_14),
.Y(n_167)
);

OAI21x1_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_176),
.B(n_35),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_91),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_173),
.Y(n_208)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_49),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_98),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_127),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_127),
.Y(n_179)
);

AND2x4_ASAP7_75t_SL g176 ( 
.A(n_115),
.B(n_49),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_185),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_203),
.B1(n_172),
.B2(n_161),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_115),
.C(n_121),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_188),
.C(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_213),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_106),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_138),
.B(n_106),
.C(n_97),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_189),
.B(n_150),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_121),
.C(n_87),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_97),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_123),
.B1(n_108),
.B2(n_118),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_87),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_167),
.B(n_135),
.Y(n_230)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_140),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_218),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_149),
.B1(n_162),
.B2(n_153),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_238),
.B1(n_243),
.B2(n_248),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_182),
.B1(n_180),
.B2(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_142),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_139),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_198),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_230),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_178),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_159),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_241),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_209),
.B1(n_186),
.B2(n_191),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_153),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_202),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_163),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_153),
.B(n_168),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_245),
.B(n_199),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_171),
.B1(n_98),
.B2(n_108),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_246),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_182),
.B(n_189),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_169),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_157),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_183),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_184),
.A2(n_155),
.B1(n_123),
.B2(n_176),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_253),
.B1(n_260),
.B2(n_248),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_261),
.C(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_202),
.B1(n_199),
.B2(n_176),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_254),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_230),
.B1(n_222),
.B2(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_265),
.B1(n_267),
.B2(n_241),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_258),
.B(n_247),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_219),
.A2(n_224),
.B1(n_232),
.B2(n_239),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_218),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_231),
.B(n_227),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_242),
.B1(n_238),
.B2(n_226),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_156),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_151),
.B1(n_211),
.B2(n_204),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_148),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_275),
.C(n_193),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_236),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_223),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_146),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_160),
.B1(n_196),
.B2(n_204),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_278),
.A2(n_192),
.B(n_160),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_279),
.A2(n_291),
.B1(n_293),
.B2(n_275),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_280),
.A2(n_285),
.B1(n_292),
.B2(n_266),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_281),
.B(n_303),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_245),
.B(n_222),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_245),
.B1(n_231),
.B2(n_240),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_249),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_295),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_233),
.B1(n_229),
.B2(n_211),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_220),
.B1(n_228),
.B2(n_212),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_253),
.A2(n_228),
.B1(n_207),
.B2(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_183),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_207),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_300),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_157),
.B(n_143),
.C(n_160),
.D(n_192),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_272),
.B(n_198),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_274),
.B(n_170),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_263),
.B1(n_276),
.B2(n_254),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_305),
.A2(n_24),
.B1(n_3),
.B2(n_5),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_286),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_252),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_314),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_312),
.A2(n_292),
.B1(n_326),
.B2(n_324),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_257),
.B1(n_270),
.B2(n_264),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_324),
.B1(n_325),
.B2(n_328),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_260),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g315 ( 
.A(n_285),
.B(n_257),
.C(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_300),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_258),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_320),
.C(n_295),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_268),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_261),
.B1(n_24),
.B2(n_6),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_302),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_280),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_338),
.C(n_346),
.Y(n_357)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_310),
.C(n_319),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_311),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_323),
.B(n_297),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_342),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_311),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_312),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_321),
.B(n_294),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_327),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_284),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_345),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_293),
.C(n_284),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_291),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_329),
.C(n_318),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_329),
.C(n_322),
.Y(n_359)
);

FAx1_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_308),
.CI(n_307),
.CON(n_350),
.SN(n_350)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_356),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_332),
.B1(n_336),
.B2(n_348),
.Y(n_366)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_308),
.B(n_315),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_358),
.A2(n_365),
.B(n_325),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_337),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_363),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_332),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_341),
.A2(n_298),
.B(n_305),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_366),
.B(n_372),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_355),
.B(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_369),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_370),
.C(n_375),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_346),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_337),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_358),
.B(n_349),
.CI(n_338),
.CON(n_371),
.SN(n_371)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_374),
.B(n_376),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_347),
.C(n_336),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_298),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_353),
.A2(n_328),
.B1(n_299),
.B2(n_8),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_365),
.C(n_353),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_381),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_351),
.C(n_350),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_364),
.B1(n_361),
.B2(n_356),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_383),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_352),
.B1(n_354),
.B2(n_350),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_352),
.C(n_354),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_389),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_6),
.C(n_7),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_371),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_390),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_375),
.C(n_371),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_395),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_386),
.A2(n_377),
.B(n_378),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_397),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_8),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_393),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_9),
.C(n_10),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_388),
.B(n_11),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_10),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_399),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_396),
.B(n_10),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_404),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_401),
.A2(n_394),
.B(n_398),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_406),
.A2(n_407),
.B(n_393),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_402),
.A2(n_399),
.B(n_395),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_409),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_405),
.A2(n_403),
.B(n_400),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_411),
.A2(n_410),
.B(n_408),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_412),
.B(n_11),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_11),
.C(n_12),
.Y(n_414)
);


endmodule