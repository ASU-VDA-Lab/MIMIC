module real_jpeg_26145_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_346, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_346;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_1),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_67),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_47),
.C(n_50),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_130),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_1),
.B(n_30),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_1),
.A2(n_104),
.B1(n_209),
.B2(n_213),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_42),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_4),
.A2(n_26),
.B1(n_58),
.B2(n_65),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_7),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_127),
.Y(n_273)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_9),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_134),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_134),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_69),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_14),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_125),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_125),
.Y(n_202)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_20),
.A2(n_73),
.B1(n_329),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_20),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_44),
.C(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_24),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_25),
.A2(n_30),
.B(n_38),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_25),
.A2(n_38),
.B(n_81),
.Y(n_274)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_27),
.A2(n_62),
.B(n_131),
.C(n_153),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g225 ( 
.A(n_27),
.B(n_130),
.CON(n_225),
.SN(n_225)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_29),
.B(n_63),
.C(n_66),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g226 ( 
.A(n_29),
.B(n_32),
.C(n_34),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_30),
.A2(n_38),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_30),
.A2(n_38),
.B1(n_169),
.B2(n_225),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_30),
.A2(n_38),
.B1(n_80),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_31),
.A2(n_144),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_31),
.A2(n_37),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_33),
.A2(n_36),
.B(n_224),
.C(n_226),
.Y(n_223)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_34),
.B(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_38),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_38),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_73),
.C(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_43),
.A2(n_44),
.B1(n_79),
.B2(n_332),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_45),
.A2(n_49),
.B1(n_184),
.B2(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_45),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_45),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_49),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_49),
.B(n_130),
.Y(n_207)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_51),
.B(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_117),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_53),
.B(n_182),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_61),
.B(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_68),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_67),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_60),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_60),
.A2(n_67),
.B1(n_141),
.B2(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_61),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_67),
.B(n_294),
.Y(n_293)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_73),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_73),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_76),
.B(n_130),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_78),
.B(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_79),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_88),
.A2(n_139),
.B(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_326),
.A3(n_338),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_303),
.B(n_325),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_277),
.B(n_302),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_171),
.B(n_258),
.C(n_276),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_155),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_100),
.B(n_155),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_135),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_120),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_102),
.B(n_120),
.C(n_135),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_103),
.B(n_114),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B(n_110),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_104),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_104),
.A2(n_202),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_104),
.A2(n_110),
.B(n_191),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_104),
.A2(n_191),
.B(n_213),
.Y(n_283)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_109),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_105),
.B(n_111),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_105),
.A2(n_163),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_107),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_113),
.B(n_130),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_116),
.B(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_117),
.A2(n_182),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_117),
.A2(n_182),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_128),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_123),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_122),
.Y(n_286)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_145),
.B2(n_154),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_138),
.B(n_142),
.C(n_154),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_139),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_156),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_160),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_164),
.B(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_257),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_252),
.B(n_256),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_236),
.B(n_251),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_219),
.B(n_235),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_198),
.B(n_218),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_180),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_193),
.C(n_196),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_205),
.B(n_217),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_204),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_216),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_234),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_234),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_230),
.C(n_231),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_246),
.C(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_260),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_269),
.C(n_275),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_268),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_268),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_272),
.C(n_274),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_273),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_279),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_301),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_288),
.B1(n_299),
.B2(n_300),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_300),
.C(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_287),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_283),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_313),
.B(n_317),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_295),
.C(n_298),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_304),
.B(n_305),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_312),
.B1(n_320),
.B2(n_321),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_310),
.B(n_311),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_328),
.B1(n_333),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_320),
.C(n_324),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_335),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_335),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.C(n_334),
.Y(n_327)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_339),
.B(n_340),
.Y(n_343)
);


endmodule