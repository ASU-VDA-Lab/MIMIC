module real_jpeg_28153_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_313, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_313;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_46),
.Y(n_94)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_0),
.Y(n_256)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_5),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_159),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_159),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_159),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_6),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_6),
.A2(n_29),
.B(n_66),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_68),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_6),
.A2(n_35),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_35),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_77),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_93),
.B1(n_252),
.B2(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_6),
.A2(n_28),
.B(n_268),
.Y(n_267)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_42),
.B1(n_60),
.B2(n_61),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_8),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_9),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_136),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_9),
.A2(n_46),
.B1(n_48),
.B2(n_136),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_136),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_11),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_103),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_103),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_11),
.A2(n_46),
.B1(n_48),
.B2(n_103),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_12),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_152),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_152),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_152),
.Y(n_246)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_15),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_55),
.Y(n_112)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_63),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_17),
.A2(n_46),
.B1(n_48),
.B2(n_63),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_22),
.B(n_119),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_56),
.CI(n_82),
.CON(n_22),
.SN(n_22)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_23),
.A2(n_24),
.B(n_43),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_38),
.B2(n_41),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_25),
.A2(n_32),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_25),
.A2(n_32),
.B1(n_168),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_25),
.A2(n_32),
.B1(n_201),
.B2(n_267),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_31),
.C(n_32),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_28),
.A2(n_33),
.A3(n_36),
.B1(n_269),
.B2(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_29),
.B(n_163),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_33),
.Y(n_278)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_36),
.B1(n_49),
.B2(n_51),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_35),
.A2(n_48),
.A3(n_51),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_35),
.B(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_39),
.A2(n_75),
.B1(n_77),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_54),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_45),
.B(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_44),
.A2(n_45),
.B1(n_88),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_44),
.A2(n_45),
.B1(n_133),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_44),
.A2(n_45),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_44),
.A2(n_45),
.B1(n_226),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_44),
.A2(n_45),
.B1(n_193),
.B2(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_45),
.B(n_163),
.Y(n_253)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_46),
.B(n_49),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_46),
.B(n_258),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_72),
.B2(n_81),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_58),
.B1(n_106),
.B2(n_114),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_73),
.C(n_80),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_64),
.B1(n_71),
.B2(n_101),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_61),
.A2(n_69),
.B(n_163),
.C(n_164),
.Y(n_162)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_64),
.A2(n_71),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_68),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_65),
.A2(n_68),
.B1(n_102),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_65),
.A2(n_68),
.B1(n_135),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_65),
.A2(n_68),
.B1(n_158),
.B2(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_75),
.A2(n_77),
.B1(n_128),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_75),
.A2(n_77),
.B1(n_189),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_80),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_99),
.B(n_100),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_84),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_85),
.A2(n_86),
.B1(n_92),
.B2(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_89),
.A2(n_91),
.B1(n_148),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_89),
.A2(n_91),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_99),
.B1(n_100),
.B2(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_98),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_95),
.B1(n_131),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_93),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_93),
.A2(n_97),
.B1(n_246),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_93),
.A2(n_240),
.B1(n_241),
.B2(n_280),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_96),
.B1(n_145),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_94),
.A2(n_96),
.B1(n_166),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_94),
.A2(n_96),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_SL g241 ( 
.A(n_96),
.Y(n_241)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_97),
.B(n_163),
.Y(n_258)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_137),
.B(n_310),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_125),
.A2(n_126),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_134),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_127),
.B(n_129),
.CI(n_134),
.CON(n_174),
.SN(n_174)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_132),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_176),
.A3(n_181),
.B1(n_304),
.B2(n_309),
.C(n_313),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_139),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_171),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_140),
.B(n_171),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.C(n_170),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_141),
.B(n_170),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_150),
.C(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_146),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_155),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.C(n_167),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_167),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_161),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_165),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_174),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_177),
.B(n_178),
.Y(n_309)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_211),
.C(n_216),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_205),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_183),
.B(n_205),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_196),
.C(n_197),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_184),
.B(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_194),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_191),
.C(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_196),
.Y(n_302)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_202),
.B(n_204),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_203),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_212),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_213),
.B(n_214),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_298),
.B(n_303),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_284),
.B(n_297),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_262),
.B(n_283),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_242),
.B(n_261),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_221),
.B(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_249),
.B(n_260),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_248),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_254),
.B(n_259),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_275),
.B1(n_281),
.B2(n_282),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_274),
.C(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_275),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_293),
.C(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);


endmodule