module real_aes_7699_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g504 ( .A1(n_0), .A2(n_168), .B(n_505), .C(n_508), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_1), .B(n_500), .Y(n_509) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_88), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g166 ( .A(n_3), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_4), .B(n_169), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_468), .B(n_544), .Y(n_543) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_6), .A2(n_176), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_7), .A2(n_35), .B1(n_156), .B2(n_204), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_8), .B(n_176), .Y(n_184) );
AND2x6_ASAP7_75t_L g171 ( .A(n_9), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_10), .A2(n_171), .B(n_473), .C(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_11), .B(n_36), .Y(n_124) );
INVx1_ASAP7_75t_L g150 ( .A(n_12), .Y(n_150) );
INVx1_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_14), .B(n_152), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_15), .B(n_169), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_16), .B(n_143), .Y(n_250) );
AO32x2_ASAP7_75t_L g220 ( .A1(n_17), .A2(n_142), .A3(n_176), .B1(n_195), .B2(n_221), .Y(n_220) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_18), .A2(n_39), .B1(n_127), .B2(n_746), .C1(n_747), .C2(n_749), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_19), .B(n_156), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_20), .B(n_143), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_21), .A2(n_53), .B1(n_156), .B2(n_204), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_22), .A2(n_80), .B1(n_152), .B2(n_156), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_23), .B(n_156), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_24), .A2(n_195), .B(n_473), .C(n_491), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_25), .A2(n_195), .B(n_473), .C(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_26), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_27), .B(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_28), .A2(n_468), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_29), .B(n_197), .Y(n_238) );
INVx2_ASAP7_75t_L g154 ( .A(n_30), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_31), .A2(n_471), .B(n_475), .C(n_481), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_32), .B(n_156), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_33), .B(n_197), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_34), .B(n_215), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_36), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_37), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_38), .Y(n_521) );
INVx1_ASAP7_75t_L g746 ( .A(n_39), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_40), .B(n_169), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_41), .B(n_468), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_42), .A2(n_130), .B1(n_131), .B2(n_452), .Y(n_129) );
INVx1_ASAP7_75t_L g452 ( .A(n_42), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_42), .A2(n_44), .B1(n_452), .B2(n_758), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_43), .A2(n_471), .B(n_481), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_44), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_45), .B(n_156), .Y(n_179) );
INVx1_ASAP7_75t_L g506 ( .A(n_46), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_47), .A2(n_89), .B1(n_204), .B2(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g537 ( .A(n_48), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_49), .B(n_156), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_50), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_51), .B(n_468), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_52), .B(n_164), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_54), .A2(n_58), .B1(n_152), .B2(n_156), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_55), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_56), .B(n_156), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_57), .B(n_156), .Y(n_212) );
INVx1_ASAP7_75t_L g172 ( .A(n_59), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_60), .B(n_468), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_61), .B(n_500), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_62), .A2(n_158), .B(n_164), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_63), .B(n_156), .Y(n_167) );
INVx1_ASAP7_75t_L g146 ( .A(n_64), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_65), .A2(n_101), .B1(n_112), .B2(n_759), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_67), .B(n_169), .Y(n_479) );
AO32x2_ASAP7_75t_L g201 ( .A1(n_68), .A2(n_176), .A3(n_195), .B1(n_202), .B2(n_207), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_69), .B(n_170), .Y(n_518) );
INVx1_ASAP7_75t_L g191 ( .A(n_70), .Y(n_191) );
INVx1_ASAP7_75t_L g233 ( .A(n_71), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_72), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_73), .B(n_478), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_74), .A2(n_473), .B(n_481), .C(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_75), .B(n_152), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_76), .Y(n_545) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_78), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_79), .B(n_477), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_81), .B(n_204), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_82), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_83), .B(n_152), .Y(n_237) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_85), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_86), .B(n_194), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_87), .B(n_152), .Y(n_180) );
OR2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g455 ( .A(n_88), .B(n_122), .Y(n_455) );
INVx2_ASAP7_75t_L g459 ( .A(n_88), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_90), .A2(n_99), .B1(n_152), .B2(n_153), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_91), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g476 ( .A(n_92), .Y(n_476) );
INVxp67_ASAP7_75t_L g548 ( .A(n_93), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_94), .B(n_152), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g514 ( .A(n_96), .Y(n_514) );
INVx1_ASAP7_75t_L g572 ( .A(n_97), .Y(n_572) );
AND2x2_ASAP7_75t_L g539 ( .A(n_98), .B(n_197), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_104), .Y(n_760) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_126), .B1(n_752), .B2(n_754), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g753 ( .A(n_117), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_118), .A2(n_120), .B(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_121), .B(n_459), .Y(n_751) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g458 ( .A(n_122), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI22x1_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_453), .B1(n_456), .B2(n_460), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_129), .A2(n_453), .B1(n_458), .B2(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_130), .A2(n_131), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_418), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_322), .C(n_406), .Y(n_132) );
NAND4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_265), .C(n_287), .D(n_303), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_198), .B1(n_224), .B2(n_243), .C(n_251), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_174), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_137), .B(n_243), .Y(n_277) );
NAND4xp25_ASAP7_75t_L g317 ( .A(n_137), .B(n_305), .C(n_318), .D(n_320), .Y(n_317) );
INVxp67_ASAP7_75t_L g434 ( .A(n_137), .Y(n_434) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g316 ( .A(n_138), .B(n_254), .Y(n_316) );
AND2x2_ASAP7_75t_L g340 ( .A(n_138), .B(n_174), .Y(n_340) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g307 ( .A(n_139), .B(n_242), .Y(n_307) );
AND2x2_ASAP7_75t_L g347 ( .A(n_139), .B(n_328), .Y(n_347) );
AND2x2_ASAP7_75t_L g364 ( .A(n_139), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_139), .B(n_175), .Y(n_388) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g241 ( .A(n_140), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g259 ( .A(n_140), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g271 ( .A(n_140), .B(n_175), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_140), .B(n_185), .Y(n_293) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_148), .B(n_173), .Y(n_140) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_141), .A2(n_186), .B(n_196), .Y(n_185) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_142), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_144), .B(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_162), .B(n_171), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .C(n_158), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_151), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_151), .A2(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
INVx1_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
INVx3_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_156), .Y(n_574) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
AND2x6_ASAP7_75t_L g473 ( .A(n_157), .B(n_474), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_158), .A2(n_572), .B(n_573), .C(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_159), .A2(n_236), .B(n_237), .Y(n_235) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g478 ( .A(n_160), .Y(n_478) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g170 ( .A(n_161), .Y(n_170) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
AND2x2_ASAP7_75t_L g469 ( .A(n_161), .B(n_165), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_161), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_167), .C(n_168), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_L g190 ( .A1(n_163), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_163), .A2(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_168), .A2(n_182), .B(n_183), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_168), .A2(n_194), .B1(n_222), .B2(n_223), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_168), .A2(n_194), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_169), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_169), .A2(n_188), .B(n_189), .Y(n_187) );
O2A1O1Ixp5_ASAP7_75t_SL g231 ( .A1(n_169), .A2(n_232), .B(n_233), .C(n_234), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_169), .B(n_548), .Y(n_547) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_170), .A2(n_194), .B1(n_203), .B2(n_206), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_171), .A2(n_178), .B(n_181), .Y(n_177) );
BUFx3_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_171), .A2(n_211), .B(n_216), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_171), .A2(n_231), .B(n_235), .Y(n_230) );
AND2x4_ASAP7_75t_L g468 ( .A(n_171), .B(n_469), .Y(n_468) );
INVx4_ASAP7_75t_SL g482 ( .A(n_171), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_171), .B(n_469), .Y(n_515) );
AND2x2_ASAP7_75t_L g274 ( .A(n_174), .B(n_275), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_174), .A2(n_324), .B1(n_327), .B2(n_329), .C(n_333), .Y(n_323) );
AND2x2_ASAP7_75t_L g382 ( .A(n_174), .B(n_347), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_174), .B(n_364), .Y(n_416) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_185), .Y(n_174) );
INVx3_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
AND2x2_ASAP7_75t_L g291 ( .A(n_175), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g345 ( .A(n_175), .B(n_260), .Y(n_345) );
AND2x2_ASAP7_75t_L g403 ( .A(n_175), .B(n_404), .Y(n_403) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_184), .Y(n_175) );
INVx4_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_176), .A2(n_524), .B(n_525), .Y(n_523) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_176), .Y(n_542) );
AND2x2_ASAP7_75t_L g243 ( .A(n_185), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g260 ( .A(n_185), .Y(n_260) );
INVx1_ASAP7_75t_L g315 ( .A(n_185), .Y(n_315) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_185), .Y(n_321) );
AND2x2_ASAP7_75t_L g366 ( .A(n_185), .B(n_242), .Y(n_366) );
OR2x2_ASAP7_75t_L g405 ( .A(n_185), .B(n_244), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B(n_195), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_193), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx4_ASAP7_75t_L g507 ( .A(n_194), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g264 ( .A(n_195), .B(n_245), .C(n_246), .Y(n_264) );
INVx2_ASAP7_75t_L g207 ( .A(n_197), .Y(n_207) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_197), .A2(n_210), .B(n_219), .Y(n_209) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_230), .B(n_238), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_197), .A2(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g497 ( .A(n_197), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_197), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_198), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
AND2x2_ASAP7_75t_L g401 ( .A(n_199), .B(n_398), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_199), .B(n_383), .Y(n_433) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g332 ( .A(n_200), .B(n_256), .Y(n_332) );
AND2x2_ASAP7_75t_L g381 ( .A(n_200), .B(n_227), .Y(n_381) );
INVx1_ASAP7_75t_L g427 ( .A(n_200), .Y(n_427) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
AND2x2_ASAP7_75t_L g282 ( .A(n_201), .B(n_256), .Y(n_282) );
INVx1_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
AND2x2_ASAP7_75t_L g305 ( .A(n_201), .B(n_220), .Y(n_305) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_205), .Y(n_480) );
INVx2_ASAP7_75t_L g508 ( .A(n_205), .Y(n_508) );
INVx1_ASAP7_75t_L g494 ( .A(n_207), .Y(n_494) );
AND2x2_ASAP7_75t_L g373 ( .A(n_208), .B(n_281), .Y(n_373) );
INVx2_ASAP7_75t_L g438 ( .A(n_208), .Y(n_438) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AND2x2_ASAP7_75t_L g255 ( .A(n_209), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g268 ( .A(n_209), .B(n_228), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_209), .B(n_227), .Y(n_296) );
INVx1_ASAP7_75t_L g302 ( .A(n_209), .Y(n_302) );
INVx1_ASAP7_75t_L g319 ( .A(n_209), .Y(n_319) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_209), .Y(n_331) );
INVx2_ASAP7_75t_L g399 ( .A(n_209), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g256 ( .A(n_220), .Y(n_256) );
BUFx2_ASAP7_75t_L g353 ( .A(n_220), .Y(n_353) );
AND2x2_ASAP7_75t_L g398 ( .A(n_220), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_226), .B(n_335), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_226), .A2(n_397), .B(n_411), .Y(n_421) );
AND2x2_ASAP7_75t_L g446 ( .A(n_226), .B(n_332), .Y(n_446) );
BUFx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g368 ( .A(n_228), .Y(n_368) );
AND2x2_ASAP7_75t_L g397 ( .A(n_228), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_229), .Y(n_281) );
INVx2_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_229), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g254 ( .A(n_240), .Y(n_254) );
OR2x2_ASAP7_75t_L g267 ( .A(n_240), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g335 ( .A(n_240), .B(n_331), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_240), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g436 ( .A(n_240), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_240), .B(n_373), .Y(n_448) );
AND2x2_ASAP7_75t_L g327 ( .A(n_241), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_241), .B(n_243), .Y(n_350) );
INVx2_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
AND2x2_ASAP7_75t_L g290 ( .A(n_242), .B(n_263), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_242), .B(n_315), .Y(n_371) );
AND2x2_ASAP7_75t_L g285 ( .A(n_243), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g432 ( .A(n_243), .Y(n_432) );
AND2x2_ASAP7_75t_L g444 ( .A(n_243), .B(n_307), .Y(n_444) );
AND2x2_ASAP7_75t_L g270 ( .A(n_244), .B(n_260), .Y(n_270) );
INVx1_ASAP7_75t_L g365 ( .A(n_244), .Y(n_365) );
AO21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_249), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_245), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g500 ( .A(n_245), .Y(n_500) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_245), .A2(n_513), .B(n_520), .Y(n_512) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_245), .A2(n_569), .B(n_576), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_245), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g263 ( .A(n_250), .B(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_257), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_254), .B(n_301), .Y(n_310) );
OR2x2_ASAP7_75t_L g442 ( .A(n_254), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_300), .Y(n_359) );
AND2x2_ASAP7_75t_L g367 ( .A(n_255), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g426 ( .A(n_255), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g450 ( .A(n_255), .B(n_297), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_256), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g437 ( .A(n_256), .B(n_300), .Y(n_437) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g289 ( .A(n_259), .B(n_290), .Y(n_289) );
INVxp67_ASAP7_75t_L g451 ( .A(n_259), .Y(n_451) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
AND2x2_ASAP7_75t_L g337 ( .A(n_262), .B(n_270), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_262), .B(n_405), .Y(n_431) );
INVx2_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
INVx3_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
OR2x2_ASAP7_75t_L g356 ( .A(n_263), .B(n_357), .Y(n_356) );
AOI311xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .A3(n_271), .B(n_272), .C(n_283), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_266), .A2(n_304), .B(n_306), .C(n_308), .Y(n_303) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g288 ( .A(n_268), .Y(n_288) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_270), .B(n_286), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_270), .B(n_271), .Y(n_439) );
AND2x2_ASAP7_75t_L g361 ( .A(n_271), .B(n_275), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B(n_278), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g419 ( .A(n_275), .B(n_307), .Y(n_419) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_276), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g313 ( .A(n_276), .Y(n_313) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g349 ( .A(n_282), .Y(n_349) );
AND2x4_ASAP7_75t_L g411 ( .A(n_282), .B(n_380), .Y(n_411) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI222xp33_ASAP7_75t_L g362 ( .A1(n_285), .A2(n_351), .B1(n_363), .B2(n_367), .C1(n_369), .C2(n_373), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_291), .C(n_294), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_288), .B(n_332), .Y(n_355) );
INVx1_ASAP7_75t_L g377 ( .A(n_290), .Y(n_377) );
INVx1_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
OR2x2_ASAP7_75t_L g376 ( .A(n_293), .B(n_377), .Y(n_376) );
OAI21xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_301), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_295), .B(n_313), .C(n_314), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_295), .A2(n_332), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_300), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g409 ( .A(n_300), .Y(n_409) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
INVx2_ASAP7_75t_L g383 ( .A(n_301), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_305), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g357 ( .A(n_307), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_312), .B2(n_316), .C(n_317), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_311), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g445 ( .A(n_311), .Y(n_445) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g326 ( .A(n_318), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_318), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g384 ( .A(n_318), .B(n_332), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_318), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g417 ( .A(n_318), .B(n_352), .Y(n_417) );
BUFx3_ASAP7_75t_L g380 ( .A(n_319), .Y(n_380) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND5xp2_ASAP7_75t_L g322 ( .A(n_323), .B(n_341), .C(n_362), .D(n_374), .E(n_389), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI32xp33_ASAP7_75t_L g414 ( .A1(n_326), .A2(n_353), .A3(n_369), .B1(n_415), .B2(n_417), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_328), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g338 ( .A(n_332), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B1(n_338), .B2(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_348), .B1(n_350), .B2(n_351), .C(n_354), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g413 ( .A(n_345), .B(n_364), .Y(n_413) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_350), .A2(n_411), .B1(n_429), .B2(n_434), .C(n_435), .Y(n_428) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g372 ( .A(n_364), .Y(n_372) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_382), .B2(n_383), .C1(n_384), .C2(n_385), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_430), .B1(n_432), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_395), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_400), .B(n_402), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B(n_412), .C(n_414), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_422), .C(n_447), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_419), .Y(n_423) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_428), .C(n_440), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B(n_439), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g748 ( .A(n_460), .Y(n_748) );
OR3x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_660), .C(n_703), .Y(n_460) );
NAND5xp2_ASAP7_75t_L g461 ( .A(n_462), .B(n_587), .C(n_617), .D(n_634), .E(n_649), .Y(n_461) );
AOI221xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_510), .B1(n_550), .B2(n_556), .C(n_560), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_485), .Y(n_463) );
OR2x2_ASAP7_75t_L g565 ( .A(n_464), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g622 ( .A(n_464), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_464), .B(n_558), .Y(n_639) );
OR2x2_ASAP7_75t_L g651 ( .A(n_464), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_464), .B(n_610), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_464), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_464), .B(n_588), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_464), .B(n_596), .Y(n_702) );
AND2x2_ASAP7_75t_L g734 ( .A(n_464), .B(n_498), .Y(n_734) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_464), .Y(n_742) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_465), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g562 ( .A(n_465), .B(n_540), .Y(n_562) );
BUFx2_ASAP7_75t_L g584 ( .A(n_465), .Y(n_584) );
AND2x2_ASAP7_75t_L g613 ( .A(n_465), .B(n_486), .Y(n_613) );
AND2x2_ASAP7_75t_L g668 ( .A(n_465), .B(n_566), .Y(n_668) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_483), .Y(n_465) );
BUFx2_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_472), .A2(n_482), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_472), .A2(n_482), .B(n_545), .C(n_546), .Y(n_544) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_479), .C(n_480), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_480), .B(n_537), .C(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_485), .B(n_622), .Y(n_631) );
OAI32xp33_ASAP7_75t_L g645 ( .A1(n_485), .A2(n_581), .A3(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_485), .B(n_647), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_485), .B(n_565), .Y(n_688) );
INVx1_ASAP7_75t_SL g717 ( .A(n_485), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_485), .B(n_512), .C(n_668), .D(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .Y(n_485) );
INVx5_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_499), .Y(n_588) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_486), .Y(n_667) );
AND2x2_ASAP7_75t_L g737 ( .A(n_486), .B(n_684), .Y(n_737) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_490), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g610 ( .A(n_498), .B(n_559), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_498), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g644 ( .A(n_498), .B(n_566), .Y(n_644) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g558 ( .A(n_499), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_568), .Y(n_596) );
AND2x2_ASAP7_75t_L g605 ( .A(n_499), .B(n_567), .Y(n_605) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_509), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_510), .A2(n_674), .B1(n_676), .B2(n_678), .C1(n_681), .C2(n_682), .Y(n_673) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_529), .Y(n_510) );
AND2x2_ASAP7_75t_L g606 ( .A(n_511), .B(n_607), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_511), .B(n_584), .C(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
INVx5_ASAP7_75t_SL g555 ( .A(n_512), .Y(n_555) );
OAI322xp33_ASAP7_75t_L g560 ( .A1(n_512), .A2(n_561), .A3(n_563), .B1(n_564), .B2(n_578), .C1(n_581), .C2(n_583), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_512), .B(n_553), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_512), .B(n_541), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g553 ( .A(n_522), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_522), .B(n_531), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_529), .B(n_591), .Y(n_646) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g625 ( .A(n_530), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
OR2x2_ASAP7_75t_L g554 ( .A(n_531), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_531), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g593 ( .A(n_531), .B(n_541), .Y(n_593) );
AND2x2_ASAP7_75t_L g616 ( .A(n_531), .B(n_553), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_531), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_531), .B(n_591), .Y(n_632) );
AND2x2_ASAP7_75t_L g640 ( .A(n_531), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_531), .B(n_600), .Y(n_690) );
INVx5_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g580 ( .A(n_532), .B(n_555), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_532), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g607 ( .A(n_532), .B(n_541), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_532), .B(n_654), .Y(n_695) );
OR2x2_ASAP7_75t_L g711 ( .A(n_532), .B(n_655), .Y(n_711) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_532), .B(n_672), .Y(n_718) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_532), .Y(n_725) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_L g579 ( .A(n_540), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g629 ( .A(n_540), .B(n_553), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_540), .B(n_555), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_540), .B(n_591), .Y(n_713) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_541), .B(n_555), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_541), .B(n_553), .Y(n_601) );
OR2x2_ASAP7_75t_L g655 ( .A(n_541), .B(n_553), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_541), .B(n_552), .Y(n_672) );
INVxp67_ASAP7_75t_L g694 ( .A(n_541), .Y(n_694) );
AND2x2_ASAP7_75t_L g721 ( .A(n_541), .B(n_591), .Y(n_721) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_541), .Y(n_728) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_552), .B(n_602), .Y(n_675) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_555), .Y(n_591) );
OR2x2_ASAP7_75t_L g658 ( .A(n_553), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
OR2x2_ASAP7_75t_L g663 ( .A(n_554), .B(n_655), .Y(n_663) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g563 ( .A(n_558), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_558), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g564 ( .A(n_559), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_559), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_559), .B(n_566), .Y(n_598) );
INVx2_ASAP7_75t_L g643 ( .A(n_559), .Y(n_643) );
AND2x2_ASAP7_75t_L g656 ( .A(n_559), .B(n_596), .Y(n_656) );
AND2x2_ASAP7_75t_L g681 ( .A(n_559), .B(n_605), .Y(n_681) );
INVx1_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
INVx2_ASAP7_75t_SL g620 ( .A(n_565), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_567), .Y(n_586) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g684 ( .A(n_568), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g653 ( .A(n_580), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_580), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_580), .A2(n_662), .B1(n_664), .B2(n_669), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_580), .B(n_672), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_581), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g615 ( .A(n_582), .Y(n_615) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g597 ( .A(n_584), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_584), .B(n_588), .Y(n_648) );
AND2x2_ASAP7_75t_L g671 ( .A(n_584), .B(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g647 ( .A(n_586), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_594), .C(n_608), .Y(n_587) );
INVx1_ASAP7_75t_L g611 ( .A(n_588), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g719 ( .A1(n_588), .A2(n_720), .B1(n_722), .B2(n_723), .C(n_726), .Y(n_719) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g738 ( .A(n_591), .Y(n_738) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g687 ( .A(n_593), .B(n_626), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_599), .C(n_603), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_601), .A2(n_602), .A3(n_665), .B1(n_702), .B2(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
AND2x2_ASAP7_75t_L g744 ( .A(n_604), .B(n_643), .Y(n_744) );
AND2x2_ASAP7_75t_L g691 ( .A(n_605), .B(n_643), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_605), .B(n_613), .Y(n_709) );
AOI31xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .A3(n_612), .B(n_614), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_610), .B(n_622), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_610), .B(n_620), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_610), .A2(n_640), .B1(n_730), .B2(n_733), .C(n_735), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g635 ( .A(n_615), .B(n_636), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_624), .B1(n_627), .B2(n_630), .C1(n_632), .C2(n_633), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g700 ( .A(n_619), .Y(n_700) );
INVx1_ASAP7_75t_L g722 ( .A(n_622), .Y(n_722) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_625), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g641 ( .A(n_626), .Y(n_641) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B1(n_640), .B2(n_642), .C(n_645), .Y(n_634) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g679 ( .A(n_637), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g731 ( .A(n_637), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g706 ( .A(n_642), .Y(n_706) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g670 ( .A(n_643), .Y(n_670) );
INVx1_ASAP7_75t_L g652 ( .A(n_644), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_647), .B(n_734), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_656), .B2(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g743 ( .A(n_656), .Y(n_743) );
INVxp33_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_658), .B(n_702), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g692 ( .A1(n_659), .A2(n_693), .A3(n_694), .B1(n_695), .B2(n_696), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_673), .C(n_685), .D(n_697), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NAND2xp33_ASAP7_75t_SL g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_668), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
CKINVDCx16_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_682), .A2(n_698), .B1(n_715), .B2(n_718), .C(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g733 ( .A(n_684), .B(n_734), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_689), .B2(n_691), .C(n_692), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_694), .B(n_725), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_704), .B(n_714), .C(n_729), .D(n_740), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B(n_710), .C(n_712), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g745 ( .A(n_732), .Y(n_745) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_744), .B(n_745), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
endmodule