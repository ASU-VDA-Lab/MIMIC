module fake_jpeg_18938_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_44),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_21),
.B(n_22),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_42),
.Y(n_81)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_23),
.B1(n_19),
.B2(n_30),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_23),
.B1(n_19),
.B2(n_41),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_42),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_81),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_78),
.B1(n_38),
.B2(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_41),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_38),
.B1(n_58),
.B2(n_51),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_42),
.B(n_39),
.C(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_39),
.B1(n_34),
.B2(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_42),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_38),
.B1(n_57),
.B2(n_40),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_36),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_36),
.B(n_24),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_79),
.B(n_75),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_60),
.B1(n_53),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_101),
.B1(n_78),
.B2(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_49),
.B1(n_58),
.B2(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_73),
.B1(n_66),
.B2(n_87),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_111),
.B1(n_86),
.B2(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_72),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_113),
.B1(n_52),
.B2(n_40),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_31),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_140),
.B1(n_97),
.B2(n_96),
.Y(n_146)
);

OAI21x1_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_96),
.B(n_81),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_120),
.B(n_126),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_124),
.B(n_138),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_100),
.B(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_136),
.B1(n_142),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_86),
.B1(n_75),
.B2(n_73),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_132),
.B1(n_139),
.B2(n_89),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_63),
.B1(n_70),
.B2(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_73),
.B1(n_31),
.B2(n_16),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_101),
.B1(n_97),
.B2(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_40),
.B1(n_52),
.B2(n_32),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_113),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_94),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_140),
.B1(n_117),
.B2(n_128),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_100),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_90),
.C(n_94),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_25),
.C(n_88),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_90),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_112),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_126),
.B(n_135),
.C(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_143),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_166),
.B(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_109),
.A3(n_107),
.B1(n_27),
.B2(n_32),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_28),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_91),
.B(n_27),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_99),
.B1(n_106),
.B2(n_95),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_106),
.B(n_1),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_87),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_171),
.B(n_21),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_151),
.B1(n_166),
.B2(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_184),
.B1(n_189),
.B2(n_190),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_152),
.C(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_185),
.B(n_197),
.Y(n_203)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_143),
.B1(n_93),
.B2(n_125),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_93),
.B1(n_87),
.B2(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_88),
.B1(n_69),
.B2(n_28),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_199),
.B1(n_148),
.B2(n_172),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_196),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_153),
.A3(n_169),
.B1(n_160),
.B2(n_159),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_176),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_21),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_212),
.C(n_223),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_188),
.B1(n_190),
.B2(n_189),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_208),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_150),
.B1(n_169),
.B2(n_163),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_210),
.B1(n_214),
.B2(n_191),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_213),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_159),
.B1(n_170),
.B2(n_164),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_156),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_211),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_165),
.B1(n_155),
.B2(n_26),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_155),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_25),
.C(n_26),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_15),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_2),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_208),
.B1(n_219),
.B2(n_223),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_183),
.B1(n_187),
.B2(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_240),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_183),
.B1(n_199),
.B2(n_182),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_192),
.C(n_175),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_239),
.C(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_173),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_196),
.B1(n_177),
.B2(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_175),
.C(n_173),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_243),
.B1(n_231),
.B2(n_230),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_217),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_209),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_249),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_207),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_204),
.B(n_191),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_250),
.B(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_235),
.B(n_233),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_239),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_256),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_214),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_241),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_8),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_269),
.B1(n_270),
.B2(n_13),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_224),
.B(n_226),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_267),
.B(n_6),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_225),
.C(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_266),
.C(n_7),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_232),
.C(n_229),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_201),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_7),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_245),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_249),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_262),
.B(n_282),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_256),
.B1(n_253),
.B2(n_257),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_248),
.B(n_7),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_263),
.B(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_291)
);

OAI221xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_8),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_265),
.C(n_260),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_260),
.C(n_262),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_268),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_278),
.B(n_284),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_299),
.B(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_300),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_9),
.B(n_11),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_11),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_12),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_12),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_292),
.C(n_12),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_296),
.B(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_298),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_13),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_13),
.Y(n_311)
);


endmodule