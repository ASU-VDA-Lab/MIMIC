module real_jpeg_24336_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_2),
.A2(n_19),
.B1(n_26),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_30),
.B1(n_32),
.B2(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_30),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_62),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_30),
.C(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_34),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_19),
.B1(n_26),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_9),
.A2(n_22),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_9),
.A2(n_19),
.B1(n_26),
.B2(n_64),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_30),
.B1(n_32),
.B2(n_64),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_74),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_65),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_65),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_42),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_21),
.C(n_25),
.Y(n_17)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_18),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_18),
.A2(n_22),
.B1(n_27),
.B2(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_19),
.A2(n_26),
.B1(n_50),
.B2(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_21),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_24),
.CON(n_21),
.SN(n_21)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_26),
.C(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_24),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_36),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_32),
.B1(n_50),
.B2(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_33),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_34),
.A2(n_37),
.B1(n_91),
.B2(n_99),
.Y(n_107)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_35),
.Y(n_92)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_57),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_48),
.B1(n_53),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_53),
.B1(n_67),
.B2(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.C(n_70),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_87),
.B(n_110),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_96),
.B(n_109),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_94),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_105),
.B(n_108),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_106),
.B(n_107),
.Y(n_108)
);


endmodule