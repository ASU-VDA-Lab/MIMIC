module fake_jpeg_31679_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_24),
.B(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_68),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_24),
.A2(n_14),
.B(n_5),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_5),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_89),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_2),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_34),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_94),
.Y(n_156)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_99),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_45),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_46),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_30),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_102),
.A2(n_107),
.B1(n_125),
.B2(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_26),
.B1(n_40),
.B2(n_38),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_40),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_26),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_36),
.B(n_41),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_27),
.C(n_19),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_45),
.B1(n_49),
.B2(n_48),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_53),
.B(n_30),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_145),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_63),
.B(n_42),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_55),
.B(n_47),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_66),
.A2(n_38),
.B1(n_42),
.B2(n_48),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_41),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_43),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_84),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_62),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_163),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_74),
.B1(n_96),
.B2(n_75),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_162),
.A2(n_179),
.B1(n_158),
.B2(n_122),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_173),
.Y(n_227)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_85),
.B1(n_83),
.B2(n_76),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_167),
.A2(n_204),
.B1(n_125),
.B2(n_120),
.Y(n_232)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_43),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

OR2x4_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_44),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_181),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_95),
.B1(n_91),
.B2(n_48),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_82),
.B1(n_88),
.B2(n_59),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_49),
.C(n_44),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_183),
.B(n_208),
.Y(n_234)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_153),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_196),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_114),
.Y(n_187)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_197),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g193 ( 
.A(n_130),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_46),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_207),
.B1(n_155),
.B2(n_156),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.Y(n_211)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_111),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_44),
.B(n_33),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_132),
.A2(n_147),
.B1(n_123),
.B2(n_127),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_102),
.A2(n_49),
.B1(n_99),
.B2(n_94),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_129),
.B1(n_122),
.B2(n_138),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_146),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_155),
.Y(n_216)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_216),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_168),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_141),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_120),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_232),
.A2(n_188),
.B1(n_229),
.B2(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_205),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_137),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_237),
.B(n_246),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_187),
.B(n_33),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_245),
.B1(n_185),
.B2(n_129),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_121),
.B1(n_138),
.B2(n_133),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_164),
.B(n_104),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_31),
.B(n_21),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_33),
.B(n_31),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_182),
.C(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_254),
.C(n_208),
.Y(n_313)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_168),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_273),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_195),
.B1(n_184),
.B2(n_174),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_182),
.C(n_169),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_272),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_233),
.B1(n_213),
.B2(n_223),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_188),
.B1(n_190),
.B2(n_167),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_262),
.B1(n_275),
.B2(n_281),
.Y(n_293)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_211),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_265),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_211),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_219),
.B1(n_233),
.B2(n_246),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_160),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_187),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_19),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_177),
.B1(n_121),
.B2(n_124),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_278),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_214),
.A2(n_192),
.B(n_163),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_240),
.B(n_210),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_176),
.Y(n_278)
);

BUFx4f_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_216),
.B(n_199),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_240),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_215),
.A2(n_166),
.B1(n_198),
.B2(n_191),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_225),
.A2(n_171),
.B1(n_202),
.B2(n_170),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_295),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_214),
.A3(n_243),
.B1(n_247),
.B2(n_221),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_289),
.A2(n_270),
.B(n_276),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_294),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_262),
.A2(n_241),
.B1(n_222),
.B2(n_231),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_221),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_297),
.B(n_308),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_257),
.A2(n_222),
.B1(n_238),
.B2(n_231),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_222),
.B1(n_213),
.B2(n_226),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_272),
.A2(n_223),
.B1(n_226),
.B2(n_189),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_283),
.B(n_252),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_250),
.B(n_210),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_224),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_309),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_250),
.B(n_217),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_311),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_312),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.C(n_277),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_248),
.C(n_254),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_255),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_339),
.C(n_346),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_316),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_263),
.Y(n_320)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_255),
.B(n_274),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_328),
.B(n_345),
.Y(n_364)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_310),
.B(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_336),
.B(n_299),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_290),
.A2(n_252),
.B(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_333),
.B(n_220),
.Y(n_384)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_275),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_300),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_286),
.A2(n_280),
.B(n_270),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_310),
.B(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_259),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_340),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_212),
.C(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_344),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_291),
.B(n_224),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_279),
.C(n_288),
.Y(n_367)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_286),
.A2(n_256),
.B(n_267),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_286),
.C(n_306),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_212),
.B1(n_260),
.B2(n_194),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_349),
.Y(n_381)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_293),
.A2(n_258),
.B1(n_242),
.B2(n_249),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_350),
.A2(n_288),
.B1(n_314),
.B2(n_258),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_319),
.B(n_328),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_359),
.B1(n_345),
.B2(n_324),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_284),
.B1(n_292),
.B2(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

AOI32xp33_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_316),
.A3(n_301),
.B1(n_302),
.B2(n_295),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_330),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_287),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_377),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_329),
.B(n_279),
.CI(n_302),
.CON(n_362),
.SN(n_362)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_375),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_314),
.C(n_307),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_368),
.C(n_341),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_331),
.B(n_279),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_366),
.B(n_376),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_367),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_307),
.C(n_299),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_370),
.A2(n_373),
.B(n_330),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_230),
.Y(n_372)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_220),
.B(n_298),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_201),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_337),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_378),
.B(n_349),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_266),
.Y(n_382)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_384),
.B(n_348),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_392),
.C(n_398),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_386),
.A2(n_369),
.B1(n_379),
.B2(n_380),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_401),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_397),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_336),
.C(n_351),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_364),
.A2(n_370),
.B(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_375),
.A2(n_347),
.B1(n_319),
.B2(n_350),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_362),
.Y(n_422)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_363),
.B(n_344),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_347),
.C(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_323),
.C(n_335),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_406),
.C(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_371),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_407),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_334),
.C(n_230),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_408),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_409),
.B(n_381),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_261),
.C(n_186),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_244),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_412),
.B(n_380),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_352),
.Y(n_421)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_392),
.B(n_352),
.CI(n_384),
.CON(n_416),
.SN(n_416)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_364),
.C(n_355),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_423),
.C(n_429),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_422),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_362),
.C(n_374),
.Y(n_423)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_395),
.C(n_389),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_413),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_427),
.A2(n_394),
.B1(n_402),
.B2(n_390),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_382),
.C(n_369),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_405),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_381),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_435),
.C(n_325),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_365),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_437),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_410),
.C(n_401),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_322),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_414),
.A2(n_388),
.B1(n_399),
.B2(n_408),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_450),
.B1(n_454),
.B2(n_419),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_389),
.B(n_409),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_443),
.A2(n_435),
.B(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_436),
.Y(n_445)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_431),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_452),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_432),
.A2(n_390),
.B(n_387),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_449),
.A2(n_420),
.B(n_416),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_421),
.A2(n_325),
.B1(n_322),
.B2(n_249),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_456),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_415),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g454 ( 
.A1(n_423),
.A2(n_244),
.B1(n_207),
.B2(n_200),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_429),
.B(n_126),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_448),
.B1(n_438),
.B2(n_134),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_463),
.B(n_448),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_418),
.C(n_417),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_466),
.C(n_467),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_418),
.C(n_417),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_433),
.C(n_106),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_106),
.C(n_126),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_455),
.C(n_446),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_443),
.B(n_27),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_471),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_443),
.B(n_21),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_21),
.Y(n_473)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_440),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_478),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_468),
.B(n_453),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_459),
.B(n_449),
.Y(n_479)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_441),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_481),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_441),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_439),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_483),
.B(n_486),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_50),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_134),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_460),
.C(n_465),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_SL g490 ( 
.A(n_485),
.B(n_463),
.C(n_461),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_493),
.Y(n_505)
);

NOR2x1_ASAP7_75t_SL g492 ( 
.A(n_474),
.B(n_460),
.Y(n_492)
);

AOI31xp67_ASAP7_75t_L g500 ( 
.A1(n_492),
.A2(n_496),
.A3(n_484),
.B(n_476),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_481),
.A2(n_465),
.B(n_482),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_467),
.C(n_469),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_489),
.Y(n_501)
);

AOI21x1_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_496),
.B(n_499),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_502),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_475),
.Y(n_502)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_78),
.A3(n_65),
.B1(n_46),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_503)
);

AOI321xp33_ASAP7_75t_SL g508 ( 
.A1(n_503),
.A2(n_504),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_78),
.A3(n_65),
.B1(n_46),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_498),
.C(n_490),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_5),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_506),
.C(n_46),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_509),
.A2(n_510),
.B(n_505),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_512),
.Y(n_513)
);

AOI322xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_507),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_7),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_9),
.C(n_12),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_12),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_13),
.Y(n_517)
);


endmodule