module fake_jpeg_12923_n_398 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_398);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_398;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_57),
.B(n_75),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_63),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g154 ( 
.A(n_59),
.Y(n_154)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_12),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_66),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_20),
.B(n_4),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_6),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_91),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_24),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_96),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_33),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_33),
.A2(n_7),
.B(n_8),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_97),
.B(n_98),
.C(n_44),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_7),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx5_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_32),
.B(n_9),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_12),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_41),
.Y(n_143)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_108),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_37),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_61),
.B1(n_69),
.B2(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_111),
.A2(n_132),
.B1(n_142),
.B2(n_150),
.Y(n_218)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_32),
.Y(n_117)
);

NAND4xp25_ASAP7_75t_L g217 ( 
.A(n_117),
.B(n_154),
.C(n_116),
.D(n_142),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_45),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_119),
.B(n_130),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_67),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_56),
.B1(n_42),
.B2(n_43),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_41),
.B1(n_53),
.B2(n_52),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_144),
.B1(n_44),
.B2(n_30),
.Y(n_191)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_73),
.A2(n_48),
.B1(n_28),
.B2(n_54),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_172),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_74),
.A2(n_53),
.B1(n_52),
.B2(n_47),
.Y(n_144)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_60),
.A2(n_28),
.B1(n_54),
.B2(n_36),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_36),
.B1(n_46),
.B2(n_43),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_168),
.B1(n_59),
.B2(n_90),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_76),
.A2(n_28),
.B1(n_51),
.B2(n_38),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_156),
.A2(n_170),
.B1(n_126),
.B2(n_113),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_98),
.B(n_47),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_45),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_167),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_81),
.A2(n_35),
.B1(n_46),
.B2(n_42),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_100),
.A2(n_51),
.B1(n_30),
.B2(n_35),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_111),
.A2(n_106),
.B1(n_104),
.B2(n_94),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_175),
.A2(n_190),
.B1(n_193),
.B2(n_220),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_179),
.Y(n_230)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_131),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_38),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_196),
.Y(n_241)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_185),
.B(n_195),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_186),
.B(n_189),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_115),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_85),
.B1(n_113),
.B2(n_165),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_93),
.B1(n_86),
.B2(n_29),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_83),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_13),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_83),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_197),
.B(n_206),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_138),
.B1(n_163),
.B2(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_13),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_204),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_212),
.Y(n_233)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_14),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_117),
.A2(n_90),
.B1(n_92),
.B2(n_16),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_205),
.A2(n_214),
.B(n_224),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_17),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_17),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_213),
.B(n_215),
.Y(n_273)
);

OR2x4_ASAP7_75t_L g214 ( 
.A(n_114),
.B(n_129),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_125),
.B(n_152),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_137),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_216),
.B(n_219),
.Y(n_264)
);

NAND2x1_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_205),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_134),
.B(n_146),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_150),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_222),
.B(n_227),
.Y(n_269)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_226),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_135),
.A2(n_171),
.B1(n_174),
.B2(n_141),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_126),
.A2(n_135),
.B1(n_171),
.B2(n_166),
.Y(n_225)
);

AOI22x1_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_183),
.B1(n_217),
.B2(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_120),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_174),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_141),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_221),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_154),
.A2(n_159),
.B(n_136),
.C(n_138),
.Y(n_229)
);

AOI22x1_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_221),
.B1(n_226),
.B2(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_239),
.B1(n_269),
.B2(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_163),
.B1(n_222),
.B2(n_227),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_242),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_184),
.B(n_181),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_252),
.C(n_258),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_249),
.A2(n_232),
.B(n_233),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_191),
.A2(n_182),
.B1(n_193),
.B2(n_204),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_253),
.B1(n_254),
.B2(n_262),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_196),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_200),
.A2(n_224),
.B1(n_186),
.B2(n_214),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_184),
.A2(n_211),
.B1(n_192),
.B2(n_178),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_255),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_201),
.C(n_198),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_208),
.A2(n_203),
.A3(n_198),
.B1(n_202),
.B2(n_188),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_177),
.B(n_202),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_212),
.A2(n_180),
.B1(n_187),
.B2(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_194),
.A2(n_222),
.B1(n_227),
.B2(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_268),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_176),
.B(n_179),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_266),
.Y(n_274)
);

AO22x1_ASAP7_75t_SL g268 ( 
.A1(n_218),
.A2(n_222),
.B1(n_227),
.B2(n_217),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_238),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_283),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_282),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_279),
.B1(n_297),
.B2(n_296),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_271),
.B(n_249),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_278),
.A2(n_286),
.B(n_300),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_239),
.A2(n_234),
.B1(n_268),
.B2(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_244),
.B(n_264),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_248),
.B(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_248),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_286),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_254),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_235),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_272),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_248),
.A2(n_243),
.B1(n_242),
.B2(n_255),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_237),
.A2(n_273),
.B(n_258),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_247),
.A2(n_255),
.B(n_267),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_231),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_241),
.A2(n_230),
.B(n_232),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_288),
.B(n_282),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_240),
.C(n_235),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_284),
.C(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_275),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_240),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_316),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_262),
.B(n_270),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_306),
.A2(n_289),
.B(n_296),
.C(n_290),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_309),
.A2(n_314),
.B1(n_322),
.B2(n_274),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_310),
.A2(n_283),
.B(n_299),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_231),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_313),
.B(n_319),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_278),
.B(n_298),
.C(n_287),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_281),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_279),
.B1(n_297),
.B2(n_285),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_274),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_301),
.B(n_291),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_335),
.B(n_339),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_337),
.Y(n_346)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

AO22x1_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_310),
.B1(n_323),
.B2(n_315),
.Y(n_351)
);

AO221x1_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_303),
.B1(n_294),
.B2(n_299),
.C(n_295),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_325),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_343),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_305),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_323),
.B1(n_307),
.B2(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_357),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_318),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_316),
.C(n_315),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_352),
.C(n_327),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_325),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_350),
.B(n_353),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_351),
.A2(n_318),
.B(n_336),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_317),
.C(n_326),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_332),
.Y(n_353)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_362),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_354),
.A2(n_329),
.B(n_339),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_361),
.B(n_365),
.Y(n_370)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_369),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_354),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_349),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_368),
.A2(n_355),
.B1(n_340),
.B2(n_344),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_327),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_347),
.C(n_352),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_372),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_335),
.C(n_308),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_375),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_367),
.A2(n_357),
.B1(n_306),
.B2(n_322),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_370),
.B(n_361),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_365),
.B(n_320),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_343),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_358),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_375),
.C(n_366),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_371),
.B(n_369),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_374),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_385),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_370),
.A2(n_360),
.B(n_367),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_374),
.C(n_384),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_390),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_377),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_356),
.C(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_391),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_393),
.B1(n_388),
.B2(n_386),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_351),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_379),
.C(n_314),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_396),
.B(n_397),
.Y(n_398)
);


endmodule