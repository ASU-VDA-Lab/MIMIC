module fake_netlist_6_4284_n_1986 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1986);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1986;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_67),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_8),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_63),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_31),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_29),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_68),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_113),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_31),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_59),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_64),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_96),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_92),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_58),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_70),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_44),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_126),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_86),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_142),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_137),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_64),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_104),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_72),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_79),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_118),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_88),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_125),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_71),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_123),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_85),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_147),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_141),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_52),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_52),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_8),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_45),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_94),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_115),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_183),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_171),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_149),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_3),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_179),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_103),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_63),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_162),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_89),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_73),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_121),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_166),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_51),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_164),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_28),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_95),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_60),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_93),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_54),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_161),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_18),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_49),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_131),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_135),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_143),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_75),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_51),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_74),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_134),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_100),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_34),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

BUFx8_ASAP7_75t_SL g309 ( 
.A(n_98),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_128),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_119),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_151),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_44),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_20),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_48),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_114),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_150),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_163),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_155),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_34),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_26),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_20),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_146),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_152),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_76),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_169),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_12),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_132),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_154),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_173),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_30),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_33),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_139),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_185),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_12),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_111),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_110),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_90),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_124),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_167),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_160),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_60),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_0),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_45),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_37),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_116),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_186),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_9),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_129),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_97),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_39),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_11),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_40),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_182),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_23),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_11),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_32),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_14),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_24),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_105),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_80),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_159),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_170),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_43),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_61),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_57),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_24),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_50),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_156),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_27),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_18),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_133),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_81),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_62),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_77),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_83),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_42),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_3),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_22),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_309),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_351),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_359),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_248),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_197),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_249),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_244),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_196),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_244),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_244),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_244),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_244),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_293),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_293),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_296),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_294),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_293),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_293),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_293),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_253),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_253),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_205),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_205),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_203),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_198),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_247),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_250),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_201),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_215),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_251),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_302),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_266),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_252),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_221),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_254),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_266),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_231),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_268),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_305),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_255),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_270),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_232),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_241),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_246),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_203),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_273),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_206),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_333),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_283),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_206),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_306),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_333),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_336),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_284),
.Y(n_459)
);

INVxp33_ASAP7_75t_SL g460 ( 
.A(n_208),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_266),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_256),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_267),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_288),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_333),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_208),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_269),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_333),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_292),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_295),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_298),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_230),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_303),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_271),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_313),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_209),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_275),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_321),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_347),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_209),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_333),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_442),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_390),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_401),
.B(n_277),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_401),
.B(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_403),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_404),
.B(n_305),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_405),
.B(n_277),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

CKINVDCx8_ASAP7_75t_R g491 ( 
.A(n_402),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_398),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_406),
.B(n_194),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_394),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_406),
.B(n_194),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_407),
.B(n_207),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

CKINVDCx11_ASAP7_75t_R g501 ( 
.A(n_426),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_400),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_442),
.B(n_199),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_404),
.B(n_343),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_472),
.A2(n_349),
.B1(n_331),
.B2(n_376),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_411),
.B(n_207),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_421),
.B(n_423),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_433),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_410),
.A2(n_384),
.B1(n_220),
.B2(n_376),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_228),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_439),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_389),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_387),
.A2(n_257),
.B(n_226),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_439),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_445),
.A2(n_384),
.B1(n_220),
.B2(n_373),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_387),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_439),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_229),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_439),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_431),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_461),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_388),
.Y(n_539)
);

CKINVDCx8_ASAP7_75t_R g540 ( 
.A(n_446),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_421),
.B(n_199),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_395),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_461),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_396),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_396),
.B(n_343),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_397),
.B(n_210),
.Y(n_552)
);

CKINVDCx8_ASAP7_75t_R g553 ( 
.A(n_446),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_386),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_397),
.B(n_210),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_423),
.B(n_241),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_434),
.B(n_211),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_399),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_551),
.A2(n_447),
.B1(n_409),
.B2(n_480),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_483),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_499),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_501),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_527),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_482),
.B(n_438),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_532),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

BUFx8_ASAP7_75t_SL g573 ( 
.A(n_494),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_507),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_507),
.B(n_482),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_527),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_539),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_392),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_521),
.B(n_392),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_499),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_541),
.B(n_416),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_534),
.B(n_432),
.Y(n_585)
);

NOR2x1p5_ASAP7_75t_L g586 ( 
.A(n_484),
.B(n_214),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_539),
.Y(n_589)
);

INVxp67_ASAP7_75t_R g590 ( 
.A(n_500),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_490),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_559),
.B(n_432),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_552),
.B(n_480),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_496),
.B(n_462),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_547),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_555),
.Y(n_604)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_503),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_550),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_507),
.B(n_463),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_510),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_458),
.C(n_427),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_420),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_487),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_504),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_552),
.B(n_467),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_493),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_493),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_527),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_424),
.Y(n_621)
);

BUFx4f_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_424),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_502),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_502),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_537),
.B(n_474),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_517),
.B(n_415),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_518),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_505),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_560),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_556),
.B(n_451),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_505),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_509),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_517),
.B(n_415),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_556),
.B(n_477),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_540),
.B(n_454),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_551),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_557),
.B(n_348),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_551),
.B(n_488),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_495),
.B(n_460),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_513),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_513),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_546),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_516),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_551),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_488),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_519),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_530),
.A2(n_476),
.B1(n_466),
.B2(n_356),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_522),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_522),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_540),
.B(n_241),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_553),
.B(n_211),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_529),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_553),
.B(n_530),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_518),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_495),
.B(n_441),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_520),
.B(n_213),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_486),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_491),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_506),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_542),
.A2(n_257),
.B1(n_279),
.B2(n_226),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_542),
.B(n_512),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_488),
.B(n_386),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_520),
.B(n_213),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_488),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_497),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_486),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_511),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_497),
.B(n_498),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_511),
.B(n_425),
.Y(n_680)
);

BUFx6f_ASAP7_75t_SL g681 ( 
.A(n_511),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_526),
.A2(n_368),
.B1(n_327),
.B2(n_453),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_491),
.B(n_216),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_508),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_518),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_518),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_491),
.B(n_216),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_498),
.B(n_386),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_514),
.B(n_456),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_514),
.B(n_417),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_508),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_485),
.A2(n_350),
.B1(n_362),
.B2(n_335),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_508),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_485),
.A2(n_358),
.B1(n_380),
.B2(n_323),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_492),
.B(n_280),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_523),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_SL g697 ( 
.A(n_489),
.B(n_383),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_525),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_489),
.B(n_224),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_525),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_525),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_492),
.A2(n_375),
.B1(n_337),
.B2(n_332),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_525),
.B(n_224),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_492),
.B(n_515),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_492),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_523),
.B(n_214),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_515),
.B(n_225),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_523),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_525),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_515),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_538),
.A2(n_357),
.B1(n_372),
.B2(n_364),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_515),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_525),
.Y(n_713)
);

OAI221xp5_ASAP7_75t_L g714 ( 
.A1(n_694),
.A2(n_324),
.B1(n_354),
.B2(n_361),
.C(n_377),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_677),
.B(n_538),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_638),
.B(n_538),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_665),
.A2(n_366),
.B1(n_279),
.B2(n_334),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_573),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_678),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_595),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_619),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_608),
.B(n_336),
.Y(n_722)
);

BUFx5_ASAP7_75t_L g723 ( 
.A(n_641),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_644),
.B(n_225),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_678),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_595),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_651),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_650),
.B(n_266),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_665),
.B(n_543),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_675),
.B(n_543),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_650),
.B(n_266),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_675),
.A2(n_366),
.B1(n_334),
.B2(n_310),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_608),
.B(n_543),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_690),
.B(n_545),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_673),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_688),
.A2(n_219),
.B(n_338),
.C(n_330),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_673),
.B(n_193),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_622),
.B(n_310),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_622),
.B(n_310),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_674),
.B(n_234),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_690),
.B(n_545),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_599),
.B(n_234),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_615),
.B(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_633),
.B(n_235),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_627),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_567),
.A2(n_310),
.B1(n_195),
.B2(n_312),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_564),
.B(n_548),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_627),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_664),
.A2(n_227),
.B1(n_373),
.B2(n_370),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_637),
.Y(n_754)
);

NAND2x1p5_ASAP7_75t_L g755 ( 
.A(n_575),
.B(n_200),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_622),
.B(n_310),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_607),
.B(n_299),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_564),
.B(n_548),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_566),
.B(n_548),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_235),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_566),
.A2(n_204),
.B(n_218),
.C(n_217),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_568),
.B(n_300),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_604),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_569),
.B(n_549),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_676),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_660),
.B(n_429),
.C(n_425),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_633),
.B(n_697),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_643),
.A2(n_533),
.B(n_528),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_663),
.B(n_236),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_672),
.B(n_430),
.C(n_429),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_637),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_621),
.B(n_430),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_567),
.A2(n_353),
.B1(n_261),
.B2(n_258),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_569),
.B(n_549),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_680),
.B(n_435),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_641),
.B(n_202),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_680),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_641),
.B(n_212),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_572),
.B(n_549),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_680),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_567),
.A2(n_620),
.B(n_577),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_671),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_689),
.A2(n_304),
.B1(n_320),
.B2(n_311),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_613),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_572),
.B(n_222),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_575),
.B(n_223),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_699),
.B(n_236),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_654),
.B(n_289),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_585),
.B(n_289),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_676),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_578),
.B(n_233),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_695),
.A2(n_533),
.B(n_528),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_578),
.B(n_237),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_621),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_647),
.B(n_435),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_589),
.B(n_238),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_676),
.B(n_243),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_574),
.A2(n_704),
.B(n_620),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_589),
.B(n_592),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_639),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_609),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_583),
.B(n_443),
.C(n_440),
.Y(n_803)
);

NAND3x1_ASAP7_75t_L g804 ( 
.A(n_682),
.B(n_443),
.C(n_440),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_592),
.B(n_274),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_645),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_580),
.B(n_325),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_571),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_623),
.A2(n_382),
.B1(n_360),
.B2(n_301),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_598),
.B(n_325),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_645),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_594),
.B(n_278),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_562),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_579),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_594),
.B(n_281),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_565),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_646),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_597),
.B(n_285),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_642),
.B(n_326),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_597),
.B(n_602),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_602),
.B(n_291),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_646),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_579),
.B(n_444),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_623),
.A2(n_319),
.B1(n_318),
.B2(n_317),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_603),
.B(n_297),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_649),
.Y(n_827)
);

AND2x4_ASAP7_75t_SL g828 ( 
.A(n_611),
.B(n_444),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_603),
.B(n_528),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_606),
.B(n_528),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_649),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_606),
.B(n_528),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_618),
.B(n_528),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_533),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_623),
.B(n_448),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_629),
.B(n_533),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_611),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_655),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_629),
.B(n_533),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_642),
.B(n_326),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_613),
.B(n_316),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_642),
.B(n_328),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_631),
.B(n_533),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_562),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_631),
.B(n_328),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_655),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_611),
.B(n_448),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_632),
.B(n_535),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_605),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_632),
.B(n_535),
.Y(n_850)
);

AOI221xp5_ASAP7_75t_L g851 ( 
.A1(n_692),
.A2(n_365),
.B1(n_227),
.B2(n_339),
.C(n_345),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_667),
.B(n_412),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_656),
.B(n_535),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_561),
.B(n_262),
.C(n_263),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_570),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_702),
.B(n_329),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_656),
.B(n_535),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_659),
.B(n_535),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_570),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_659),
.Y(n_860)
);

BUFx6f_ASAP7_75t_SL g861 ( 
.A(n_670),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_662),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_571),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_577),
.B(n_329),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_577),
.A2(n_339),
.B1(n_345),
.B2(n_370),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_642),
.B(n_332),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_623),
.B(n_337),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_662),
.B(n_535),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_620),
.B(n_536),
.Y(n_869)
);

NOR2x1p5_ASAP7_75t_L g870 ( 
.A(n_666),
.B(n_365),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_707),
.B(n_536),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_586),
.B(n_450),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_612),
.B(n_536),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_612),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_614),
.B(n_340),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_614),
.B(n_340),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_616),
.B(n_341),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_683),
.B(n_687),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_616),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_601),
.B(n_341),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_576),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_617),
.B(n_536),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_666),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_719),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_816),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_725),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_783),
.B(n_617),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_874),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_791),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_879),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_720),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_L g892 ( 
.A1(n_745),
.A2(n_670),
.B(n_658),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_781),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_801),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_806),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_811),
.Y(n_896)
);

AND2x2_ASAP7_75t_SL g897 ( 
.A(n_749),
.B(n_610),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_732),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_791),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_817),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_785),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_791),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_823),
.B(n_624),
.Y(n_903)
);

BUFx4f_ASAP7_75t_L g904 ( 
.A(n_819),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_773),
.A2(n_670),
.B1(n_669),
.B2(n_648),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_827),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_831),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_773),
.A2(n_670),
.B1(n_669),
.B2(n_648),
.Y(n_908)
);

BUFx4f_ASAP7_75t_SL g909 ( 
.A(n_849),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_L g910 ( 
.A(n_723),
.B(n_586),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_838),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_732),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_726),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_791),
.B(n_624),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_846),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_723),
.B(n_625),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_860),
.B(n_625),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_878),
.B(n_630),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_862),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_878),
.B(n_782),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_744),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_SL g922 ( 
.A1(n_883),
.A2(n_565),
.B1(n_242),
.B2(n_239),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_767),
.B(n_626),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_813),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_796),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_745),
.B(n_590),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_715),
.B(n_630),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_718),
.Y(n_928)
);

CKINVDCx6p67_ASAP7_75t_R g929 ( 
.A(n_847),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_751),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_727),
.A2(n_681),
.B1(n_640),
.B2(n_703),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_721),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_735),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_851),
.B(n_865),
.C(n_724),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_800),
.B(n_634),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_737),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_742),
.B(n_657),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_821),
.B(n_634),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_865),
.B(n_259),
.C(n_245),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_777),
.A2(n_681),
.B1(n_706),
.B2(n_653),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_752),
.B(n_635),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_828),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_749),
.B(n_635),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_795),
.B(n_652),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_780),
.A2(n_681),
.B1(n_652),
.B2(n_653),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_734),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_750),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_758),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_723),
.B(n_705),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_808),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_763),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_SL g953 ( 
.A(n_789),
.B(n_264),
.C(n_260),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_736),
.B(n_705),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_717),
.A2(n_711),
.B(n_450),
.C(n_455),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_717),
.A2(n_733),
.B1(n_754),
.B2(n_748),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_759),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_814),
.B(n_342),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_764),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_765),
.B(n_628),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_847),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_723),
.B(n_710),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_774),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_779),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_824),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_819),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_771),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_819),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_810),
.A2(n_265),
.B1(n_276),
.B2(n_286),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_743),
.B(n_710),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_775),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_847),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_760),
.B(n_712),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_808),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_740),
.A2(n_712),
.B1(n_669),
.B2(n_590),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_863),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_753),
.B(n_352),
.C(n_342),
.Y(n_977)
);

CKINVDCx11_ASAP7_75t_R g978 ( 
.A(n_872),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_760),
.B(n_669),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_775),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_772),
.B(n_576),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_716),
.B(n_582),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_864),
.A2(n_713),
.B1(n_709),
.B2(n_581),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_746),
.B(n_582),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_869),
.A2(n_701),
.B(n_628),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_742),
.B(n_563),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_747),
.B(n_563),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_765),
.B(n_344),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_837),
.B(n_455),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_872),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_802),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_835),
.B(n_459),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_829),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_861),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_722),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_844),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_863),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_804),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_861),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_863),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_830),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_790),
.B(n_459),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_855),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_SL g1004 ( 
.A(n_854),
.B(n_287),
.C(n_290),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_723),
.B(n_571),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_729),
.B(n_584),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_859),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_880),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_733),
.A2(n_584),
.B1(n_593),
.B2(n_696),
.Y(n_1010)
);

NOR2x2_ASAP7_75t_L g1011 ( 
.A(n_790),
.B(n_667),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_881),
.Y(n_1012)
);

AND2x6_ASAP7_75t_L g1013 ( 
.A(n_730),
.B(n_668),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_875),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_810),
.B(n_593),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_832),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_833),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_786),
.B(n_563),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_792),
.B(n_581),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_864),
.A2(n_668),
.B1(n_708),
.B2(n_696),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_794),
.B(n_581),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_863),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_834),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_740),
.A2(n_679),
.B1(n_708),
.B2(n_693),
.Y(n_1024)
);

NOR2x2_ASAP7_75t_L g1025 ( 
.A(n_807),
.B(n_679),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_875),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_SL g1027 ( 
.A(n_741),
.B(n_344),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_836),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_766),
.B(n_464),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_741),
.A2(n_684),
.B1(n_693),
.B2(n_691),
.Y(n_1030)
);

AO21x1_ASAP7_75t_L g1031 ( 
.A1(n_756),
.A2(n_691),
.B(n_684),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_839),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_852),
.Y(n_1033)
);

AOI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_880),
.A2(n_385),
.B(n_307),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_852),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_852),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_852),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_723),
.B(n_571),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_797),
.B(n_588),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_805),
.B(n_588),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_739),
.B(n_799),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_845),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_876),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_848),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_812),
.B(n_591),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_852),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_850),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_755),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_853),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_739),
.B(n_571),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_756),
.A2(n_714),
.B1(n_807),
.B2(n_770),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_815),
.B(n_591),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_769),
.B(n_591),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_818),
.B(n_661),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_776),
.A2(n_713),
.B1(n_709),
.B2(n_661),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_822),
.B(n_826),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_755),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_787),
.B(n_661),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_857),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_787),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_858),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_868),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_809),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_873),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_845),
.B(n_685),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_788),
.B(n_685),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_856),
.A2(n_470),
.B1(n_475),
.B2(n_473),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_876),
.B(n_877),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_778),
.B(n_798),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_889),
.Y(n_1072)
);

AOI33xp33_ASAP7_75t_L g1073 ( 
.A1(n_967),
.A2(n_470),
.A3(n_478),
.B1(n_473),
.B2(n_471),
.B3(n_464),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_934),
.A2(n_877),
.B(n_738),
.C(n_798),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_886),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_889),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_SL g1077 ( 
.A1(n_1031),
.A2(n_768),
.B(n_871),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_901),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_889),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_885),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1009),
.B(n_820),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_937),
.B(n_841),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_932),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_SL g1084 ( 
.A1(n_1034),
.A2(n_731),
.B(n_728),
.C(n_478),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_893),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1002),
.B(n_947),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_924),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_901),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_937),
.B(n_925),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_916),
.A2(n_701),
.B(n_628),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_966),
.B(n_867),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_948),
.B(n_867),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_940),
.A2(n_803),
.B(n_762),
.C(n_761),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_899),
.B(n_701),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1042),
.A2(n_793),
.B(n_757),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_889),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_897),
.A2(n_842),
.B1(n_840),
.B2(n_820),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_966),
.B(n_825),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_928),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_924),
.Y(n_1100)
);

BUFx12f_ASAP7_75t_L g1101 ( 
.A(n_978),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_926),
.B(n_923),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_968),
.B(n_866),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_909),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_920),
.A2(n_866),
.B(n_842),
.C(n_840),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_894),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_994),
.B(n_308),
.C(n_314),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_909),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_923),
.A2(n_784),
.B1(n_346),
.B2(n_367),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_925),
.B(n_315),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_892),
.A2(n_698),
.B(n_381),
.C(n_379),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_897),
.A2(n_346),
.B1(n_379),
.B2(n_352),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_995),
.A2(n_355),
.B1(n_378),
.B2(n_367),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_902),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_884),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_SL g1116 ( 
.A(n_977),
.B(n_375),
.C(n_369),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_899),
.B(n_355),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_895),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_956),
.A2(n_469),
.B1(n_471),
.B2(n_475),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_968),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_949),
.B(n_698),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_888),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_965),
.B(n_369),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_902),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1042),
.A2(n_636),
.B(n_596),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_378),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_899),
.B(n_596),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_922),
.B(n_969),
.C(n_998),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_996),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_974),
.A2(n_636),
.B(n_596),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_974),
.A2(n_636),
.B(n_596),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1043),
.B(n_596),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1003),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1043),
.A2(n_469),
.B(n_452),
.C(n_412),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_636),
.B(n_686),
.Y(n_1135)
);

AOI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1068),
.A2(n_959),
.B1(n_963),
.B2(n_957),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_899),
.B(n_636),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1005),
.A2(n_412),
.B(n_437),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_989),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1026),
.B(n_700),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1008),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1007),
.Y(n_1142)
);

OR2x6_ASAP7_75t_SL g1143 ( 
.A(n_999),
.B(n_417),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_896),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_961),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_902),
.B(n_418),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_964),
.B(n_452),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_974),
.A2(n_686),
.B(n_587),
.Y(n_1148)
);

NOR2xp67_ASAP7_75t_L g1149 ( 
.A(n_943),
.B(n_82),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1014),
.B(n_1044),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1064),
.A2(n_418),
.B(n_419),
.C(n_465),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1064),
.A2(n_419),
.B(n_468),
.C(n_465),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1052),
.A2(n_468),
.B(n_437),
.C(n_457),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_900),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_902),
.B(n_465),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_887),
.A2(n_686),
.B(n_587),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1061),
.B(n_481),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_992),
.B(n_1061),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_956),
.A2(n_481),
.B1(n_468),
.B2(n_457),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_938),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_906),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1071),
.A2(n_481),
.B(n_457),
.C(n_437),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1052),
.A2(n_436),
.B1(n_686),
.B2(n_587),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1069),
.A2(n_436),
.B(n_554),
.C(n_536),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1071),
.A2(n_436),
.B(n_554),
.C(n_536),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_SL g1166 ( 
.A1(n_990),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_933),
.B(n_4),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_R g1168 ( 
.A(n_978),
.B(n_191),
.Y(n_1168)
);

INVx8_ASAP7_75t_L g1169 ( 
.A(n_989),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_938),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_931),
.B(n_700),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_904),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_992),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_987),
.A2(n_554),
.B(n_587),
.C(n_9),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_907),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_977),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.C(n_13),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_971),
.A2(n_980),
.B1(n_987),
.B2(n_992),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_989),
.Y(n_1178)
);

NOR3xp33_ASAP7_75t_L g1179 ( 
.A(n_1049),
.B(n_5),
.C(n_10),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_979),
.A2(n_1049),
.B1(n_1058),
.B2(n_1057),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_935),
.B(n_700),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1029),
.B(n_13),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1038),
.A2(n_554),
.B(n_189),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_938),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1012),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_891),
.Y(n_1186)
);

NAND2xp33_ASAP7_75t_R g1187 ( 
.A(n_953),
.B(n_174),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_929),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_913),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_1027),
.A2(n_165),
.B(n_148),
.C(n_145),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_939),
.B(n_554),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_942),
.B(n_15),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1038),
.A2(n_985),
.B(n_944),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_927),
.A2(n_554),
.B(n_140),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_905),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_921),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1058),
.B(n_138),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_R g1198 ( 
.A(n_904),
.B(n_120),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_936),
.B(n_112),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_936),
.B(n_16),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1066),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_911),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_918),
.A2(n_21),
.B(n_23),
.C(n_25),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_915),
.B(n_919),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_918),
.A2(n_25),
.B(n_27),
.C(n_30),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_984),
.A2(n_102),
.B(n_101),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1029),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_972),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_982),
.A2(n_99),
.B(n_91),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_898),
.A2(n_66),
.B(n_37),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_993),
.B(n_35),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_SL g1212 ( 
.A1(n_905),
.A2(n_38),
.B(n_40),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_954),
.A2(n_970),
.B(n_1006),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_973),
.B(n_981),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_945),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_930),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_898),
.A2(n_38),
.B(n_42),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_986),
.B(n_46),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_912),
.A2(n_66),
.B(n_50),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_975),
.A2(n_47),
.B(n_53),
.C(n_55),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_903),
.A2(n_47),
.B(n_55),
.C(n_56),
.Y(n_1221)
);

AO32x2_ASAP7_75t_L g1222 ( 
.A1(n_1047),
.A2(n_56),
.A3(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1066),
.A2(n_986),
.B(n_1054),
.C(n_946),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_972),
.B(n_62),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_938),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_950),
.A2(n_65),
.B(n_962),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1051),
.A2(n_65),
.B(n_1015),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_917),
.A2(n_1004),
.B(n_890),
.C(n_955),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_908),
.A2(n_1068),
.B1(n_1022),
.B2(n_1010),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1020),
.A2(n_1024),
.B(n_1030),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_951),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1001),
.B(n_1017),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1023),
.B(n_1028),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1089),
.B(n_1041),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1086),
.B(n_1045),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1095),
.A2(n_914),
.B(n_1051),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1125),
.A2(n_914),
.B(n_1020),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1138),
.A2(n_1024),
.B(n_1030),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1193),
.A2(n_1039),
.B(n_1019),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1231),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1097),
.A2(n_908),
.B1(n_1022),
.B2(n_941),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1214),
.B(n_1092),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1081),
.B(n_958),
.Y(n_1243)
);

AOI211x1_ASAP7_75t_L g1244 ( 
.A1(n_1195),
.A2(n_1067),
.B(n_991),
.C(n_1062),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1223),
.A2(n_1054),
.A3(n_1063),
.B(n_1021),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1092),
.B(n_958),
.Y(n_1246)
);

INVx3_ASAP7_75t_SL g1247 ( 
.A(n_1099),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1158),
.B(n_1004),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1077),
.A2(n_960),
.B(n_1070),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1078),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1104),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1136),
.A2(n_1040),
.B(n_1055),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1213),
.A2(n_1018),
.B(n_1046),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_SL g1254 ( 
.A1(n_1228),
.A2(n_1059),
.B(n_1047),
.Y(n_1254)
);

AO21x1_ASAP7_75t_L g1255 ( 
.A1(n_1218),
.A2(n_910),
.B(n_1053),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1075),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1213),
.A2(n_1016),
.B(n_1032),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1080),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1182),
.B(n_1207),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1083),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1215),
.B(n_953),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1090),
.A2(n_983),
.B(n_1065),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1181),
.A2(n_1060),
.B(n_1050),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1229),
.A2(n_1048),
.A3(n_955),
.B(n_952),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1181),
.A2(n_951),
.B(n_976),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1085),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1227),
.A2(n_997),
.B(n_1056),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1106),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1195),
.A2(n_1176),
.B1(n_1068),
.B2(n_1116),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1102),
.B(n_988),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1180),
.A2(n_1233),
.B1(n_1232),
.B2(n_1177),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1231),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1087),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1088),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1105),
.A2(n_951),
.B(n_976),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1230),
.A2(n_951),
.B(n_976),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1128),
.A2(n_1037),
.B1(n_1036),
.B2(n_1035),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1191),
.A2(n_1013),
.B(n_1037),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1100),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1110),
.B(n_988),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1150),
.B(n_1204),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1226),
.A2(n_1013),
.B(n_997),
.Y(n_1282)
);

INVx3_ASAP7_75t_SL g1283 ( 
.A(n_1141),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1230),
.A2(n_976),
.B(n_1000),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1082),
.B(n_1000),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1229),
.A2(n_1013),
.A3(n_1025),
.B(n_1011),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1204),
.B(n_1013),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1118),
.B(n_1013),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1144),
.B(n_1000),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1191),
.A2(n_1033),
.B(n_1035),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1192),
.B(n_1000),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1115),
.B(n_1033),
.Y(n_1292)
);

AOI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1171),
.A2(n_1156),
.B(n_1163),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1074),
.A2(n_1033),
.B(n_1035),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1169),
.B(n_1091),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1130),
.A2(n_1033),
.B(n_1035),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1154),
.B(n_1036),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1147),
.A2(n_1036),
.B(n_1037),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1164),
.A2(n_1036),
.B(n_1037),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1131),
.A2(n_1183),
.B(n_1084),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1231),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1111),
.A2(n_1157),
.B(n_1093),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_1153),
.B(n_1163),
.Y(n_1303)
);

NOR4xp25_ASAP7_75t_L g1304 ( 
.A(n_1220),
.B(n_1208),
.C(n_1201),
.D(n_1221),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1123),
.B(n_1126),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_R g1306 ( 
.A(n_1188),
.B(n_1108),
.Y(n_1306)
);

AO21x1_ASAP7_75t_L g1307 ( 
.A1(n_1203),
.A2(n_1205),
.B(n_1211),
.Y(n_1307)
);

AO32x2_ASAP7_75t_L g1308 ( 
.A1(n_1119),
.A2(n_1159),
.A3(n_1166),
.B1(n_1222),
.B2(n_1139),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1161),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1211),
.A2(n_1132),
.B(n_1174),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1175),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1155),
.A2(n_1159),
.B(n_1094),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1202),
.B(n_1122),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1231),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1109),
.A2(n_1200),
.B(n_1212),
.C(n_1167),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1179),
.A2(n_1194),
.B1(n_1210),
.B2(n_1219),
.C(n_1217),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1121),
.A2(n_1135),
.B(n_1148),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1076),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1119),
.A2(n_1224),
.B1(n_1112),
.B2(n_1151),
.C(n_1098),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1129),
.B(n_1185),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1165),
.A2(n_1134),
.B(n_1121),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1133),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1094),
.A2(n_1206),
.B(n_1209),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1146),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1142),
.B(n_1186),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1152),
.A2(n_1196),
.B(n_1216),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1091),
.A2(n_1103),
.B1(n_1098),
.B2(n_1189),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1145),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1155),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1073),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1140),
.B(n_1091),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1113),
.B(n_1103),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1155),
.A2(n_1199),
.B(n_1146),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1076),
.Y(n_1334)
);

AOI221x1_ASAP7_75t_L g1335 ( 
.A1(n_1222),
.A2(n_1072),
.B1(n_1079),
.B2(n_1124),
.C(n_1190),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1146),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1127),
.A2(n_1137),
.B(n_1162),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1178),
.B(n_1173),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1120),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1096),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1072),
.A2(n_1079),
.B(n_1124),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1197),
.A2(n_1117),
.B(n_1103),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1343)
);

AOI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1149),
.A2(n_1187),
.B(n_1170),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1101),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1107),
.A2(n_1168),
.B(n_1198),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1169),
.B(n_1096),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1170),
.A2(n_1184),
.B(n_1114),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1184),
.A2(n_1114),
.B(n_1076),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1160),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1160),
.A2(n_1225),
.B(n_1222),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1160),
.A2(n_1225),
.B(n_1143),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1225),
.B(n_1089),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1075),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1223),
.A2(n_920),
.B(n_1092),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1081),
.B(n_1009),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1075),
.Y(n_1360)
);

CKINVDCx14_ASAP7_75t_R g1361 ( 
.A(n_1099),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1195),
.A2(n_934),
.B1(n_897),
.B2(n_1097),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1218),
.A2(n_977),
.B1(n_892),
.B2(n_1227),
.C(n_1229),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1075),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1075),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1223),
.A2(n_920),
.B(n_791),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1223),
.A2(n_1229),
.A3(n_1031),
.B(n_1164),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1077),
.A2(n_1095),
.B(n_1223),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1097),
.A2(n_654),
.B(n_682),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1223),
.A2(n_934),
.B(n_920),
.C(n_1197),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1092),
.B(n_925),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1074),
.A2(n_937),
.B(n_892),
.C(n_878),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1087),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1092),
.B(n_1214),
.Y(n_1380)
);

NAND2x1_ASAP7_75t_L g1381 ( 
.A(n_1096),
.B(n_889),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1172),
.B(n_966),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1097),
.A2(n_654),
.B(n_682),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1077),
.A2(n_1095),
.B(n_1223),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1125),
.A2(n_1138),
.B(n_1095),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1158),
.B(n_925),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_L g1388 ( 
.A(n_1082),
.B(n_937),
.C(n_934),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1389)
);

OAI22x1_ASAP7_75t_L g1390 ( 
.A1(n_1177),
.A2(n_1009),
.B1(n_937),
.B2(n_1081),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1077),
.A2(n_1095),
.B(n_1223),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1099),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1223),
.A2(n_920),
.B(n_1092),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1125),
.A2(n_1138),
.B(n_1095),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1089),
.B(n_1086),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_920),
.Y(n_1398)
);

NOR2x1_ASAP7_75t_SL g1399 ( 
.A(n_1271),
.B(n_1240),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1361),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1293),
.A2(n_1275),
.B(n_1236),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1295),
.B(n_1329),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1286),
.B(n_1362),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1240),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1305),
.A2(n_1362),
.B1(n_1242),
.B2(n_1395),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1250),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1273),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1278),
.A2(n_1262),
.B(n_1371),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1354),
.A2(n_1389),
.B(n_1376),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1256),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1266),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1334),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1305),
.A2(n_1378),
.B(n_1315),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1274),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1268),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1373),
.A2(n_1383),
.B1(n_1390),
.B2(n_1396),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1311),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1354),
.A2(n_1389),
.B(n_1376),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1397),
.A2(n_1398),
.B(n_1323),
.Y(n_1421)
);

XOR2xp5_ASAP7_75t_L g1422 ( 
.A(n_1258),
.B(n_1327),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1249),
.A2(n_1284),
.B(n_1276),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1276),
.A2(n_1284),
.B(n_1237),
.Y(n_1424)
);

AO21x1_ASAP7_75t_L g1425 ( 
.A1(n_1388),
.A2(n_1310),
.B(n_1302),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1251),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1388),
.A2(n_1319),
.B1(n_1269),
.B2(n_1270),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1328),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1279),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_R g1430 ( 
.A(n_1345),
.B(n_1382),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1379),
.Y(n_1431)
);

BUFx2_ASAP7_75t_SL g1432 ( 
.A(n_1339),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1319),
.A2(n_1269),
.B1(n_1270),
.B2(n_1261),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1355),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1363),
.A2(n_1393),
.B(n_1356),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1281),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1360),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1248),
.A2(n_1246),
.B1(n_1280),
.B2(n_1330),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1300),
.A2(n_1239),
.B(n_1275),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1364),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1365),
.B(n_1369),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1366),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1307),
.A2(n_1243),
.B1(n_1358),
.B2(n_1332),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1370),
.B(n_1375),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1298),
.A2(n_1265),
.B(n_1303),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_SL g1446 ( 
.A1(n_1285),
.A2(n_1380),
.B(n_1294),
.C(n_1288),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1313),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1335),
.A2(n_1255),
.B(n_1303),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1334),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1264),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1260),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1264),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1320),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1387),
.B(n_1377),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1290),
.A2(n_1282),
.B(n_1253),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1367),
.A2(n_1253),
.B(n_1312),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1234),
.A2(n_1235),
.B1(n_1336),
.B2(n_1277),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1380),
.B(n_1304),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1374),
.A2(n_1257),
.B(n_1263),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1254),
.A2(n_1238),
.B(n_1257),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1263),
.A2(n_1316),
.B(n_1285),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1259),
.A2(n_1241),
.B1(n_1386),
.B2(n_1346),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1296),
.A2(n_1351),
.B(n_1337),
.Y(n_1463)
);

AO32x2_ASAP7_75t_L g1464 ( 
.A1(n_1308),
.A2(n_1286),
.A3(n_1245),
.B1(n_1368),
.B2(n_1391),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1291),
.A2(n_1331),
.B1(n_1324),
.B2(n_1287),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1325),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1240),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1322),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1289),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

AOI22x1_ASAP7_75t_L g1471 ( 
.A1(n_1337),
.A2(n_1326),
.B1(n_1352),
.B2(n_1324),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1342),
.A2(n_1252),
.B(n_1267),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1382),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1299),
.A2(n_1252),
.B(n_1321),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1299),
.A2(n_1321),
.B(n_1341),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1297),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1372),
.A2(n_1391),
.B(n_1384),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1245),
.B(n_1286),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1286),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1308),
.B(n_1245),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1336),
.A2(n_1295),
.B1(n_1338),
.B2(n_1247),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1245),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1348),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1333),
.A2(n_1352),
.B(n_1381),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_SL g1485 ( 
.A1(n_1347),
.A2(n_1301),
.B(n_1350),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1368),
.A2(n_1292),
.B(n_1318),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1283),
.A2(n_1343),
.B1(n_1244),
.B2(n_1318),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1340),
.A2(n_1301),
.B(n_1334),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1308),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1308),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1340),
.B(n_1334),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1368),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1240),
.A2(n_1272),
.B(n_1314),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1272),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1306),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1272),
.A2(n_1314),
.B(n_1368),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1314),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1251),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1392),
.A2(n_1305),
.B1(n_934),
.B2(n_1362),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1392),
.A2(n_1306),
.B(n_1283),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1260),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1502)
);

INVxp33_ASAP7_75t_L g1503 ( 
.A(n_1386),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1305),
.A2(n_1009),
.B1(n_1097),
.B2(n_1362),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_L g1506 ( 
.A1(n_1305),
.A2(n_937),
.B(n_1009),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1309),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1305),
.B(n_1009),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1309),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1309),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1295),
.B(n_1329),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1309),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1260),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1260),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1309),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1309),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1305),
.B(n_1271),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1361),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1286),
.B(n_1362),
.Y(n_1523)
);

AO22x2_ASAP7_75t_L g1524 ( 
.A1(n_1363),
.A2(n_1335),
.B1(n_1195),
.B2(n_1388),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1335),
.A2(n_1255),
.A3(n_1363),
.B(n_1354),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1305),
.A2(n_937),
.B(n_1378),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1240),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1335),
.A2(n_1376),
.B(n_1354),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1286),
.B(n_1362),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1245),
.B(n_1286),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1309),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1250),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1258),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1354),
.A2(n_1389),
.B(n_1376),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1305),
.A2(n_934),
.B1(n_1362),
.B2(n_937),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1309),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1309),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1305),
.B(n_1009),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1309),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1305),
.A2(n_937),
.B1(n_1009),
.B2(n_1362),
.C(n_934),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1385),
.A2(n_1394),
.B(n_1317),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1240),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1334),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1309),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1240),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1260),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1309),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1309),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_1454),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1444),
.B(n_1436),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1503),
.B(n_1470),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1462),
.B(n_1438),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1417),
.B(n_1441),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1483),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1504),
.B(n_1507),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1483),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1456),
.A2(n_1521),
.B(n_1526),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1403),
.B(n_1512),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1521),
.A2(n_1505),
.B(n_1506),
.C(n_1414),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1541),
.A2(n_1418),
.B(n_1536),
.C(n_1406),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1447),
.B(n_1499),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1453),
.B(n_1466),
.Y(n_1563)
);

NOR2xp67_ASAP7_75t_L g1564 ( 
.A(n_1495),
.B(n_1534),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1509),
.A2(n_1539),
.B1(n_1433),
.B2(n_1427),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_1425),
.A2(n_1458),
.B(n_1435),
.C(n_1461),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1434),
.Y(n_1567)
);

AOI221x1_ASAP7_75t_SL g1568 ( 
.A1(n_1457),
.A2(n_1440),
.B1(n_1419),
.B2(n_1416),
.C(n_1412),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1465),
.B(n_1443),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1451),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1422),
.A2(n_1481),
.B1(n_1487),
.B2(n_1495),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1439),
.A2(n_1477),
.B(n_1474),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1403),
.B(n_1512),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1403),
.B(n_1512),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1437),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1458),
.B(n_1517),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1469),
.B(n_1476),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1459),
.A2(n_1425),
.B(n_1496),
.C(n_1523),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1399),
.A2(n_1430),
.B(n_1491),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1422),
.A2(n_1400),
.B1(n_1522),
.B2(n_1524),
.Y(n_1581)
);

O2A1O1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1446),
.A2(n_1501),
.B(n_1516),
.C(n_1547),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1404),
.A2(n_1523),
.B(n_1530),
.C(n_1410),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1404),
.A2(n_1530),
.B(n_1410),
.C(n_1420),
.Y(n_1584)
);

O2A1O1Ixp5_ASAP7_75t_L g1585 ( 
.A1(n_1472),
.A2(n_1482),
.B(n_1402),
.C(n_1492),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1468),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1524),
.A2(n_1415),
.B1(n_1428),
.B2(n_1473),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1508),
.B(n_1510),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1439),
.A2(n_1474),
.B(n_1424),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1473),
.B(n_1511),
.Y(n_1590)
);

O2A1O1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1446),
.A2(n_1485),
.B(n_1442),
.C(n_1411),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1432),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1513),
.B(n_1519),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1407),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1424),
.A2(n_1423),
.B(n_1445),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1407),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1426),
.Y(n_1597)
);

O2A1O1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1485),
.A2(n_1498),
.B(n_1548),
.C(n_1545),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1492),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1524),
.A2(n_1471),
.B1(n_1533),
.B2(n_1522),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1520),
.B(n_1532),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1533),
.A2(n_1400),
.B1(n_1426),
.B2(n_1549),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1537),
.B(n_1540),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1408),
.B(n_1431),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1429),
.B(n_1431),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1478),
.B(n_1531),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1478),
.B(n_1531),
.Y(n_1607)
);

OA21x2_ASAP7_75t_L g1608 ( 
.A1(n_1423),
.A2(n_1445),
.B(n_1421),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1497),
.B(n_1494),
.Y(n_1609)
);

NAND2x1_ASAP7_75t_L g1610 ( 
.A(n_1488),
.B(n_1486),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1484),
.A2(n_1455),
.B(n_1479),
.C(n_1480),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1484),
.B(n_1467),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1455),
.A2(n_1479),
.B(n_1480),
.C(n_1450),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1543),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1491),
.A2(n_1486),
.B(n_1544),
.Y(n_1615)
);

A2O1A1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1450),
.A2(n_1452),
.B(n_1500),
.C(n_1493),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1525),
.B(n_1452),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1528),
.B(n_1500),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1528),
.B(n_1546),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1486),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1543),
.A2(n_1544),
.B1(n_1413),
.B2(n_1449),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1413),
.A2(n_1449),
.B(n_1448),
.C(n_1535),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1464),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1535),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1460),
.B(n_1463),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1405),
.B(n_1475),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1401),
.A2(n_1514),
.B(n_1542),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1525),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1463),
.A2(n_1489),
.B(n_1490),
.C(n_1525),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1543),
.B(n_1464),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1448),
.A2(n_1529),
.B1(n_1472),
.B2(n_1525),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1525),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1401),
.A2(n_1502),
.B(n_1515),
.Y(n_1633)
);

BUFx4_ASAP7_75t_R g1634 ( 
.A(n_1464),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1409),
.A2(n_1515),
.B(n_1518),
.C(n_1527),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1518),
.A2(n_1305),
.B(n_1526),
.C(n_1521),
.Y(n_1636)
);

OAI22x1_ASAP7_75t_L g1637 ( 
.A1(n_1521),
.A2(n_1009),
.B1(n_1305),
.B2(n_1458),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1444),
.B(n_1454),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1536),
.A2(n_1009),
.B1(n_1539),
.B2(n_1509),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1434),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1536),
.A2(n_1009),
.B1(n_1539),
.B2(n_1509),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1526),
.A2(n_1305),
.B(n_1521),
.C(n_937),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1526),
.A2(n_1305),
.B(n_1521),
.C(n_937),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1444),
.B(n_1454),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1526),
.A2(n_1305),
.B(n_1521),
.C(n_937),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1407),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1526),
.B(n_1521),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1536),
.A2(n_1009),
.B1(n_1539),
.B2(n_1509),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1434),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1536),
.A2(n_1009),
.B1(n_1539),
.B2(n_1509),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1414),
.A2(n_1526),
.B(n_1305),
.C(n_1541),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1503),
.B(n_1386),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1439),
.A2(n_1477),
.B(n_1335),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1503),
.B(n_1386),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1583),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1597),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1583),
.B(n_1584),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1599),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1642),
.A2(n_1645),
.B(n_1643),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1635),
.A2(n_1631),
.B(n_1558),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1566),
.A2(n_1585),
.B(n_1579),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1612),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1618),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1615),
.B(n_1579),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1612),
.B(n_1626),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1644),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1584),
.B(n_1550),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1613),
.A2(n_1620),
.B(n_1611),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1606),
.B(n_1607),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1617),
.B(n_1629),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1554),
.B(n_1556),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1577),
.Y(n_1673)
);

NAND2x1_ASAP7_75t_L g1674 ( 
.A(n_1615),
.B(n_1580),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1654),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1611),
.B(n_1629),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1651),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1570),
.Y(n_1679)
);

AO21x2_ASAP7_75t_L g1680 ( 
.A1(n_1624),
.A2(n_1616),
.B(n_1622),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1647),
.B(n_1651),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1559),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1590),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_L g1684 ( 
.A(n_1572),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1626),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1610),
.B(n_1625),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1616),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_L g1688 ( 
.A(n_1561),
.B(n_1565),
.C(n_1560),
.D(n_1648),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1567),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1636),
.A2(n_1650),
.B(n_1641),
.Y(n_1690)
);

OR2x6_ASAP7_75t_L g1691 ( 
.A(n_1625),
.B(n_1591),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1576),
.B(n_1640),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1649),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1646),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1609),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1628),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1571),
.B(n_1594),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1632),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1587),
.B(n_1623),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1559),
.B(n_1574),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1555),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1555),
.A2(n_1557),
.B(n_1627),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1589),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1625),
.B(n_1555),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1557),
.A2(n_1627),
.B(n_1633),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1604),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1605),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1690),
.A2(n_1581),
.B(n_1600),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1669),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1568),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1662),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1562),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1582),
.B(n_1569),
.C(n_1553),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1705),
.Y(n_1716)
);

OAI222xp33_ASAP7_75t_L g1717 ( 
.A1(n_1678),
.A2(n_1578),
.B1(n_1563),
.B2(n_1598),
.C1(n_1634),
.C2(n_1574),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1670),
.B(n_1653),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1705),
.Y(n_1719)
);

BUFx4f_ASAP7_75t_L g1720 ( 
.A(n_1664),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1656),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1670),
.B(n_1573),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1657),
.B(n_1573),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1706),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1707),
.A2(n_1704),
.B(n_1687),
.Y(n_1727)
);

AOI322xp5_ASAP7_75t_L g1728 ( 
.A1(n_1681),
.A2(n_1597),
.A3(n_1634),
.B1(n_1572),
.B2(n_1596),
.C1(n_1592),
.C2(n_1637),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1665),
.B(n_1589),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1698),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1665),
.B(n_1589),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1673),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1677),
.B(n_1595),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1689),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1689),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1677),
.B(n_1595),
.Y(n_1736)
);

OR2x6_ASAP7_75t_L g1737 ( 
.A(n_1664),
.B(n_1608),
.Y(n_1737)
);

AOI33xp33_ASAP7_75t_L g1738 ( 
.A1(n_1688),
.A2(n_1708),
.A3(n_1709),
.B1(n_1603),
.B2(n_1593),
.B3(n_1695),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1658),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1658),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1698),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1586),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1734),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1710),
.A2(n_1659),
.B1(n_1693),
.B2(n_1699),
.C(n_1687),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1710),
.A2(n_1666),
.B1(n_1664),
.B2(n_1661),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1734),
.Y(n_1746)
);

AOI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1715),
.A2(n_1717),
.B1(n_1712),
.B2(n_1672),
.C1(n_1720),
.C2(n_1679),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1735),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1711),
.B(n_1702),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1715),
.A2(n_1664),
.B1(n_1702),
.B2(n_1674),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1714),
.B(n_1671),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1712),
.A2(n_1664),
.B1(n_1674),
.B2(n_1691),
.Y(n_1752)
);

OR2x6_ASAP7_75t_SL g1753 ( 
.A(n_1714),
.B(n_1718),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1702),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1720),
.A2(n_1661),
.B1(n_1684),
.B2(n_1676),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1732),
.B(n_1742),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1720),
.A2(n_1691),
.B1(n_1682),
.B2(n_1661),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1716),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1663),
.Y(n_1759)
);

NOR4xp25_ASAP7_75t_L g1760 ( 
.A(n_1738),
.B(n_1683),
.C(n_1588),
.D(n_1601),
.Y(n_1760)
);

NOR4xp25_ASAP7_75t_SL g1761 ( 
.A(n_1726),
.B(n_1703),
.C(n_1675),
.D(n_1700),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1720),
.A2(n_1661),
.B1(n_1684),
.B2(n_1660),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1720),
.A2(n_1684),
.B1(n_1660),
.B2(n_1575),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1723),
.A2(n_1660),
.B1(n_1680),
.B2(n_1691),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1721),
.A2(n_1680),
.B1(n_1691),
.B2(n_1701),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_R g1766 ( 
.A(n_1726),
.B(n_1696),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1735),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1730),
.Y(n_1768)
);

OAI211xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1728),
.A2(n_1697),
.B(n_1709),
.C(n_1663),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1726),
.A2(n_1682),
.B1(n_1696),
.B2(n_1701),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1742),
.B(n_1696),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1725),
.A2(n_1721),
.B1(n_1722),
.B2(n_1733),
.C(n_1736),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1716),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1728),
.A2(n_1686),
.B1(n_1564),
.B2(n_1692),
.C(n_1685),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1713),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1738),
.B(n_1686),
.C(n_1668),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1722),
.B(n_1694),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1741),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1722),
.B(n_1685),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1718),
.B(n_1686),
.C(n_1668),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1713),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1737),
.A2(n_1614),
.B1(n_1621),
.B2(n_1619),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1718),
.B(n_1739),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1713),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1758),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_SL g1788 ( 
.A(n_1744),
.B(n_1724),
.C(n_1725),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1782),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1766),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1768),
.B(n_1771),
.Y(n_1791)
);

INVx4_ASAP7_75t_SL g1792 ( 
.A(n_1782),
.Y(n_1792)
);

OAI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1747),
.A2(n_1724),
.B(n_1725),
.Y(n_1793)
);

CKINVDCx14_ASAP7_75t_R g1794 ( 
.A(n_1766),
.Y(n_1794)
);

OR2x6_ASAP7_75t_L g1795 ( 
.A(n_1777),
.B(n_1737),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1779),
.B(n_1739),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1753),
.B(n_1729),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1784),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1745),
.A2(n_1737),
.B(n_1668),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

INVx4_ASAP7_75t_SL g1802 ( 
.A(n_1776),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

BUFx8_ASAP7_75t_L g1804 ( 
.A(n_1785),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1767),
.Y(n_1805)
);

OA21x2_ASAP7_75t_L g1806 ( 
.A1(n_1781),
.A2(n_1764),
.B(n_1765),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1764),
.A2(n_1727),
.B(n_1719),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1759),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1774),
.B(n_1724),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1780),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1778),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1756),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1749),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1760),
.B(n_1719),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1754),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1770),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1772),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1751),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1786),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1786),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1801),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1797),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1790),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1797),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1790),
.B(n_1773),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1814),
.B(n_1765),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1794),
.B(n_1731),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1814),
.B(n_1740),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1803),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1812),
.B(n_1772),
.Y(n_1830)
);

NOR2x1_ASAP7_75t_SL g1831 ( 
.A(n_1795),
.B(n_1737),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1794),
.B(n_1731),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1798),
.B(n_1731),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1793),
.A2(n_1745),
.B1(n_1769),
.B2(n_1775),
.Y(n_1834)
);

NOR2xp67_ASAP7_75t_L g1835 ( 
.A(n_1788),
.B(n_1762),
.Y(n_1835)
);

OR2x6_ASAP7_75t_L g1836 ( 
.A(n_1800),
.B(n_1783),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1801),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1803),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1805),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1788),
.B(n_1762),
.C(n_1755),
.D(n_1763),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_R g1842 ( 
.A(n_1804),
.B(n_1816),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1805),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1793),
.B(n_1752),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1805),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1799),
.B(n_1811),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1787),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1791),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1791),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1806),
.B(n_1755),
.C(n_1763),
.Y(n_1850)
);

INVxp33_ASAP7_75t_L g1851 ( 
.A(n_1842),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1819),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1823),
.B(n_1834),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1818),
.B(n_1796),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1823),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_SL g1856 ( 
.A(n_1844),
.B(n_1800),
.C(n_1761),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1819),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1820),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1835),
.A2(n_1750),
.B(n_1816),
.C(n_1807),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1820),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1822),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1835),
.A2(n_1806),
.B1(n_1795),
.B2(n_1757),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1823),
.B(n_1817),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1792),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1818),
.B(n_1809),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1841),
.A2(n_1806),
.B1(n_1795),
.B2(n_1817),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1822),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1830),
.B(n_1813),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1827),
.B(n_1792),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1825),
.B(n_1813),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1826),
.B(n_1813),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1824),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1832),
.B(n_1792),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1825),
.B(n_1815),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1843),
.B(n_1815),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1846),
.B(n_1809),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1832),
.B(n_1792),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1843),
.B(n_1815),
.Y(n_1878)
);

AND2x4_ASAP7_75t_SL g1879 ( 
.A(n_1839),
.B(n_1808),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1821),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1845),
.B(n_1802),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1826),
.B(n_1810),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1831),
.B(n_1792),
.Y(n_1883)
);

OAI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1841),
.A2(n_1850),
.B1(n_1836),
.B2(n_1795),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1821),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1821),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1824),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1852),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1857),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1879),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1879),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1858),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1855),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1860),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1882),
.B(n_1846),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1864),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1870),
.B(n_1874),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1855),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1871),
.B(n_1828),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1854),
.B(n_1828),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1864),
.B(n_1831),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1869),
.B(n_1829),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1869),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1881),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1853),
.B(n_1845),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1906)
);

AND2x4_ASAP7_75t_SL g1907 ( 
.A(n_1881),
.B(n_1789),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1881),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1861),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1877),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1877),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1876),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1876),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1911),
.B(n_1851),
.Y(n_1915)
);

AOI21xp33_ASAP7_75t_L g1916 ( 
.A1(n_1896),
.A2(n_1851),
.B(n_1884),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1913),
.Y(n_1917)
);

XOR2xp5_ASAP7_75t_L g1918 ( 
.A(n_1905),
.B(n_1856),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1911),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1912),
.B(n_1866),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1913),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1913),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1898),
.B(n_1875),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1890),
.B(n_1878),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1890),
.Y(n_1927)
);

A2O1A1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1897),
.A2(n_1850),
.B(n_1859),
.C(n_1862),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1906),
.A2(n_1859),
.B(n_1836),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1904),
.B(n_1868),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1906),
.B(n_1883),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1908),
.B(n_1883),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1904),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1914),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1928),
.B(n_1901),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1919),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1918),
.A2(n_1897),
.B1(n_1836),
.B2(n_1891),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1927),
.B(n_1902),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1915),
.B(n_1891),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_1908),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1933),
.B(n_1902),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1916),
.B(n_1909),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1920),
.B(n_1909),
.Y(n_1943)
);

OAI21xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1918),
.A2(n_1901),
.B(n_1895),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1917),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1935),
.A2(n_1928),
.B1(n_1929),
.B2(n_1921),
.C(n_1925),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1944),
.B(n_1923),
.C(n_1922),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_SL g1948 ( 
.A(n_1937),
.B(n_1930),
.C(n_1926),
.Y(n_1948)
);

NAND3xp33_ASAP7_75t_SL g1949 ( 
.A(n_1937),
.B(n_1942),
.C(n_1938),
.Y(n_1949)
);

NOR2x1p5_ASAP7_75t_SL g1950 ( 
.A(n_1936),
.B(n_1917),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1939),
.A2(n_1932),
.B(n_1931),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1940),
.B(n_1934),
.Y(n_1952)
);

AOI211xp5_ASAP7_75t_L g1953 ( 
.A1(n_1943),
.A2(n_1924),
.B(n_1932),
.C(n_1893),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1945),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1946),
.A2(n_1941),
.B(n_1893),
.C(n_1909),
.Y(n_1955)
);

AOI322xp5_ASAP7_75t_L g1956 ( 
.A1(n_1949),
.A2(n_1892),
.A3(n_1910),
.B1(n_1888),
.B2(n_1889),
.C1(n_1894),
.C2(n_1914),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1951),
.A2(n_1909),
.B1(n_1902),
.B2(n_1907),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1950),
.Y(n_1958)
);

AND4x2_ASAP7_75t_L g1959 ( 
.A(n_1948),
.B(n_1907),
.C(n_1893),
.D(n_1902),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1958),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1957),
.B(n_1953),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1959),
.B(n_1954),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1956),
.B(n_1952),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1955),
.B(n_1947),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1957),
.B(n_1907),
.Y(n_1965)
);

AOI321xp33_ASAP7_75t_L g1966 ( 
.A1(n_1964),
.A2(n_1910),
.A3(n_1888),
.B1(n_1889),
.B2(n_1892),
.C(n_1894),
.Y(n_1966)
);

AOI221x1_ASAP7_75t_L g1967 ( 
.A1(n_1960),
.A2(n_1867),
.B1(n_1872),
.B2(n_1887),
.C(n_1885),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1963),
.B(n_1895),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1965),
.Y(n_1969)
);

NOR2x1_ASAP7_75t_L g1970 ( 
.A(n_1960),
.B(n_1900),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1970),
.B(n_1961),
.Y(n_1971)
);

OAI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1968),
.A2(n_1962),
.B1(n_1900),
.B2(n_1899),
.Y(n_1972)
);

NOR2x1p5_ASAP7_75t_L g1973 ( 
.A(n_1966),
.B(n_1899),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1972),
.B(n_1969),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1974),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1971),
.B(n_1973),
.C(n_1967),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1975),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1977),
.Y(n_1978)
);

OAI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1976),
.A2(n_1854),
.B(n_1880),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_SL g1980 ( 
.A1(n_1978),
.A2(n_1979),
.B1(n_1865),
.B2(n_1836),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1886),
.B1(n_1885),
.B2(n_1880),
.C(n_1848),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1886),
.B(n_1865),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1849),
.B(n_1848),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_SL g1984 ( 
.A1(n_1983),
.A2(n_1849),
.B(n_1838),
.Y(n_1984)
);

AOI221xp5_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1829),
.B1(n_1838),
.B2(n_1847),
.C(n_1837),
.Y(n_1985)
);

OA22x2_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1847),
.B1(n_1840),
.B2(n_1837),
.Y(n_1986)
);


endmodule