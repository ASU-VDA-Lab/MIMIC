module fake_netlist_5_2451_n_1116 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1116);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1116;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_194;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_785;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_633;
wire n_307;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_186;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_1045;
wire n_297;
wire n_1079;
wire n_833;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_482;
wire n_342;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_866;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_239;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_1027;
wire n_971;
wire n_490;
wire n_805;
wire n_910;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_952;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_868;
wire n_803;
wire n_1092;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_73),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_61),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_20),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_21),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_96),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_22),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_93),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_86),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_25),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_142),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_107),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_23),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_83),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_137),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_48),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_156),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_49),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_146),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_170),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_152),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_77),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_154),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_35),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_78),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_117),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_178),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_11),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_108),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_181),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_179),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_183),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_194),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_206),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_182),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_187),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_191),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_196),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_199),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_198),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_210),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_207),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_189),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_201),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_192),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_212),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_218),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_233),
.B1(n_238),
.B2(n_247),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_193),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_195),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_250),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_203),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_258),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_278),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_248),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_204),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_251),
.B(n_209),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_213),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_274),
.A2(n_246),
.B1(n_245),
.B2(n_241),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_215),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_240),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_217),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_293),
.A2(n_220),
.B(n_219),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_254),
.A2(n_229),
.B1(n_237),
.B2(n_236),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_295),
.A2(n_224),
.B(n_198),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_262),
.A2(n_226),
.B(n_223),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_271),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_332),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_292),
.Y(n_357)
);

AO21x2_ASAP7_75t_L g358 ( 
.A1(n_345),
.A2(n_224),
.B(n_198),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_336),
.B(n_271),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_290),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_335),
.C(n_305),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_290),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_309),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

AO21x2_ASAP7_75t_L g380 ( 
.A1(n_345),
.A2(n_224),
.B(n_228),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_254),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_336),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_282),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_336),
.B(n_340),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_336),
.B(n_267),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_333),
.B(n_282),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_341),
.B(n_234),
.C(n_231),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_340),
.B(n_272),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_344),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

CKINVDCx6p67_ASAP7_75t_R g417 ( 
.A(n_339),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_318),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_318),
.Y(n_419)
);

NOR2x1p5_ASAP7_75t_L g420 ( 
.A(n_354),
.B(n_235),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_352),
.B(n_289),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_354),
.B(n_288),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_318),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_319),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_297),
.Y(n_431)
);

XOR2x2_ASAP7_75t_L g432 ( 
.A(n_362),
.B(n_303),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_400),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_417),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_323),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

XNOR2x2_ASAP7_75t_L g442 ( 
.A(n_383),
.B(n_303),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_378),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_297),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_344),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_325),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_352),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_327),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_388),
.B(n_369),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_372),
.B(n_325),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_372),
.A2(n_341),
.B(n_314),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_417),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_422),
.B(n_348),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_391),
.B(n_341),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_364),
.B(n_353),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_359),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_359),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_360),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_360),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_409),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_374),
.B(n_375),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_401),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_368),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_361),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_361),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_363),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_374),
.B(n_306),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_406),
.B(n_289),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_363),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_367),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_368),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_375),
.B(n_306),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_370),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_370),
.B(n_348),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_376),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_406),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_376),
.B(n_353),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_381),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_402),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_405),
.B(n_340),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_380),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_389),
.B(n_381),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_436),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_481),
.A2(n_306),
.B(n_324),
.C(n_314),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_457),
.B(n_353),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_481),
.A2(n_353),
.B1(n_316),
.B2(n_306),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_435),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_453),
.B(n_340),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_476),
.B(n_314),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_434),
.B(n_351),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_456),
.B(n_346),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_442),
.A2(n_351),
.B1(n_349),
.B2(n_358),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_439),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_449),
.B(n_346),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_314),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_434),
.B(n_346),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_440),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_429),
.B(n_324),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_455),
.A2(n_324),
.B(n_351),
.C(n_342),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_477),
.Y(n_538)
);

NAND2x1_ASAP7_75t_L g539 ( 
.A(n_452),
.B(n_366),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_438),
.B(n_324),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_348),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_491),
.B(n_389),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_447),
.B(n_348),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_474),
.B(n_338),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_395),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_348),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_395),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_350),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_507),
.B(n_346),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_458),
.B(n_397),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_489),
.A2(n_349),
.B1(n_358),
.B2(n_350),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_489),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_514),
.A2(n_380),
.B1(n_358),
.B2(n_224),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_479),
.B(n_350),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_461),
.A2(n_316),
.B1(n_397),
.B2(n_408),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_459),
.B(n_384),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_486),
.B(n_350),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_460),
.B(n_384),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_486),
.B(n_350),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_462),
.B(n_384),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_432),
.B(n_342),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_446),
.B(n_347),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_431),
.B(n_343),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_496),
.B(n_347),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_452),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_502),
.B(n_343),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_480),
.A2(n_385),
.B1(n_366),
.B2(n_377),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_463),
.B(n_385),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_464),
.B(n_347),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_467),
.B(n_385),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_508),
.A2(n_302),
.B(n_425),
.C(n_423),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_469),
.B(n_366),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_366),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_445),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_452),
.B(n_302),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_472),
.B(n_377),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_508),
.A2(n_316),
.B1(n_425),
.B2(n_423),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_487),
.A2(n_380),
.B1(n_224),
.B2(n_316),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_473),
.B(n_302),
.Y(n_585)
);

O2A1O1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_533),
.A2(n_518),
.B(n_537),
.C(n_517),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_533),
.B(n_471),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_471),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_534),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_566),
.B(n_433),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_SL g592 ( 
.A(n_536),
.B(n_433),
.C(n_239),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_524),
.B(n_504),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_525),
.B(n_522),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_548),
.A2(n_448),
.B1(n_451),
.B2(n_450),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_551),
.B(n_484),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_487),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_520),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_527),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_550),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

BUFx12f_ASAP7_75t_SL g603 ( 
.A(n_545),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_568),
.Y(n_604)
);

CKINVDCx6p67_ASAP7_75t_R g605 ( 
.A(n_534),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_535),
.B(n_483),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_571),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_545),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_550),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_531),
.A2(n_540),
.B1(n_580),
.B2(n_542),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_547),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_528),
.B(n_485),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_559),
.B(n_484),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_541),
.B(n_488),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_528),
.B(n_493),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_569),
.B(n_571),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_562),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_572),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_544),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_585),
.B(n_305),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_R g627 ( 
.A(n_543),
.B(n_505),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_572),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_546),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_549),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_494),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_581),
.B(n_552),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_553),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_515),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_572),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_563),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_555),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_523),
.B(n_331),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_SL g641 ( 
.A(n_532),
.B(n_511),
.C(n_498),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_574),
.Y(n_642)
);

NOR3xp33_ASAP7_75t_SL g643 ( 
.A(n_526),
.B(n_511),
.C(n_499),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_579),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_SL g647 ( 
.A(n_575),
.B(n_500),
.C(n_495),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_582),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_570),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_530),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_573),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_586),
.A2(n_577),
.B(n_519),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_598),
.B(n_512),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_605),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_629),
.B(n_555),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_598),
.B(n_513),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_586),
.A2(n_583),
.B(n_560),
.Y(n_657)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_651),
.A2(n_490),
.B(n_475),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_607),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_625),
.B(n_468),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_624),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_591),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_595),
.B(n_630),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_607),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_598),
.B(n_506),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_617),
.A2(n_501),
.B(n_506),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_634),
.A2(n_557),
.B(n_584),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_634),
.A2(n_584),
.B(n_557),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_608),
.A2(n_594),
.B(n_635),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_608),
.A2(n_398),
.B(n_509),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_638),
.A2(n_592),
.B1(n_620),
.B2(n_609),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_638),
.B(n_509),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_644),
.A2(n_465),
.B(n_503),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_638),
.B(n_224),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_637),
.A2(n_398),
.B(n_392),
.Y(n_676)
);

AOI21x1_ASAP7_75t_L g677 ( 
.A1(n_615),
.A2(n_503),
.B(n_418),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_468),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_640),
.A2(n_398),
.B(n_392),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_607),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_642),
.A2(n_398),
.B(n_392),
.Y(n_681)
);

OAI21x1_ASAP7_75t_SL g682 ( 
.A1(n_615),
.A2(n_418),
.B(n_414),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_600),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_645),
.A2(n_392),
.B(n_492),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_638),
.A2(n_492),
.B(n_427),
.C(n_419),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_633),
.A2(n_392),
.B(n_386),
.Y(n_686)
);

AOI21x1_ASAP7_75t_SL g687 ( 
.A1(n_619),
.A2(n_316),
.B(n_414),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_386),
.B(n_377),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_612),
.A2(n_377),
.B1(n_386),
.B2(n_396),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_331),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_621),
.A2(n_396),
.B(n_386),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_590),
.B(n_319),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_622),
.B(n_329),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_396),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_592),
.A2(n_632),
.B1(n_597),
.B2(n_603),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_619),
.A2(n_427),
.A3(n_419),
.B(n_307),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_621),
.A2(n_392),
.B(n_396),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_627),
.B(n_330),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_597),
.B(n_329),
.Y(n_699)
);

NAND2x1_ASAP7_75t_L g700 ( 
.A(n_593),
.B(n_316),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_649),
.A2(n_407),
.B(n_399),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_589),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_650),
.A2(n_407),
.B(n_399),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_587),
.A2(n_307),
.B1(n_328),
.B2(n_329),
.C(n_330),
.Y(n_704)
);

AOI21xp33_ASAP7_75t_L g705 ( 
.A1(n_588),
.A2(n_328),
.B(n_330),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_611),
.B(n_330),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_648),
.A2(n_407),
.B(n_399),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_606),
.A2(n_614),
.B(n_613),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_646),
.B(n_316),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_636),
.B(n_31),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_611),
.B(n_330),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_646),
.B(n_0),
.Y(n_712)
);

NAND2x1_ASAP7_75t_L g713 ( 
.A(n_682),
.B(n_623),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_661),
.B(n_663),
.Y(n_714)
);

OA21x2_ASAP7_75t_L g715 ( 
.A1(n_652),
.A2(n_641),
.B(n_643),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_654),
.Y(n_716)
);

AO31x2_ASAP7_75t_L g717 ( 
.A1(n_685),
.A2(n_623),
.A3(n_628),
.B(n_618),
.Y(n_717)
);

AO32x2_ASAP7_75t_L g718 ( 
.A1(n_689),
.A2(n_628),
.A3(n_641),
.B1(n_647),
.B2(n_643),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_655),
.B(n_602),
.Y(n_719)
);

OA21x2_ASAP7_75t_L g720 ( 
.A1(n_691),
.A2(n_647),
.B(n_596),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_706),
.B(n_639),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_672),
.A2(n_631),
.B(n_616),
.Y(n_722)
);

OAI22x1_ASAP7_75t_L g723 ( 
.A1(n_653),
.A2(n_632),
.B1(n_631),
.B2(n_599),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_692),
.Y(n_724)
);

BUFx8_ASAP7_75t_L g725 ( 
.A(n_710),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_712),
.B(n_616),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_683),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_SL g728 ( 
.A1(n_671),
.A2(n_702),
.B1(n_695),
.B2(n_669),
.C(n_690),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_660),
.B(n_601),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_675),
.A2(n_710),
.B1(n_656),
.B2(n_653),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_672),
.A2(n_610),
.B(n_601),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_668),
.A2(n_610),
.B(n_626),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_662),
.B(n_626),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_665),
.B(n_656),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_694),
.B(n_626),
.Y(n_735)
);

CKINVDCx11_ASAP7_75t_R g736 ( 
.A(n_659),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_667),
.A2(n_657),
.B(n_675),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_670),
.A2(n_312),
.B(n_416),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_659),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_705),
.A2(n_312),
.B(n_416),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_699),
.B(n_32),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_659),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_693),
.B(n_33),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_711),
.B(n_0),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_664),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_665),
.A2(n_312),
.B1(n_416),
.B2(n_3),
.Y(n_746)
);

CKINVDCx6p67_ASAP7_75t_R g747 ( 
.A(n_664),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_678),
.B(n_1),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_708),
.Y(n_749)
);

AO21x2_ASAP7_75t_L g750 ( 
.A1(n_658),
.A2(n_36),
.B(n_34),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_664),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_SL g752 ( 
.A(n_698),
.B(n_2),
.C(n_3),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_709),
.B(n_2),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_680),
.B(n_4),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_704),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_696),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_677),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_673),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_688),
.A2(n_38),
.B(n_37),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_680),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_696),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_673),
.B(n_7),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_676),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_696),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_679),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

AO31x2_ASAP7_75t_L g767 ( 
.A1(n_684),
.A2(n_686),
.A3(n_681),
.B(n_697),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_700),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_674),
.A2(n_40),
.B(n_39),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_666),
.A2(n_113),
.A3(n_176),
.B(n_174),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_707),
.A2(n_177),
.B(n_43),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_703),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_772)
);

OA21x2_ASAP7_75t_L g773 ( 
.A1(n_701),
.A2(n_44),
.B(n_42),
.Y(n_773)
);

AO31x2_ASAP7_75t_L g774 ( 
.A1(n_652),
.A2(n_114),
.A3(n_172),
.B(n_171),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_663),
.B(n_12),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_652),
.A2(n_111),
.A3(n_169),
.B(n_168),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_662),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_691),
.A2(n_110),
.B(n_163),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_672),
.B(n_13),
.Y(n_779)
);

AOI21xp33_ASAP7_75t_L g780 ( 
.A1(n_655),
.A2(n_14),
.B(n_16),
.Y(n_780)
);

BUFx2_ASAP7_75t_R g781 ( 
.A(n_661),
.Y(n_781)
);

AO31x2_ASAP7_75t_L g782 ( 
.A1(n_652),
.A2(n_109),
.A3(n_162),
.B(n_161),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_725),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_780),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_737),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_752),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_753),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_725),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_745),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_777),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_755),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_766),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_756),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_733),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_736),
.Y(n_796)
);

CKINVDCx11_ASAP7_75t_R g797 ( 
.A(n_716),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_714),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_R g799 ( 
.A1(n_724),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_743),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_719),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_764),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_730),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_721),
.B(n_47),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_723),
.Y(n_805)
);

INVx3_ASAP7_75t_SL g806 ( 
.A(n_747),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_726),
.B(n_50),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_779),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_739),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_745),
.Y(n_810)
);

INVx6_ASAP7_75t_L g811 ( 
.A(n_734),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_734),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_746),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_815)
);

CKINVDCx6p67_ASAP7_75t_R g816 ( 
.A(n_754),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_751),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_741),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_781),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_757),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_761),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_728),
.B(n_63),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_735),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_729),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_775),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_717),
.Y(n_826)
);

CKINVDCx11_ASAP7_75t_R g827 ( 
.A(n_768),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_760),
.Y(n_828)
);

INVx4_ASAP7_75t_SL g829 ( 
.A(n_774),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_765),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_758),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_SL g832 ( 
.A1(n_715),
.A2(n_722),
.B1(n_748),
.B2(n_750),
.Y(n_832)
);

INVx6_ASAP7_75t_L g833 ( 
.A(n_768),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_744),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_717),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_713),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_770),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_762),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_770),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_715),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_840)
);

BUFx4_ASAP7_75t_R g841 ( 
.A(n_718),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_718),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_720),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_713),
.Y(n_844)
);

BUFx2_ASAP7_75t_SL g845 ( 
.A(n_731),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_720),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_774),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_823),
.B(n_90),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_812),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_794),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_802),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_825),
.A2(n_763),
.B(n_772),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_798),
.B(n_732),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_805),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_790),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_820),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_821),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_826),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_799),
.A2(n_771),
.B1(n_769),
.B2(n_773),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_835),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_839),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_793),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_792),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_847),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_836),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_824),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_842),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_846),
.B(n_776),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_837),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_791),
.A2(n_773),
.B1(n_740),
.B2(n_776),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_844),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_844),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_829),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_792),
.B(n_778),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_795),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_834),
.B(n_782),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_829),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_829),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_841),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_811),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_845),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_822),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_822),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_832),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_792),
.B(n_759),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_828),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_789),
.B(n_738),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_834),
.B(n_782),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_791),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_792),
.B(n_767),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_811),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_843),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_809),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_806),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_872),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_849),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_851),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_897),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_855),
.B(n_843),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_895),
.A2(n_786),
.B1(n_800),
.B2(n_785),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_856),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_892),
.Y(n_906)
);

HB1xp67_ASAP7_75t_SL g907 ( 
.A(n_850),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_879),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_856),
.Y(n_909)
);

OA21x2_ASAP7_75t_L g910 ( 
.A1(n_885),
.A2(n_807),
.B(n_840),
.Y(n_910)
);

INVxp67_ASAP7_75t_R g911 ( 
.A(n_877),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_869),
.B(n_804),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_851),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_894),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_869),
.B(n_801),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_892),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_852),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_885),
.B(n_814),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_897),
.B(n_797),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_894),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_857),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_857),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_868),
.B(n_767),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_879),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_882),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_872),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_862),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_891),
.B(n_817),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_882),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_898),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_928),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_917),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_898),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_902),
.B(n_850),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_917),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_928),
.Y(n_937)
);

OR2x6_ASAP7_75t_L g938 ( 
.A(n_908),
.B(n_893),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_901),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_926),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_899),
.B(n_900),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_899),
.B(n_891),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_901),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_919),
.B(n_877),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_908),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_911),
.B(n_880),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_913),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_919),
.B(n_889),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_911),
.B(n_880),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_913),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_925),
.B(n_889),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_925),
.B(n_893),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_918),
.Y(n_953)
);

OAI211xp5_ASAP7_75t_SL g954 ( 
.A1(n_906),
.A2(n_853),
.B(n_854),
.C(n_860),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_918),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_951),
.B(n_915),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_915),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_937),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_937),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_916),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_944),
.B(n_930),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_938),
.B(n_898),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_946),
.B(n_949),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_932),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_954),
.A2(n_895),
.B1(n_903),
.B2(n_904),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_945),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_948),
.B(n_929),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_SL g968 ( 
.A(n_949),
.B(n_902),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_932),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_940),
.B(n_929),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_947),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_912),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_963),
.B(n_952),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_961),
.B(n_942),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_962),
.B(n_945),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_963),
.B(n_938),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_967),
.B(n_942),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_956),
.B(n_938),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_956),
.B(n_938),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_941),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_966),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_971),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_957),
.B(n_914),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_957),
.B(n_931),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_980),
.B(n_965),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_974),
.B(n_960),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_982),
.B(n_920),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_968),
.C(n_848),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_977),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_975),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_960),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_985),
.A2(n_975),
.B1(n_968),
.B2(n_904),
.C(n_935),
.Y(n_993)
);

AO221x2_ASAP7_75t_L g994 ( 
.A1(n_988),
.A2(n_907),
.B1(n_964),
.B2(n_969),
.C(n_958),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_991),
.B(n_783),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_987),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_988),
.B(n_973),
.Y(n_997)
);

NOR2x1_ASAP7_75t_L g998 ( 
.A(n_990),
.B(n_796),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_998),
.B(n_992),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_996),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_997),
.B(n_986),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_995),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_989),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_993),
.B(n_979),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_998),
.B(n_978),
.Y(n_1005)
);

CKINVDCx16_ASAP7_75t_R g1006 ( 
.A(n_995),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_997),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_997),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1000),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_SL g1010 ( 
.A1(n_1003),
.A2(n_819),
.B1(n_903),
.B2(n_979),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1000),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1002),
.B(n_984),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1006),
.A2(n_819),
.B1(n_788),
.B2(n_976),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1002),
.B(n_984),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_999),
.B(n_1005),
.Y(n_1015)
);

NAND4xp25_ASAP7_75t_L g1016 ( 
.A(n_1007),
.B(n_976),
.C(n_784),
.D(n_890),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_1008),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_SL g1018 ( 
.A1(n_1012),
.A2(n_1014),
.B1(n_1004),
.B2(n_1010),
.C(n_1001),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1011),
.B(n_1004),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_787),
.C(n_825),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_1013),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_962),
.B1(n_959),
.B2(n_958),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_1013),
.Y(n_1023)
);

XNOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_803),
.Y(n_1024)
);

AOI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_1021),
.A2(n_807),
.B(n_838),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1023),
.B(n_972),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_827),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_972),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_1017),
.A2(n_815),
.B(n_871),
.C(n_818),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1020),
.A2(n_962),
.B1(n_808),
.B2(n_959),
.C(n_830),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1022),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1026),
.B(n_1024),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_1027),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1031),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1029),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1025),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1030),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1026),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1026),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_SL g1041 ( 
.A(n_1031),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1026),
.Y(n_1042)
);

NAND4xp75_ASAP7_75t_L g1043 ( 
.A(n_1039),
.B(n_910),
.C(n_874),
.D(n_878),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1040),
.A2(n_921),
.B(n_914),
.C(n_883),
.Y(n_1044)
);

OA22x2_ASAP7_75t_L g1045 ( 
.A1(n_1035),
.A2(n_810),
.B1(n_864),
.B2(n_931),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1034),
.B(n_810),
.C(n_831),
.Y(n_1046)
);

NAND4xp25_ASAP7_75t_L g1047 ( 
.A(n_1032),
.B(n_864),
.C(n_912),
.D(n_884),
.Y(n_1047)
);

NAND4xp75_ASAP7_75t_L g1048 ( 
.A(n_1038),
.B(n_910),
.C(n_874),
.D(n_878),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_1034),
.B(n_921),
.C(n_914),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1042),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1033),
.B(n_864),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1037),
.B(n_883),
.C(n_884),
.Y(n_1052)
);

NOR4xp25_ASAP7_75t_L g1053 ( 
.A(n_1036),
.B(n_953),
.C(n_933),
.D(n_950),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1050),
.B(n_1034),
.C(n_1041),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_1049),
.B(n_914),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_1051),
.B(n_914),
.C(n_921),
.Y(n_1056)
);

NOR4xp25_ASAP7_75t_L g1057 ( 
.A(n_1046),
.B(n_955),
.C(n_950),
.D(n_943),
.Y(n_1057)
);

NAND4xp25_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_881),
.C(n_887),
.D(n_896),
.Y(n_1058)
);

NOR5xp2_ASAP7_75t_L g1059 ( 
.A(n_1045),
.B(n_862),
.C(n_865),
.D(n_861),
.E(n_859),
.Y(n_1059)
);

AOI211xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1044),
.A2(n_867),
.B(n_881),
.C(n_934),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1052),
.B(n_921),
.C(n_896),
.Y(n_1061)
);

AO221x1_ASAP7_75t_L g1062 ( 
.A1(n_1054),
.A2(n_1053),
.B1(n_1048),
.B2(n_1043),
.C(n_921),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1055),
.A2(n_887),
.B(n_888),
.Y(n_1063)
);

OAI211xp5_ASAP7_75t_SL g1064 ( 
.A1(n_1060),
.A2(n_881),
.B(n_941),
.C(n_863),
.Y(n_1064)
);

AOI221xp5_ASAP7_75t_L g1065 ( 
.A1(n_1057),
.A2(n_931),
.B1(n_934),
.B2(n_939),
.C(n_943),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1056),
.A2(n_934),
.B1(n_939),
.B2(n_955),
.C(n_936),
.Y(n_1066)
);

NAND5xp2_ASAP7_75t_L g1067 ( 
.A(n_1059),
.B(n_875),
.C(n_886),
.D(n_865),
.E(n_100),
.Y(n_1067)
);

OAI211xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1061),
.A2(n_863),
.B(n_876),
.C(n_936),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1058),
.Y(n_1069)
);

AOI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_894),
.B(n_893),
.C(n_876),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_1069),
.B(n_1063),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1067),
.B(n_97),
.C(n_98),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_L g1073 ( 
.A(n_1064),
.B(n_99),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_1062),
.Y(n_1074)
);

NAND3x1_ASAP7_75t_L g1075 ( 
.A(n_1065),
.B(n_927),
.C(n_898),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1070),
.B(n_922),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1068),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1066),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1069),
.B(n_101),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1062),
.B(n_922),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1072),
.B(n_894),
.Y(n_1081)
);

XOR2x2_ASAP7_75t_L g1082 ( 
.A(n_1079),
.B(n_104),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_1080),
.B(n_105),
.C(n_106),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_SL g1084 ( 
.A(n_1074),
.B(n_875),
.C(n_886),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1073),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_1071),
.B(n_833),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1077),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1078),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1076),
.B(n_115),
.C(n_116),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_1075),
.B(n_888),
.C(n_894),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_1071),
.Y(n_1091)
);

AND3x4_ASAP7_75t_L g1092 ( 
.A(n_1072),
.B(n_873),
.C(n_833),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_1085),
.B(n_875),
.C(n_886),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_833),
.B1(n_888),
.B2(n_866),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1088),
.A2(n_1087),
.B1(n_1086),
.B2(n_1092),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1081),
.A2(n_910),
.B1(n_888),
.B2(n_866),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1082),
.A2(n_910),
.B(n_923),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1083),
.Y(n_1098)
);

XNOR2xp5_ASAP7_75t_L g1099 ( 
.A(n_1089),
.B(n_118),
.Y(n_1099)
);

AO22x2_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_1084),
.B1(n_1090),
.B2(n_927),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_923),
.B1(n_909),
.B2(n_905),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1095),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1094),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1093),
.A2(n_861),
.B1(n_859),
.B2(n_924),
.Y(n_1104)
);

OAI22x1_ASAP7_75t_L g1105 ( 
.A1(n_1096),
.A2(n_858),
.B1(n_870),
.B2(n_924),
.Y(n_1105)
);

XNOR2xp5_ASAP7_75t_L g1106 ( 
.A(n_1102),
.B(n_1097),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1100),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1103),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_1105),
.B1(n_1104),
.B2(n_1101),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1109),
.A2(n_1107),
.B(n_1106),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_1110),
.Y(n_1111)
);

AO22x2_ASAP7_75t_L g1112 ( 
.A1(n_1111),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1112),
.B(n_858),
.Y(n_1113)
);

AO221x2_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.C(n_132),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_140),
.B(n_141),
.C(n_145),
.Y(n_1116)
);


endmodule