module real_jpeg_12178_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_296, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_296;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_215;
wire n_221;
wire n_292;
wire n_288;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_3),
.A2(n_37),
.B1(n_60),
.B2(n_63),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_68),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_7),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_134),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_134),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_10),
.A2(n_60),
.B1(n_63),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_79),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_79),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_12),
.A2(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_70),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_13),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_65),
.B(n_161),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_152),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_44),
.B(n_49),
.C(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_13),
.B(n_109),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_33),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_13),
.B(n_54),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_13),
.A2(n_63),
.B(n_73),
.C(n_223),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_14),
.A2(n_46),
.B1(n_60),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_46),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_14),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_15),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_102),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_16),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_271),
.B1(n_293),
.B2(n_294),
.Y(n_19)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_124),
.B(n_270),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_22),
.B(n_103),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.C(n_87),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_23),
.B(n_81),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_57),
.C(n_71),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_256)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_28),
.A2(n_33),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_28),
.A2(n_33),
.B1(n_141),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_28),
.A2(n_33),
.B1(n_93),
.B2(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_28),
.A2(n_33),
.B1(n_155),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_28),
.A2(n_33),
.B1(n_152),
.B2(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_28),
.A2(n_33),
.B1(n_201),
.B2(n_208),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_29),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_32),
.A2(n_35),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_32),
.A2(n_91),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_36),
.A2(n_50),
.B(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_51),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_45),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_44),
.B(n_76),
.Y(n_153)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_45),
.A2(n_63),
.A3(n_75),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_54),
.B1(n_85),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_47),
.A2(n_54),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_47),
.A2(n_54),
.B1(n_96),
.B2(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_47),
.A2(n_54),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_47),
.A2(n_54),
.B1(n_187),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_47),
.A2(n_54),
.B(n_111),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_51),
.A2(n_97),
.B1(n_145),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_58),
.A2(n_59),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_58),
.A2(n_59),
.B1(n_120),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_60),
.B(n_152),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_162),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_61),
.B(n_63),
.Y(n_176)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_66),
.B(n_152),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_72),
.A2(n_77),
.B1(n_136),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_109),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_73),
.A2(n_109),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_73),
.A2(n_108),
.B1(n_109),
.B2(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_77),
.A2(n_133),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_83),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_83),
.A2(n_119),
.B(n_121),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_87),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.C(n_100),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_88),
.A2(n_89),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_90),
.B(n_94),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_98),
.B(n_100),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_99),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_101),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_123),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_112),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_112),
.A2(n_277),
.B1(n_289),
.B2(n_290),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_112),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_291)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_265),
.B(n_269),
.Y(n_124)
);

OAI221xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_252),
.B1(n_263),
.B2(n_264),
.C(n_296),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_236),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_179),
.B(n_235),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_156),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_129),
.B(n_156),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_143),
.C(n_147),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_138),
.C(n_140),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_139),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_147),
.B1(n_148),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_143),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_151),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_170),
.B2(n_178),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_157),
.B(n_171),
.C(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_159),
.B(n_165),
.C(n_169),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_172),
.B(n_175),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_229),
.B(n_234),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_217),
.B(n_228),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_197),
.B(n_216),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_205),
.B(n_215),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_203),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_214),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_238),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_247),
.C(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_261),
.C(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_292),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_291),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule