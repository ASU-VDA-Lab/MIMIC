module fake_jpeg_11508_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_18),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_58),
.Y(n_67)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_75),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_37),
.B1(n_36),
.B2(n_26),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_44),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_95),
.B1(n_97),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_82),
.B(n_90),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_32),
.B(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_91),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_32),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_31),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_20),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_100),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_106),
.Y(n_143)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_42),
.B1(n_50),
.B2(n_41),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_84),
.B1(n_80),
.B2(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_128),
.B1(n_92),
.B2(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_46),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_84),
.B1(n_85),
.B2(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_1),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_122),
.Y(n_150)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_2),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_12),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_4),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_68),
.C(n_94),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_97),
.B(n_69),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_133),
.B(n_109),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_98),
.B(n_83),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_129),
.B1(n_124),
.B2(n_119),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_92),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_80),
.B1(n_68),
.B2(n_88),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_106),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_152),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_88),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_112),
.B(n_101),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_125),
.C(n_103),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_92),
.C(n_7),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_4),
.Y(n_161)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_164),
.Y(n_183)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_110),
.CON(n_167),
.SN(n_167)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_172),
.B(n_132),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_115),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_12),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_133),
.B(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_151),
.B1(n_141),
.B2(n_149),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_143),
.B1(n_144),
.B2(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_188),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_146),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_185),
.B(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_152),
.B(n_130),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_154),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_157),
.B1(n_162),
.B2(n_171),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_194),
.B1(n_198),
.B2(n_177),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_173),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_181),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_157),
.B1(n_175),
.B2(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_158),
.B1(n_137),
.B2(n_131),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_159),
.B1(n_143),
.B2(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_159),
.B1(n_164),
.B2(n_100),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_202),
.C(n_183),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_212),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_178),
.C(n_185),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_213),
.C(n_203),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_194),
.B1(n_198),
.B2(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_189),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_122),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_183),
.C(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_218),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_204),
.B1(n_187),
.B2(n_191),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_213),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_14),
.B(n_7),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_207),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_216),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_217),
.C(n_214),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_228),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_214),
.C(n_209),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_227),
.C(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_231),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_224),
.Y(n_234)
);


endmodule