module real_jpeg_1455_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_1),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_1),
.A2(n_27),
.B1(n_71),
.B2(n_74),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_73),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_73),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_5),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_34),
.B1(n_71),
.B2(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_34),
.B1(n_59),
.B2(n_60),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_38),
.B1(n_71),
.B2(n_74),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_60),
.C(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_6),
.B(n_66),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_6),
.B(n_39),
.C(n_54),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_23),
.C(n_45),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_52),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_30),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_49),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_318),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_310),
.B(n_317),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_272),
.B(n_307),
.Y(n_14)
);

A2O1A1O1Ixp25_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_134),
.B(n_252),
.C(n_253),
.D(n_271),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_112),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_112),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_18),
.B(n_80),
.C(n_106),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_51),
.C(n_63),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_19),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_20),
.B(n_35),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_21),
.A2(n_29),
.B(n_87),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_47)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_23),
.B(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_28),
.B(n_33),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_28),
.A2(n_29),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_28),
.B(n_86),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_28),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_29),
.B(n_216),
.Y(n_230)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_30),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_31),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_32),
.B(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_48),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_36),
.B(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_37),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_37),
.B(n_49),
.Y(n_187)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_39),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_42),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI21x1_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_90),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_48),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_49),
.B(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_51),
.A2(n_63),
.B1(n_64),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_51),
.A2(n_116),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_51),
.B(n_314),
.C(n_316),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_62),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_52),
.B(n_62),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_52),
.B(n_127),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_52),
.A2(n_153),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_56),
.B(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_57),
.B(n_102),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_57),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_60),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_66),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_70),
.B(n_76),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_75),
.A2(n_264),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_75),
.B(n_95),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_105),
.B2(n_106),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_92),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_82),
.B(n_93),
.C(n_100),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_84),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_87),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_88)
);

AOI21x1_ASAP7_75t_SL g150 ( 
.A1(n_89),
.A2(n_110),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_91),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_91),
.B(n_187),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_97),
.B(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_97),
.A2(n_148),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_101),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_104),
.B(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_107),
.A2(n_108),
.B1(n_182),
.B2(n_183),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_107),
.A2(n_108),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_108),
.B(n_109),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_108),
.A2(n_260),
.B(n_262),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_133),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_114),
.B1(n_133),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_128),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_120),
.B(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_120),
.A2(n_148),
.B(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_156),
.B(n_249),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_136),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_137),
.B(n_140),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_147),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_149),
.A2(n_150),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_149),
.A2(n_150),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_150),
.B(n_280),
.C(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_150),
.B(n_304),
.C(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_153),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_160),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_162),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_230),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_193),
.B(n_248),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_190),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_185),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_178),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21x1_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_204),
.B(n_247),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_202),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_245),
.Y(n_244)
);

OAI21x1_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_242),
.B(n_246),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_224),
.B(n_241),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_221),
.C(n_223),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_231),
.B(n_240),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_228),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_236),
.B(n_239),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_255),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_258),
.C(n_266),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_265),
.B2(n_266),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_270),
.A2(n_278),
.B1(n_279),
.B2(n_289),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_270),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_276),
.C(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_290),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_275),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_281),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_293),
.C(n_297),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_285),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_306),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_320),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);


endmodule