module fake_jpeg_3706_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_13),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_49),
.Y(n_77)
);

OR2x4_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_27),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_52),
.B1(n_63),
.B2(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_3),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_24),
.B(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_3),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_4),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_11),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_49),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_101),
.C(n_60),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_86),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_82),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_60),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_79),
.B(n_74),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_73),
.B1(n_84),
.B2(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_109),
.B1(n_101),
.B2(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_84),
.B1(n_89),
.B2(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_72),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_94),
.C(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_115),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_76),
.A3(n_48),
.B1(n_64),
.B2(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_90),
.B(n_58),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_52),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.C(n_112),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_102),
.C(n_96),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_124),
.B(n_111),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_92),
.B(n_95),
.C(n_105),
.D(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_126),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_114),
.C(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

AO221x1_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_111),
.B1(n_70),
.B2(n_68),
.C(n_51),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_130),
.B1(n_118),
.B2(n_117),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_55),
.C(n_50),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_122),
.C(n_127),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_131),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_65),
.B(n_55),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_137),
.B1(n_65),
.B2(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_131),
.Y(n_142)
);


endmodule