module fake_netlist_5_1711_n_102 (n_8, n_4, n_5, n_7, n_0, n_2, n_3, n_6, n_1, n_102);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_2;
input n_3;
input n_6;
input n_1;

output n_102;

wire n_91;
wire n_82;
wire n_10;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_13;
wire n_66;
wire n_98;
wire n_60;
wire n_16;
wire n_43;
wire n_69;
wire n_9;
wire n_58;
wire n_18;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_17;
wire n_92;
wire n_19;
wire n_30;
wire n_33;
wire n_14;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_12;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_11;
wire n_15;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp67_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_11),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_9),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_18),
.B(n_23),
.Y(n_32)
);

OAI21x1_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_23),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_20),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_20),
.B(n_21),
.C(n_10),
.Y(n_35)
);

AO31x2_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_0),
.A3(n_20),
.B(n_5),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_4),
.Y(n_38)
);

AO31x2_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_4),
.A3(n_6),
.B(n_7),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_25),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_7),
.B1(n_24),
.B2(n_28),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_24),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_26),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_34),
.B(n_44),
.C(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_33),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_37),
.B1(n_41),
.B2(n_38),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_32),
.B(n_35),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_34),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_34),
.B(n_28),
.C(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_48),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_54),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_57),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_49),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g72 ( 
.A(n_64),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_63),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_63),
.B1(n_64),
.B2(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

OAI31xp33_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_62),
.A3(n_61),
.B(n_45),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_70),
.B1(n_57),
.B2(n_68),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_78),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_74),
.B1(n_77),
.B2(n_53),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_56),
.C(n_80),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_75),
.B1(n_73),
.B2(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_57),
.B1(n_52),
.B2(n_72),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_84),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_51),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

OAI211xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_51),
.B(n_50),
.C(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI322xp33_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_91),
.A3(n_90),
.B1(n_58),
.B2(n_60),
.C1(n_53),
.C2(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_93),
.B(n_90),
.Y(n_99)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_95),
.B1(n_75),
.B2(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_99),
.B1(n_75),
.B2(n_67),
.Y(n_102)
);


endmodule