module fake_ariane_1590_n_2149 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2149);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2149;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_2144;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_602;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_1789;
wire n_763;
wire n_1986;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_1579;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_346),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_378),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_21),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_573),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_562),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_541),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_527),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_24),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_387),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_565),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_170),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_350),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_117),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_423),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_449),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_193),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_192),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_325),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_106),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_406),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_180),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_154),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_421),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_121),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_463),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_9),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_190),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_34),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_104),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_127),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_171),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_428),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_241),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_567),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_537),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_400),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_4),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_150),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_54),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_255),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_390),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_557),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_88),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_569),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_570),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_285),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_158),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_145),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_480),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_114),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_228),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_560),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_382),
.Y(n_652)
);

BUFx8_ASAP7_75t_SL g653 ( 
.A(n_427),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_21),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_243),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_118),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_108),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_572),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_65),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_364),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_413),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_580),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_512),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_74),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_65),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_49),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_252),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_175),
.Y(n_669)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_47),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_296),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_352),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_568),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_181),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_578),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_418),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_253),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_333),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_259),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_113),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_407),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_183),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_425),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_517),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_334),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_268),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_353),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_184),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_419),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_368),
.Y(n_691)
);

CKINVDCx14_ASAP7_75t_R g692 ( 
.A(n_148),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_116),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_46),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_389),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_412),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_404),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_197),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_129),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_571),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_91),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_202),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_484),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_360),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_513),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_561),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_6),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_485),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_410),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_263),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_577),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_431),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_494),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_179),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_161),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_75),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_142),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_579),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_299),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_447),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_254),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_384),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_75),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_466),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_581),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_29),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_381),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_388),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_143),
.Y(n_730)
);

CKINVDCx14_ASAP7_75t_R g731 ( 
.A(n_540),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_113),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_351),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_401),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_3),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_342),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_452),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_62),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_149),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_91),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_118),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_67),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_278),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_45),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_312),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_277),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_200),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_25),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_160),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_576),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_488),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_187),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_95),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_63),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_182),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_173),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_495),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_264),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_47),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_240),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_554),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_454),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_566),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_344),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_487),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_511),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_45),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_82),
.Y(n_769)
);

BUFx8_ASAP7_75t_SL g770 ( 
.A(n_475),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_195),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_530),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_624),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_625),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_634),
.Y(n_775)
);

INVxp33_ASAP7_75t_SL g776 ( 
.A(n_599),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_654),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_679),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_636),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_642),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_628),
.B(n_1),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_670),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_649),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_653),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_667),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_680),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_707),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_724),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_727),
.Y(n_789)
);

INVxp33_ASAP7_75t_SL g790 ( 
.A(n_609),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_604),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_732),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_741),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_768),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_622),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_657),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_658),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_744),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_749),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_760),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_769),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_745),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_685),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_720),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_602),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_615),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_702),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_679),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_679),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_770),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_702),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_610),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_735),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_717),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_735),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_620),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_608),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_616),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_692),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_731),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_641),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_618),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_627),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_631),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_637),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_688),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_639),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_669),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_626),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_673),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_691),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_674),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_695),
.Y(n_836)
);

CKINVDCx14_ASAP7_75t_R g837 ( 
.A(n_711),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_698),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_660),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_706),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_718),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_686),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_686),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_721),
.Y(n_846)
);

INVxp33_ASAP7_75t_SL g847 ( 
.A(n_665),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_746),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_686),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_747),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_763),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_755),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_666),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_764),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_765),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_767),
.Y(n_856)
);

INVxp33_ASAP7_75t_SL g857 ( 
.A(n_693),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_694),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_699),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_701),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_738),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_740),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_742),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_754),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_758),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_597),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_696),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_629),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_655),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_758),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_681),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_598),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_600),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_865),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_778),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_778),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_778),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_799),
.B(n_613),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_810),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_810),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_810),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_852),
.A2(n_656),
.B1(n_652),
.B2(n_710),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_829),
.B(n_715),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_831),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_809),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_777),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_811),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_811),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_866),
.B(n_736),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_808),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_845),
.Y(n_891)
);

OAI21x1_ASAP7_75t_L g892 ( 
.A1(n_819),
.A2(n_750),
.B(n_762),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_813),
.B(n_758),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_872),
.B(n_601),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_873),
.B(n_603),
.Y(n_896)
);

OAI22x1_ASAP7_75t_R g897 ( 
.A1(n_853),
.A2(n_606),
.B1(n_607),
.B2(n_605),
.Y(n_897)
);

BUFx8_ASAP7_75t_SL g898 ( 
.A(n_806),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_814),
.Y(n_899)
);

OAI21x1_ASAP7_75t_L g900 ( 
.A1(n_820),
.A2(n_762),
.B(n_612),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_773),
.Y(n_901)
);

BUFx12f_ASAP7_75t_L g902 ( 
.A(n_784),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_823),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_858),
.B(n_611),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_775),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_811),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_839),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_779),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_822),
.A2(n_762),
.B(n_619),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_844),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_844),
.Y(n_912)
);

CKINVDCx6p67_ASAP7_75t_R g913 ( 
.A(n_802),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_818),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_832),
.B(n_614),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_870),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_812),
.B(n_621),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_859),
.B(n_623),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_825),
.B(n_762),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_785),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_870),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_870),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_787),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_782),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_776),
.B(n_790),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_774),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_860),
.B(n_630),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_789),
.Y(n_929)
);

OA21x2_ASAP7_75t_L g930 ( 
.A1(n_826),
.A2(n_635),
.B(n_633),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_783),
.B(n_638),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_791),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_864),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_803),
.Y(n_934)
);

INVx5_ASAP7_75t_L g935 ( 
.A(n_821),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_868),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_795),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_792),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_796),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_797),
.Y(n_940)
);

AOI22x1_ASAP7_75t_SL g941 ( 
.A1(n_824),
.A2(n_643),
.B1(n_644),
.B2(n_640),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_793),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_804),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_862),
.B(n_645),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_827),
.A2(n_647),
.B(n_646),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_798),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_794),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_828),
.A2(n_762),
.B(n_650),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_835),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_863),
.B(n_648),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_805),
.B(n_651),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_869),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_800),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_833),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_801),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_867),
.B(n_659),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_871),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_807),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_847),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_937),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_901),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_939),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_884),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_874),
.B(n_816),
.Y(n_965)
);

NOR2x1_ASAP7_75t_L g966 ( 
.A(n_907),
.B(n_815),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_936),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_896),
.B(n_830),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_926),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_905),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_908),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_874),
.B(n_915),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_885),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_920),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_926),
.Y(n_975)
);

AND2x6_ASAP7_75t_L g976 ( 
.A(n_931),
.B(n_834),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_923),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_931),
.B(n_836),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_929),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_936),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_939),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_924),
.B(n_837),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_932),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_891),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_953),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_893),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_894),
.B(n_817),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_878),
.B(n_780),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_892),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_953),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_952),
.Y(n_991)
);

XNOR2xp5_ASAP7_75t_L g992 ( 
.A(n_882),
.B(n_861),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_957),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_886),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_928),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_878),
.B(n_838),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_938),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_950),
.B(n_840),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_942),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_947),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_940),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_946),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_889),
.B(n_841),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_910),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_883),
.B(n_842),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_955),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_SL g1007 ( 
.A1(n_899),
.A2(n_857),
.B1(n_781),
.B2(n_786),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_877),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_911),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_875),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_879),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_954),
.Y(n_1012)
);

XOR2xp5_ASAP7_75t_L g1013 ( 
.A(n_949),
.B(n_843),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_906),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_877),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_880),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_880),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_875),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_881),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_895),
.B(n_846),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_881),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_887),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_887),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_917),
.B(n_890),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_888),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_888),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_916),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_916),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_934),
.B(n_856),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_921),
.Y(n_1030)
);

CKINVDCx8_ASAP7_75t_R g1031 ( 
.A(n_935),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_904),
.B(n_848),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_935),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_921),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_922),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_922),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_903),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_956),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_902),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_913),
.B(n_661),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_943),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_918),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_898),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_900),
.A2(n_851),
.B(n_850),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_927),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_876),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_944),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_876),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_919),
.B(n_854),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_912),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_919),
.B(n_855),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_933),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_919),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_1039),
.B(n_958),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1015),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_1029),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_1031),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_983),
.B(n_925),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_1043),
.B(n_958),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_967),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_965),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_968),
.B(n_914),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1042),
.B(n_959),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_L g1064 ( 
.A(n_1045),
.B(n_959),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_967),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1001),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_L g1067 ( 
.A(n_1047),
.B(n_762),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_1033),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_998),
.B(n_951),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_965),
.B(n_662),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_984),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1020),
.A2(n_945),
.B1(n_930),
.B2(n_697),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1038),
.B(n_941),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_985),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_986),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1012),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1052),
.B(n_941),
.Y(n_1077)
);

NOR2x1p5_ASAP7_75t_L g1078 ( 
.A(n_1037),
.B(n_897),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1029),
.B(n_909),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_980),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_985),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1003),
.B(n_945),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_973),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1002),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_969),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_976),
.A2(n_1005),
.B1(n_962),
.B2(n_971),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_990),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_988),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1006),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_982),
.B(n_930),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_969),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_994),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_974),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1032),
.B(n_948),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_976),
.B(n_663),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_996),
.B(n_0),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_976),
.B(n_664),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1024),
.B(n_668),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_977),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1008),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_975),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1005),
.B(n_671),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_964),
.B(n_912),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_979),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1041),
.B(n_672),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_1005),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_1013),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_978),
.B(n_675),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_972),
.B(n_676),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1013),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_990),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_993),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1016),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_995),
.B(n_677),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_997),
.B(n_678),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_682),
.Y(n_1119)
);

AND2x2_ASAP7_75t_SL g1120 ( 
.A(n_1040),
.B(n_0),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1017),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_966),
.B(n_683),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1007),
.A2(n_687),
.B1(n_689),
.B2(n_684),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1011),
.Y(n_1124)
);

INVxp33_ASAP7_75t_L g1125 ( 
.A(n_992),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1014),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_1010),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1010),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1000),
.B(n_690),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_987),
.B(n_700),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_960),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_961),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1049),
.B(n_1051),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_987),
.A2(n_708),
.B1(n_709),
.B2(n_704),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1053),
.B(n_712),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_963),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_981),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1053),
.B(n_713),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1018),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_992),
.B(n_1),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_1004),
.B(n_716),
.C(n_714),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1021),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1023),
.B(n_1027),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1028),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_1025),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1035),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1036),
.B(n_2),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1019),
.A2(n_722),
.B1(n_723),
.B2(n_719),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1030),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1030),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1058),
.B(n_1022),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1062),
.B(n_1026),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1069),
.B(n_1034),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1097),
.B(n_1044),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1071),
.B(n_1046),
.Y(n_1158)
);

OAI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1123),
.A2(n_1050),
.B1(n_1048),
.B2(n_989),
.C(n_753),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1066),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1093),
.B(n_989),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1075),
.B(n_725),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1060),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1093),
.B(n_726),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1065),
.A2(n_729),
.B1(n_730),
.B2(n_728),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1088),
.B(n_2),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1056),
.B(n_733),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1090),
.A2(n_739),
.B1(n_743),
.B2(n_737),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1092),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1111),
.B(n_748),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1076),
.B(n_3),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1076),
.B(n_752),
.C(n_751),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1151),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_1057),
.B(n_756),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1080),
.B(n_1094),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1100),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1129),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1089),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1064),
.B(n_759),
.C(n_757),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1063),
.B(n_761),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_771),
.B(n_772),
.C(n_766),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1105),
.B(n_4),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1120),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1106),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1115),
.B(n_5),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_1061),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1116),
.B(n_7),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1101),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1059),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1077),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1121),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1142),
.B(n_8),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1055),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1124),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1127),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1086),
.B(n_10),
.Y(n_1197)
);

AO22x2_ASAP7_75t_L g1198 ( 
.A1(n_1110),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1108),
.B(n_11),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1078),
.B2(n_1117),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1082),
.B(n_12),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1113),
.B(n_13),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1127),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1126),
.Y(n_1204)
);

BUFx5_ASAP7_75t_L g1205 ( 
.A(n_1138),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1070),
.B(n_14),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1054),
.B(n_14),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1131),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1083),
.B(n_15),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1108),
.B(n_15),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1114),
.B(n_16),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1141),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1133),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1108),
.B(n_16),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1096),
.B(n_17),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1118),
.B(n_17),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1144),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1129),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1132),
.B(n_18),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1102),
.B(n_18),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_SL g1221 ( 
.A(n_1128),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1139),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1098),
.B(n_1134),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1074),
.B(n_19),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1074),
.B(n_20),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1146),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1081),
.B(n_22),
.Y(n_1227)
);

NOR2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1068),
.B(n_23),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1081),
.B(n_23),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1148),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1085),
.B(n_24),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1145),
.Y(n_1232)
);

AND2x2_ASAP7_75t_SL g1233 ( 
.A(n_1087),
.B(n_25),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1230),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1200),
.B(n_1087),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1153),
.B(n_1109),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1155),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1173),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1161),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1178),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1221),
.Y(n_1241)
);

NOR2x2_ASAP7_75t_L g1242 ( 
.A(n_1233),
.B(n_1125),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1232),
.B(n_1112),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1178),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1190),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1154),
.B(n_1128),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1175),
.B(n_1127),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1169),
.Y(n_1248)
);

BUFx8_ASAP7_75t_L g1249 ( 
.A(n_1207),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1160),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1218),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1177),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1157),
.A2(n_1067),
.B(n_1095),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1187),
.B(n_1152),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1218),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1193),
.A2(n_1103),
.B1(n_1136),
.B2(n_1072),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1176),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1185),
.B(n_1143),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1209),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1187),
.B(n_1152),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1189),
.A2(n_1140),
.B1(n_1137),
.B2(n_1149),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_L g1262 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1203),
.B(n_1104),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1163),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1192),
.B(n_1119),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1216),
.B(n_1171),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1212),
.B(n_1130),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1220),
.Y(n_1268)
);

NOR2x2_ASAP7_75t_L g1269 ( 
.A(n_1228),
.B(n_1147),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1217),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1226),
.B(n_1147),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1179),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1227),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1166),
.B(n_1147),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1211),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1202),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1224),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1164),
.B(n_1122),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1225),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1208),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_SL g1281 ( 
.A(n_1184),
.B(n_1150),
.C(n_1135),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1198),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1194),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1229),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1172),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1206),
.B(n_1079),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1231),
.Y(n_1287)
);

INVx5_ASAP7_75t_L g1288 ( 
.A(n_1204),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1213),
.Y(n_1289)
);

BUFx4f_ASAP7_75t_L g1290 ( 
.A(n_1195),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1191),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1219),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1292)
);

NOR2x2_ASAP7_75t_L g1293 ( 
.A(n_1198),
.B(n_26),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1174),
.B(n_27),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1158),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1183),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1205),
.B(n_1170),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1162),
.B(n_28),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1214),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1188),
.Y(n_1300)
);

AND2x6_ASAP7_75t_L g1301 ( 
.A(n_1186),
.B(n_137),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1167),
.B(n_29),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1156),
.B(n_30),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1205),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1205),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1182),
.B(n_1223),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1197),
.B(n_1181),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_SL g1308 ( 
.A(n_1222),
.B(n_38),
.C(n_30),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1215),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1205),
.B(n_31),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1165),
.B(n_31),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1201),
.B(n_32),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1234),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1239),
.A2(n_1199),
.B1(n_1210),
.B2(n_1159),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1259),
.B(n_1180),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1244),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1244),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1243),
.B(n_1168),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1248),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1244),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1241),
.B(n_32),
.Y(n_1321)
);

NAND2x1_ASAP7_75t_L g1322 ( 
.A(n_1304),
.B(n_138),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1257),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1245),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1236),
.B(n_33),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1245),
.B(n_33),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1270),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1238),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1264),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1235),
.B(n_34),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1280),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1250),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1287),
.B(n_35),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1252),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1249),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1268),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1283),
.Y(n_1337)
);

OR2x2_ASAP7_75t_SL g1338 ( 
.A(n_1276),
.B(n_35),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1272),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1295),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1289),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1240),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1240),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1273),
.B(n_1237),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1275),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1251),
.B(n_139),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1288),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1255),
.B(n_140),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1291),
.B(n_36),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1288),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1258),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1246),
.B(n_37),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1266),
.B(n_39),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1288),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1247),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1255),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1263),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1290),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1300),
.B(n_1267),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1285),
.B(n_39),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1277),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1254),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1299),
.B(n_40),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1296),
.B(n_40),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1284),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1265),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_L g1367 ( 
.A(n_1292),
.B(n_41),
.C(n_42),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1286),
.B(n_41),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_42),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1278),
.B(n_43),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_1302),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1294),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1309),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1271),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1303),
.B(n_43),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1282),
.B(n_44),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1302),
.B(n_44),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1260),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1262),
.B(n_46),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1298),
.B(n_48),
.Y(n_1381)
);

AND2x6_ASAP7_75t_L g1382 ( 
.A(n_1305),
.B(n_141),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1274),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1311),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1312),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1310),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1261),
.B(n_1297),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1328),
.B(n_48),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1340),
.A2(n_1253),
.A3(n_1301),
.B(n_1281),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1359),
.B(n_1256),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1358),
.B(n_1269),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1313),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1367),
.A2(n_1308),
.B(n_1301),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1370),
.A2(n_1301),
.B(n_1293),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1325),
.A2(n_49),
.B(n_50),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1378),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1386),
.A2(n_146),
.B(n_144),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1330),
.B(n_51),
.Y(n_1399)
);

AOI221x1_ASAP7_75t_L g1400 ( 
.A1(n_1351),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1322),
.A2(n_1387),
.B(n_1373),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1366),
.B(n_53),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1319),
.A2(n_151),
.B(n_147),
.Y(n_1403)
);

AO21x1_ASAP7_75t_L g1404 ( 
.A1(n_1355),
.A2(n_55),
.B(n_56),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_SL g1405 ( 
.A(n_1320),
.Y(n_1405)
);

AO21x1_ASAP7_75t_L g1406 ( 
.A1(n_1381),
.A2(n_56),
.B(n_57),
.Y(n_1406)
);

AOI31xp67_ASAP7_75t_L g1407 ( 
.A1(n_1388),
.A2(n_153),
.A3(n_155),
.B(n_152),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1384),
.B(n_57),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1318),
.B(n_58),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1382),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1314),
.A2(n_1353),
.B(n_1385),
.C(n_1352),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1374),
.A2(n_58),
.B(n_59),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1368),
.A2(n_1339),
.B(n_1347),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1334),
.Y(n_1414)
);

AOI211x1_ASAP7_75t_L g1415 ( 
.A1(n_1363),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1365),
.B(n_1336),
.Y(n_1416)
);

AO21x1_ASAP7_75t_L g1417 ( 
.A1(n_1376),
.A2(n_60),
.B(n_61),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1360),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1323),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1332),
.A2(n_1337),
.A3(n_1327),
.B(n_1331),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1329),
.A2(n_157),
.B(n_156),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1315),
.A2(n_64),
.B(n_66),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1324),
.B(n_66),
.Y(n_1423)
);

AOI211x1_ASAP7_75t_L g1424 ( 
.A1(n_1375),
.A2(n_1364),
.B(n_1349),
.C(n_1369),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1378),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1350),
.A2(n_1354),
.A3(n_1341),
.B(n_1377),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1333),
.B(n_1345),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1383),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1326),
.A2(n_1361),
.B1(n_1344),
.B2(n_1321),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1357),
.B(n_68),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1316),
.B(n_69),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1317),
.B(n_70),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1379),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1380),
.A2(n_70),
.B(n_71),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1382),
.A2(n_162),
.B(n_159),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1346),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1342),
.Y(n_1437)
);

O2A1O1Ixp5_ASAP7_75t_L g1438 ( 
.A1(n_1348),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1344),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1362),
.Y(n_1440)
);

AOI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1326),
.A2(n_164),
.B(n_163),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1382),
.A2(n_76),
.B(n_77),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1321),
.B(n_76),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_L g1444 ( 
.A1(n_1362),
.A2(n_1338),
.B1(n_1343),
.B2(n_1356),
.C(n_1342),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1343),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1356),
.Y(n_1446)
);

AOI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1372),
.A2(n_166),
.B(n_165),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1371),
.A2(n_77),
.B(n_78),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1335),
.A2(n_78),
.B(n_79),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1386),
.A2(n_168),
.B(n_167),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1386),
.A2(n_172),
.B(n_169),
.Y(n_1451)
);

NOR4xp25_ASAP7_75t_L g1452 ( 
.A(n_1351),
.B(n_81),
.C(n_79),
.D(n_80),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1359),
.B(n_80),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1365),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1386),
.A2(n_81),
.B(n_82),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_L g1456 ( 
.A(n_1325),
.B(n_83),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1386),
.A2(n_176),
.B(n_174),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1386),
.A2(n_178),
.B(n_177),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1324),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1367),
.A2(n_83),
.B(n_84),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1340),
.A2(n_186),
.A3(n_188),
.B(n_185),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1328),
.B(n_84),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1358),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1335),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1386),
.A2(n_85),
.B(n_86),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1349),
.B(n_85),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1330),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_1467)
);

INVx4_ASAP7_75t_SL g1468 ( 
.A(n_1378),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1319),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1386),
.A2(n_191),
.B(n_189),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1386),
.A2(n_196),
.B(n_194),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1349),
.B(n_87),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1313),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1367),
.A2(n_89),
.B(n_90),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1358),
.B(n_89),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1386),
.A2(n_199),
.B(n_198),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1386),
.A2(n_90),
.B(n_92),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1359),
.B(n_92),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1386),
.A2(n_93),
.B(n_94),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1342),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1325),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1359),
.B(n_96),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1358),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1367),
.A2(n_96),
.B(n_97),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1349),
.B(n_97),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1359),
.B(n_98),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1386),
.A2(n_203),
.B(n_201),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1325),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_L g1489 ( 
.A(n_1427),
.B(n_99),
.Y(n_1489)
);

BUFx2_ASAP7_75t_R g1490 ( 
.A(n_1464),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1459),
.B(n_100),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1410),
.A2(n_101),
.B(n_102),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1391),
.B(n_101),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1401),
.A2(n_102),
.B(n_103),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1405),
.Y(n_1495)
);

INVx3_ASAP7_75t_R g1496 ( 
.A(n_1475),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1480),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1466),
.B(n_103),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1420),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1410),
.A2(n_104),
.B(n_105),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1399),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1467),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1420),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1413),
.A2(n_596),
.B(n_205),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1410),
.B(n_204),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1439),
.B(n_206),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1468),
.B(n_207),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1419),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1454),
.B(n_109),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1423),
.B(n_110),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_110),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1437),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1411),
.B(n_111),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1442),
.A2(n_1394),
.B(n_1456),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1446),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1395),
.A2(n_114),
.B1(n_111),
.B2(n_112),
.C(n_115),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1424),
.B(n_112),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1396),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1392),
.B(n_208),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_SL g1523 ( 
.A1(n_1422),
.A2(n_119),
.B(n_120),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1428),
.B(n_119),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1460),
.A2(n_120),
.B(n_121),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1463),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1474),
.A2(n_122),
.B(n_123),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1483),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1403),
.A2(n_210),
.B(n_209),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1468),
.B(n_211),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1414),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1426),
.Y(n_1532)
);

AND2x6_ASAP7_75t_L g1533 ( 
.A(n_1429),
.B(n_212),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1473),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1453),
.B(n_122),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1426),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1440),
.B(n_213),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1444),
.B(n_214),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1416),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1445),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1433),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1430),
.Y(n_1542)
);

OAI22x1_ASAP7_75t_L g1543 ( 
.A1(n_1443),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_SL g1544 ( 
.A1(n_1417),
.A2(n_124),
.B(n_125),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1431),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1432),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1478),
.B(n_126),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1441),
.B(n_215),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1482),
.B(n_126),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1484),
.A2(n_127),
.B(n_128),
.Y(n_1550)
);

CKINVDCx11_ASAP7_75t_R g1551 ( 
.A(n_1397),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1447),
.B(n_216),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1402),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1408),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1485),
.B(n_217),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1435),
.B(n_1409),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1418),
.B(n_128),
.C(n_129),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1486),
.B(n_130),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1389),
.B(n_130),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1412),
.A2(n_131),
.B(n_132),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1476),
.A2(n_1436),
.B(n_1404),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1461),
.B(n_218),
.Y(n_1562)
);

NOR2xp67_ASAP7_75t_L g1563 ( 
.A(n_1455),
.B(n_131),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1465),
.A2(n_132),
.B(n_133),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1390),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1390),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1461),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1477),
.B(n_133),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1462),
.B(n_134),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1421),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1452),
.B(n_219),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1434),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1398),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1450),
.Y(n_1574)
);

AO21x1_ASAP7_75t_L g1575 ( 
.A1(n_1481),
.A2(n_134),
.B(n_135),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1479),
.A2(n_135),
.B(n_136),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1400),
.B(n_220),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1406),
.B(n_136),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1425),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1451),
.A2(n_224),
.B(n_225),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1415),
.Y(n_1581)
);

OAI21xp33_ASAP7_75t_L g1582 ( 
.A1(n_1488),
.A2(n_226),
.B(n_227),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1448),
.B(n_229),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1449),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1457),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1517),
.A2(n_1438),
.B(n_1470),
.C(n_1458),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1539),
.B(n_1509),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1539),
.B(n_1471),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1561),
.A2(n_1487),
.B(n_1407),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1514),
.Y(n_1590)
);

O2A1O1Ixp5_ASAP7_75t_L g1591 ( 
.A1(n_1575),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_R g1592 ( 
.A(n_1515),
.B(n_236),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1495),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1516),
.A2(n_237),
.B(n_238),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1582),
.A2(n_239),
.B(n_242),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1528),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1571),
.A2(n_244),
.B(n_245),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1508),
.B(n_246),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1541),
.B(n_247),
.Y(n_1599)
);

O2A1O1Ixp5_ASAP7_75t_L g1600 ( 
.A1(n_1501),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_1600)
);

CKINVDCx8_ASAP7_75t_R g1601 ( 
.A(n_1526),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1545),
.B(n_595),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1497),
.B(n_251),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1556),
.B(n_256),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1554),
.B(n_1546),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1542),
.B(n_257),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1567),
.Y(n_1607)
);

NOR2x2_ASAP7_75t_L g1608 ( 
.A(n_1522),
.B(n_258),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1540),
.B(n_1493),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1553),
.B(n_260),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1531),
.Y(n_1611)
);

BUFx2_ASAP7_75t_SL g1612 ( 
.A(n_1526),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1525),
.A2(n_261),
.B(n_262),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1518),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1519),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1491),
.B(n_269),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1521),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1498),
.B(n_273),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1499),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1565),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1513),
.B(n_594),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1532),
.B(n_274),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1527),
.A2(n_275),
.B(n_276),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1511),
.B(n_279),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1512),
.B(n_280),
.Y(n_1625)
);

NOR2xp67_ASAP7_75t_L g1626 ( 
.A(n_1535),
.B(n_281),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1502),
.A2(n_1550),
.B(n_1520),
.C(n_1569),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1489),
.B(n_282),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1578),
.B(n_593),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1490),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1503),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1559),
.B(n_283),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1534),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1536),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1547),
.B(n_592),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1548),
.A2(n_284),
.B(n_286),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1524),
.Y(n_1638)
);

INVx3_ASAP7_75t_SL g1639 ( 
.A(n_1522),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1494),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1566),
.B(n_1507),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1506),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1585),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1496),
.B(n_287),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1530),
.B(n_288),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1551),
.B(n_289),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1537),
.B(n_290),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1573),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1572),
.B(n_291),
.Y(n_1649)
);

BUFx10_ASAP7_75t_L g1650 ( 
.A(n_1533),
.Y(n_1650)
);

NAND2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1538),
.B(n_292),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1533),
.B(n_293),
.Y(n_1652)
);

XNOR2xp5_ASAP7_75t_L g1653 ( 
.A(n_1543),
.B(n_1549),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_SL g1654 ( 
.A(n_1533),
.B(n_294),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1558),
.B(n_295),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1583),
.B(n_1557),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1570),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1581),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_SL g1659 ( 
.A(n_1505),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1577),
.B(n_591),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1574),
.B(n_1548),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1580),
.A2(n_297),
.B(n_298),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1560),
.A2(n_1570),
.B(n_1500),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1562),
.B(n_300),
.Y(n_1664)
);

INVx3_ASAP7_75t_SL g1665 ( 
.A(n_1552),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1504),
.B(n_301),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1584),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1492),
.B(n_590),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1563),
.B(n_305),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1568),
.B(n_306),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1564),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1544),
.Y(n_1672)
);

OAI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1576),
.A2(n_1579),
.B(n_1523),
.C(n_1529),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1565),
.A2(n_310),
.B(n_311),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1509),
.B(n_589),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1509),
.B(n_313),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1539),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1517),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1539),
.B(n_317),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1539),
.B(n_588),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1509),
.B(n_318),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1509),
.B(n_319),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1517),
.A2(n_320),
.B(n_321),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1509),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1514),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1509),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1501),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1517),
.A2(n_326),
.B(n_327),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1539),
.B(n_587),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1509),
.B(n_328),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1509),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1515),
.Y(n_1692)
);

BUFx4_ASAP7_75t_R g1693 ( 
.A(n_1542),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1526),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_SL g1695 ( 
.A(n_1490),
.B(n_329),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1509),
.B(n_330),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1509),
.B(n_586),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1509),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1509),
.B(n_331),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1539),
.B(n_585),
.Y(n_1700)
);

OA21x2_ASAP7_75t_L g1701 ( 
.A1(n_1565),
.A2(n_332),
.B(n_335),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1518),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1501),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1684),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1590),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1614),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1654),
.A2(n_1656),
.B(n_1663),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1587),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1611),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1634),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_339),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1619),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1601),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1641),
.B(n_340),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1691),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1698),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1609),
.B(n_341),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1632),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1605),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1658),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1685),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1635),
.Y(n_1722)
);

AO31x2_ASAP7_75t_L g1723 ( 
.A1(n_1640),
.A2(n_347),
.A3(n_343),
.B(n_345),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1639),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1643),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1694),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1648),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1607),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1589),
.A2(n_348),
.B(n_349),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1653),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1657),
.Y(n_1732)
);

OR2x6_ASAP7_75t_L g1733 ( 
.A(n_1612),
.B(n_357),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1620),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1638),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1665),
.B(n_358),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1677),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1641),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1661),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1588),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1676),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1682),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1696),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1650),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1675),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1659),
.A2(n_362),
.B1(n_359),
.B2(n_361),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1702),
.B(n_363),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1681),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1690),
.A2(n_365),
.B(n_366),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1693),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1596),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1697),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1622),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1699),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1628),
.B(n_367),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1642),
.B(n_369),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1672),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1631),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1674),
.A2(n_1701),
.B(n_1666),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1593),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1600),
.A2(n_370),
.B(n_371),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1622),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1624),
.B(n_372),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1599),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1598),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1652),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1674),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1646),
.B(n_376),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1701),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1610),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1606),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1627),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1602),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1630),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1618),
.B(n_377),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1679),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1621),
.B(n_379),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1680),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1586),
.A2(n_380),
.B(n_383),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1592),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1689),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1700),
.Y(n_1782)
);

CKINVDCx8_ASAP7_75t_R g1783 ( 
.A(n_1713),
.Y(n_1783)
);

NOR2xp67_ASAP7_75t_SL g1784 ( 
.A(n_1713),
.B(n_1688),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1720),
.B(n_1616),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1739),
.B(n_1633),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1649),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1728),
.B(n_1695),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1712),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1724),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1772),
.A2(n_1615),
.B1(n_1660),
.B2(n_1629),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1772),
.A2(n_1626),
.B1(n_1664),
.B2(n_1623),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1719),
.B(n_1655),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1758),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1712),
.Y(n_1795)
);

AO21x2_ASAP7_75t_L g1796 ( 
.A1(n_1769),
.A2(n_1604),
.B(n_1636),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1769),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1713),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1726),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1727),
.B(n_1651),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1727),
.B(n_1708),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1729),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1718),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1722),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1734),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1737),
.B(n_1644),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1738),
.B(n_1664),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1735),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1752),
.B(n_1645),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1724),
.B(n_1645),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1750),
.B(n_1625),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1745),
.B(n_1594),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1740),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1780),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1745),
.B(n_1673),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1757),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1725),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1705),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1744),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1709),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1741),
.B(n_1603),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1748),
.B(n_1647),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1754),
.B(n_1591),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1704),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1710),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1744),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1762),
.B(n_1637),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1721),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1774),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1715),
.B(n_1597),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1759),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1716),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1774),
.B(n_1613),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1742),
.B(n_1668),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1732),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1743),
.B(n_1683),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1744),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1751),
.B(n_1678),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1707),
.A2(n_1595),
.B1(n_1670),
.B2(n_1669),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1764),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1765),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1760),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1706),
.B(n_1667),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1760),
.B(n_1662),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1770),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1753),
.B(n_1671),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1778),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1711),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1771),
.B(n_1617),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1779),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1789),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1794),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1795),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1804),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1804),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1801),
.B(n_1773),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1797),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1797),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1843),
.B(n_1778),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1830),
.B(n_1736),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1839),
.Y(n_1864)
);

NOR4xp25_ASAP7_75t_SL g1865 ( 
.A(n_1820),
.B(n_1608),
.C(n_1782),
.D(n_1733),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1830),
.B(n_1782),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1810),
.B(n_1776),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1790),
.B(n_1781),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1827),
.B(n_1786),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1794),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1827),
.B(n_1755),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1817),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1817),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1803),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1827),
.B(n_1768),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1832),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1802),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1802),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1803),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1806),
.B(n_1779),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1832),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1851),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1849),
.B(n_1775),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1806),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1836),
.Y(n_1885)
);

AOI222xp33_ASAP7_75t_L g1886 ( 
.A1(n_1791),
.A2(n_1731),
.B1(n_1761),
.B2(n_1746),
.C1(n_1717),
.C2(n_1777),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1849),
.B(n_1733),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1838),
.B(n_1747),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1798),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1836),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1828),
.B(n_1756),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1805),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1889),
.B(n_1838),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1852),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1854),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1882),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1869),
.B(n_1860),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1864),
.B(n_1816),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1860),
.B(n_1811),
.Y(n_1899)
);

NOR2xp67_ASAP7_75t_L g1900 ( 
.A(n_1870),
.B(n_1851),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1861),
.B(n_1798),
.Y(n_1901)
);

AOI21xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1861),
.A2(n_1844),
.B(n_1845),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1883),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1866),
.Y(n_1904)
);

AND2x2_ASAP7_75t_SL g1905 ( 
.A(n_1887),
.B(n_1812),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1882),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1866),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1887),
.Y(n_1908)
);

NOR2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1853),
.B(n_1818),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1863),
.B(n_1824),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1853),
.B(n_1818),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1872),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1892),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1863),
.B(n_1831),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1864),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1891),
.B(n_1788),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1873),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1877),
.Y(n_1918)
);

OR2x6_ASAP7_75t_L g1919 ( 
.A(n_1891),
.B(n_1763),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1892),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1878),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1876),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1884),
.B(n_1834),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1875),
.B(n_1831),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1862),
.B(n_1828),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1868),
.B(n_1828),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1880),
.B(n_1809),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1871),
.B(n_1800),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1894),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1898),
.A2(n_1886),
.B1(n_1881),
.B2(n_1791),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1916),
.Y(n_1931)
);

OAI211xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1908),
.A2(n_1896),
.B(n_1906),
.C(n_1915),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1909),
.B(n_1865),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1919),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1894),
.Y(n_1935)
);

OAI33xp33_ASAP7_75t_L g1936 ( 
.A1(n_1896),
.A2(n_1880),
.A3(n_1793),
.B1(n_1813),
.B2(n_1855),
.B3(n_1856),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1895),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1901),
.B(n_1865),
.Y(n_1938)
);

AO21x2_ASAP7_75t_L g1939 ( 
.A1(n_1906),
.A2(n_1859),
.B(n_1858),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1895),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1919),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1923),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1914),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1910),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1905),
.A2(n_1886),
.B1(n_1850),
.B2(n_1792),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1912),
.B(n_1799),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1917),
.B(n_1840),
.C(n_1792),
.Y(n_1947)
);

OAI33xp33_ASAP7_75t_L g1948 ( 
.A1(n_1917),
.A2(n_1785),
.A3(n_1841),
.B1(n_1842),
.B2(n_1825),
.B3(n_1833),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1911),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1918),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1931),
.B(n_1897),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1931),
.B(n_1899),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1940),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1929),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1929),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1939),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1935),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1944),
.B(n_1943),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1939),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1937),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1942),
.B(n_1893),
.Y(n_1961)
);

INVx2_ASAP7_75t_SL g1962 ( 
.A(n_1938),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1946),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1949),
.B(n_1903),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1934),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1947),
.B(n_1921),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1954),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1951),
.B(n_1932),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1961),
.B(n_1924),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1966),
.B(n_1950),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1964),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1952),
.B(n_1904),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1958),
.B(n_1907),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1962),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1955),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1965),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1963),
.B(n_1945),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1960),
.Y(n_1978)
);

OAI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1963),
.A2(n_1933),
.B(n_1930),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1953),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1960),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1953),
.B(n_1925),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1969),
.B(n_1925),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1976),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1974),
.B(n_1926),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1971),
.B(n_1974),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1979),
.A2(n_1936),
.B1(n_1959),
.B2(n_1956),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_SL g1988 ( 
.A(n_1979),
.B(n_1902),
.C(n_1783),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1970),
.Y(n_1989)
);

NOR4xp25_ASAP7_75t_L g1990 ( 
.A(n_1977),
.B(n_1957),
.C(n_1941),
.D(n_1927),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1968),
.A2(n_1948),
.B1(n_1922),
.B2(n_1900),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1973),
.B(n_1916),
.Y(n_1992)
);

AND2x2_ASAP7_75t_SL g1993 ( 
.A(n_1982),
.B(n_1926),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1980),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1989),
.B(n_1972),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1993),
.B(n_1967),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1986),
.A2(n_1981),
.B(n_1978),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1990),
.A2(n_1975),
.B1(n_1920),
.B2(n_1913),
.C(n_1840),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1994),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1984),
.B(n_1928),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1985),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1983),
.B(n_1857),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1992),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1990),
.B(n_1823),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1987),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_2002),
.B(n_1991),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1997),
.A2(n_1988),
.B(n_1859),
.Y(n_2007)
);

AOI211x1_ASAP7_75t_L g2008 ( 
.A1(n_2005),
.A2(n_1888),
.B(n_1784),
.C(n_1807),
.Y(n_2008)
);

AOI21xp33_ASAP7_75t_L g2009 ( 
.A1(n_1995),
.A2(n_1749),
.B(n_1858),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2001),
.B(n_1822),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_2004),
.A2(n_1783),
.B1(n_1879),
.B2(n_1874),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2000),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1996),
.A2(n_1796),
.B1(n_1837),
.B2(n_1847),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1998),
.B(n_1847),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_2003),
.B(n_1867),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_2012),
.B(n_1999),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_2006),
.B(n_1787),
.Y(n_2017)
);

INVxp67_ASAP7_75t_L g2018 ( 
.A(n_2007),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2010),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2008),
.B(n_1835),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_SL g2021 ( 
.A(n_2015),
.B(n_2014),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2011),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2013),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2009),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2010),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_2012),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2012),
.B(n_1848),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2012),
.B(n_1848),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2010),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_2012),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2012),
.B(n_1874),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2017),
.B(n_1879),
.Y(n_2032)
);

NOR4xp25_ASAP7_75t_SL g2033 ( 
.A(n_2022),
.B(n_1846),
.C(n_1766),
.D(n_1703),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2021),
.B(n_1847),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_2028),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_2016),
.B(n_1687),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2019),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2026),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2030),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2025),
.B(n_1796),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2029),
.B(n_1885),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2027),
.B(n_1890),
.Y(n_2042)
);

NOR2xp67_ASAP7_75t_L g2043 ( 
.A(n_2018),
.B(n_385),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2023),
.B(n_1805),
.Y(n_2044)
);

NOR3xp33_ASAP7_75t_SL g2045 ( 
.A(n_2031),
.B(n_1730),
.C(n_1723),
.Y(n_2045)
);

NAND5xp2_ASAP7_75t_L g2046 ( 
.A(n_2038),
.B(n_2024),
.C(n_2020),
.D(n_1808),
.E(n_1723),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_L g2047 ( 
.A(n_2039),
.B(n_1814),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_2034),
.B(n_1814),
.Y(n_2048)
);

NOR3xp33_ASAP7_75t_L g2049 ( 
.A(n_2037),
.B(n_1723),
.C(n_1819),
.Y(n_2049)
);

NAND4xp25_ASAP7_75t_L g2050 ( 
.A(n_2036),
.B(n_1821),
.C(n_1826),
.D(n_1819),
.Y(n_2050)
);

OAI21xp33_ASAP7_75t_L g2051 ( 
.A1(n_2040),
.A2(n_1826),
.B(n_1821),
.Y(n_2051)
);

OAI31xp33_ASAP7_75t_L g2052 ( 
.A1(n_2035),
.A2(n_2044),
.A3(n_2041),
.B(n_2032),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2043),
.B(n_1829),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_2042),
.B(n_2045),
.Y(n_2054)
);

NAND3xp33_ASAP7_75t_L g2055 ( 
.A(n_2033),
.B(n_1829),
.C(n_386),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2052),
.B(n_391),
.Y(n_2056)
);

AOI211xp5_ASAP7_75t_L g2057 ( 
.A1(n_2055),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2054),
.A2(n_584),
.B1(n_397),
.B2(n_395),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_SL g2059 ( 
.A(n_2049),
.B(n_396),
.C(n_398),
.Y(n_2059)
);

AOI211xp5_ASAP7_75t_L g2060 ( 
.A1(n_2046),
.A2(n_403),
.B(n_399),
.C(n_402),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_405),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_2047),
.B(n_408),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2048),
.B(n_409),
.Y(n_2063)
);

O2A1O1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_2053),
.A2(n_2051),
.B(n_415),
.C(n_411),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2047),
.Y(n_2065)
);

NAND4xp75_ASAP7_75t_L g2066 ( 
.A(n_2052),
.B(n_417),
.C(n_414),
.D(n_416),
.Y(n_2066)
);

NOR2x1_ASAP7_75t_L g2067 ( 
.A(n_2055),
.B(n_420),
.Y(n_2067)
);

NOR3xp33_ASAP7_75t_L g2068 ( 
.A(n_2056),
.B(n_422),
.C(n_424),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2066),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_2065),
.B(n_426),
.Y(n_2070)
);

OAI21xp33_ASAP7_75t_SL g2071 ( 
.A1(n_2067),
.A2(n_429),
.B(n_430),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2060),
.B(n_432),
.Y(n_2072)
);

NAND2xp33_ASAP7_75t_L g2073 ( 
.A(n_2063),
.B(n_433),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_2061),
.Y(n_2074)
);

XNOR2x2_ASAP7_75t_L g2075 ( 
.A(n_2058),
.B(n_434),
.Y(n_2075)
);

AOI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_2057),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_2076)
);

OAI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2062),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.C(n_441),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_2064),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2059),
.B(n_442),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_SL g2080 ( 
.A(n_2065),
.B(n_443),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2067),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2058),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2071),
.B(n_453),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_2080),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2078),
.B(n_455),
.Y(n_2085)
);

NOR3xp33_ASAP7_75t_L g2086 ( 
.A(n_2074),
.B(n_456),
.C(n_457),
.Y(n_2086)
);

OAI21xp33_ASAP7_75t_L g2087 ( 
.A1(n_2069),
.A2(n_458),
.B(n_459),
.Y(n_2087)
);

NOR2x1_ASAP7_75t_SL g2088 ( 
.A(n_2070),
.B(n_460),
.Y(n_2088)
);

NOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2072),
.B(n_461),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2079),
.B(n_462),
.Y(n_2090)
);

NAND2x1p5_ASAP7_75t_L g2091 ( 
.A(n_2081),
.B(n_464),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2073),
.Y(n_2092)
);

OAI211xp5_ASAP7_75t_L g2093 ( 
.A1(n_2076),
.A2(n_465),
.B(n_467),
.C(n_468),
.Y(n_2093)
);

NAND4xp75_ASAP7_75t_L g2094 ( 
.A(n_2075),
.B(n_469),
.C(n_470),
.D(n_471),
.Y(n_2094)
);

NOR3xp33_ASAP7_75t_SL g2095 ( 
.A(n_2077),
.B(n_472),
.C(n_473),
.Y(n_2095)
);

NOR3xp33_ASAP7_75t_SL g2096 ( 
.A(n_2082),
.B(n_2068),
.C(n_474),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2069),
.B(n_476),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2074),
.Y(n_2098)
);

NOR2x1_ASAP7_75t_L g2099 ( 
.A(n_2070),
.B(n_477),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2078),
.B(n_478),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2078),
.B(n_481),
.Y(n_2101)
);

AOI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2098),
.A2(n_482),
.B1(n_483),
.B2(n_486),
.C(n_489),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2101),
.Y(n_2103)
);

NOR2x1_ASAP7_75t_L g2104 ( 
.A(n_2094),
.B(n_490),
.Y(n_2104)
);

NAND3xp33_ASAP7_75t_SL g2105 ( 
.A(n_2086),
.B(n_2100),
.C(n_2085),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2092),
.Y(n_2106)
);

NOR3xp33_ASAP7_75t_L g2107 ( 
.A(n_2097),
.B(n_491),
.C(n_492),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2088),
.Y(n_2108)
);

AND2x2_ASAP7_75t_SL g2109 ( 
.A(n_2083),
.B(n_493),
.Y(n_2109)
);

OAI211xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2084),
.A2(n_496),
.B(n_497),
.C(n_498),
.Y(n_2110)
);

AOI321xp33_ASAP7_75t_L g2111 ( 
.A1(n_2089),
.A2(n_499),
.A3(n_500),
.B1(n_501),
.B2(n_502),
.C(n_503),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2087),
.A2(n_504),
.B(n_506),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2109),
.B(n_2108),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_2106),
.B(n_2099),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2104),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_2103),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2105),
.A2(n_2093),
.B1(n_2090),
.B2(n_2091),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2112),
.B(n_2095),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2111),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2107),
.B(n_2096),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2114),
.B(n_2102),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2113),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2119),
.Y(n_2123)
);

AOI21xp33_ASAP7_75t_L g2124 ( 
.A1(n_2116),
.A2(n_2110),
.B(n_508),
.Y(n_2124)
);

OAI211xp5_ASAP7_75t_L g2125 ( 
.A1(n_2122),
.A2(n_2115),
.B(n_2117),
.C(n_2118),
.Y(n_2125)
);

OAI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2123),
.A2(n_2120),
.B1(n_510),
.B2(n_514),
.C(n_515),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2126),
.Y(n_2127)
);

NAND3xp33_ASAP7_75t_SL g2128 ( 
.A(n_2125),
.B(n_2121),
.C(n_2124),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2128),
.Y(n_2129)
);

AOI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_2127),
.A2(n_509),
.B1(n_516),
.B2(n_518),
.Y(n_2130)
);

OAI322xp33_ASAP7_75t_L g2131 ( 
.A1(n_2129),
.A2(n_519),
.A3(n_520),
.B1(n_521),
.B2(n_522),
.C1(n_523),
.C2(n_524),
.Y(n_2131)
);

AOI211xp5_ASAP7_75t_L g2132 ( 
.A1(n_2130),
.A2(n_525),
.B(n_526),
.C(n_528),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2132),
.A2(n_529),
.B1(n_531),
.B2(n_532),
.Y(n_2133)
);

OAI22x1_ASAP7_75t_L g2134 ( 
.A1(n_2131),
.A2(n_583),
.B1(n_534),
.B2(n_535),
.Y(n_2134)
);

XNOR2xp5_ASAP7_75t_L g2135 ( 
.A(n_2134),
.B(n_533),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2133),
.A2(n_536),
.B1(n_538),
.B2(n_539),
.Y(n_2136)
);

OAI222xp33_ASAP7_75t_L g2137 ( 
.A1(n_2135),
.A2(n_542),
.B1(n_543),
.B2(n_544),
.C1(n_545),
.C2(n_546),
.Y(n_2137)
);

OAI211xp5_ASAP7_75t_L g2138 ( 
.A1(n_2136),
.A2(n_547),
.B(n_548),
.C(n_549),
.Y(n_2138)
);

XNOR2xp5_ASAP7_75t_L g2139 ( 
.A(n_2135),
.B(n_550),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2135),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2139),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2140),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2138),
.Y(n_2143)
);

INVxp67_ASAP7_75t_SL g2144 ( 
.A(n_2137),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2142),
.B(n_2141),
.Y(n_2145)
);

AOI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_2144),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.C(n_555),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_2143),
.B(n_556),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2145),
.A2(n_558),
.B(n_559),
.Y(n_2148)
);

AOI211xp5_ASAP7_75t_L g2149 ( 
.A1(n_2148),
.A2(n_2147),
.B(n_2146),
.C(n_563),
.Y(n_2149)
);


endmodule