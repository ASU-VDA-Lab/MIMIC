module fake_jpeg_2198_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_11),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_30),
.A2(n_37),
.B1(n_44),
.B2(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_39),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_6),
.B1(n_17),
.B2(n_29),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_19),
.B(n_37),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_6),
.B1(n_12),
.B2(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_25),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_54),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_23),
.C(n_28),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_51),
.B1(n_48),
.B2(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_71),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_32),
.A2(n_34),
.B(n_44),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_48),
.B(n_51),
.C(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_71),
.B1(n_48),
.B2(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_91),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_66),
.B1(n_52),
.B2(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_66),
.B1(n_73),
.B2(n_62),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_81),
.Y(n_101)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_69),
.C(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_87),
.B1(n_74),
.B2(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_85),
.B(n_79),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_85),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_89),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_86),
.B(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_105),
.C(n_96),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_93),
.B(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_97),
.B1(n_101),
.B2(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_107),
.B1(n_108),
.B2(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_109),
.C(n_112),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_115),
.B(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_119),
.B(n_117),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);


endmodule