module fake_jpeg_28553_n_246 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_52),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_33),
.B1(n_25),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_61),
.B1(n_70),
.B2(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_33),
.B1(n_25),
.B2(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_36),
.B1(n_23),
.B2(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_72),
.B1(n_81),
.B2(n_47),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_18),
.B1(n_34),
.B2(n_24),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_70),
.B1(n_54),
.B2(n_65),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_49),
.B1(n_51),
.B2(n_28),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_25),
.B1(n_35),
.B2(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_28),
.B1(n_31),
.B2(n_24),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_31),
.B1(n_18),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_21),
.B1(n_18),
.B2(n_47),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_68),
.C(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_86),
.A2(n_106),
.B1(n_19),
.B2(n_4),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_34),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_43),
.B(n_1),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_99),
.B1(n_66),
.B2(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_102),
.B1(n_66),
.B2(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_21),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_67),
.B(n_77),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_46),
.B(n_19),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_56),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_13),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_139),
.B1(n_93),
.B2(n_97),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_123),
.B1(n_131),
.B2(n_109),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_135),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_87),
.B(n_92),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_152),
.B(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_85),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_85),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_160),
.B(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_90),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_89),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_88),
.C(n_103),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_127),
.C(n_129),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_87),
.B(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_102),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_161),
.B1(n_121),
.B2(n_130),
.C(n_97),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_125),
.A2(n_97),
.B1(n_110),
.B2(n_113),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_137),
.B1(n_105),
.B2(n_5),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_152),
.B(n_162),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_166),
.B(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_174),
.B1(n_182),
.B2(n_160),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_133),
.B(n_138),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_132),
.B(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_180),
.C(n_143),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_137),
.B(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_145),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_175),
.B(n_146),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_0),
.B(n_4),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_19),
.C(n_9),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_196),
.B(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_189),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_151),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_197),
.C(n_199),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_145),
.B1(n_156),
.B2(n_151),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_179),
.B(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_143),
.C(n_160),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_163),
.B(n_19),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_192),
.B(n_186),
.Y(n_221)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_172),
.C(n_166),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_170),
.C(n_176),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_192),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_185),
.B(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_221),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_208),
.C(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_228),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_230),
.C(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_204),
.C(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_224),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_201),
.B1(n_219),
.B2(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_174),
.B1(n_202),
.B2(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_182),
.Y(n_242)
);

OAI321xp33_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_216),
.A3(n_200),
.B1(n_210),
.B2(n_183),
.C(n_222),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_231),
.C(n_227),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_242),
.B(n_13),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_236),
.B(n_180),
.Y(n_243)
);

AOI321xp33_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.A3(n_6),
.B1(n_8),
.B2(n_163),
.C(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_6),
.Y(n_246)
);


endmodule