module fake_jpeg_24278_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_26),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_53),
.B(n_63),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_30),
.C(n_34),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_17),
.C(n_33),
.Y(n_90)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_72),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_67),
.Y(n_113)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_40),
.B1(n_56),
.B2(n_32),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_18),
.Y(n_115)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_29),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_31),
.B1(n_30),
.B2(n_17),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_31),
.B1(n_37),
.B2(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_92),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_49),
.B1(n_43),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_106),
.B1(n_110),
.B2(n_19),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_65),
.B(n_72),
.C(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_118),
.B1(n_0),
.B2(n_1),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_94),
.C(n_27),
.Y(n_144)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_34),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_105),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_66),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_102),
.B(n_67),
.C(n_66),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_23),
.B1(n_17),
.B2(n_18),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_111),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_43),
.B1(n_39),
.B2(n_32),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_102),
.B1(n_23),
.B2(n_38),
.Y(n_130)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_126),
.C(n_144),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_73),
.B(n_37),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_129),
.B(n_134),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_41),
.A3(n_45),
.B1(n_74),
.B2(n_19),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_131),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_45),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_127),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_51),
.B(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_154),
.B1(n_89),
.B2(n_98),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_74),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_137),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_64),
.B1(n_51),
.B2(n_41),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_145),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_67),
.B(n_29),
.C(n_36),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_103),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_38),
.B1(n_27),
.B2(n_24),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_41),
.B1(n_24),
.B2(n_21),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_67),
.C(n_28),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_113),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_156),
.B(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_158),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_124),
.B1(n_141),
.B2(n_122),
.Y(n_197)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_82),
.B1(n_117),
.B2(n_114),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_165),
.A2(n_168),
.B1(n_170),
.B2(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_169),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_97),
.B1(n_116),
.B2(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_179),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_175),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_111),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_104),
.B1(n_87),
.B2(n_97),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_184),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_87),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_187),
.B1(n_8),
.B2(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_101),
.B(n_2),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_125),
.B(n_3),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_123),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_121),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_189),
.B(n_10),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_151),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_126),
.A3(n_145),
.B1(n_143),
.B2(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_161),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_143),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_201),
.B(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_177),
.B1(n_169),
.B2(n_165),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_149),
.B(n_128),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_215),
.B(n_184),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_203),
.Y(n_219)
);

OR2x4_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_1),
.C(n_5),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_5),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_96),
.C(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_210),
.C(n_178),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_96),
.Y(n_210)
);

CKINVDCx12_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_214),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_10),
.B(n_11),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_10),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_243),
.C(n_208),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_229),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_228),
.B(n_236),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_239),
.B1(n_213),
.B2(n_198),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_193),
.B(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_180),
.B1(n_162),
.B2(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_196),
.B1(n_191),
.B2(n_206),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_157),
.B1(n_187),
.B2(n_163),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_188),
.B1(n_202),
.B2(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_192),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_161),
.B1(n_156),
.B2(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

HAxp5_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_192),
.CON(n_247),
.SN(n_247)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_250),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_195),
.C(n_205),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_259),
.Y(n_270)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_235),
.C(n_228),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_190),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_262),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_219),
.B(n_209),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_199),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_206),
.Y(n_281)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_215),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_198),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_237),
.Y(n_275)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_272),
.C(n_277),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_226),
.B(n_229),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_11),
.B(n_12),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_226),
.C(n_222),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_231),
.B1(n_232),
.B2(n_237),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_250),
.B1(n_248),
.B2(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_240),
.C(n_224),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_224),
.C(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_253),
.B(n_244),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_292),
.B(n_268),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_277),
.C(n_280),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_261),
.B1(n_257),
.B2(n_249),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_291),
.B1(n_293),
.B2(n_295),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_245),
.B(n_242),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_247),
.B1(n_171),
.B2(n_15),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_300),
.B(n_303),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_270),
.B1(n_265),
.B2(n_272),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_290),
.B1(n_294),
.B2(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_271),
.C(n_274),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_276),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_312),
.C(n_15),
.Y(n_316)
);

OAI21x1_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_295),
.B(n_287),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_305),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_284),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_308),
.B(n_307),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_15),
.B1(n_16),
.B2(n_297),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_304),
.B(n_302),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_16),
.C(n_313),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_315),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_311),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_318),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.Y(n_327)
);


endmodule