module fake_jpeg_21349_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_28),
.B1(n_15),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_8),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_16),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_10),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_14),
.B(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_46),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_64),
.Y(n_65)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_11),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_39),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_62),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_36),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_56),
.B1(n_55),
.B2(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_62),
.B1(n_49),
.B2(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_75),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_65),
.C(n_73),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.C(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_65),
.C(n_69),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_67),
.B(n_74),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_79),
.B(n_76),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_89),
.B(n_92),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_54),
.B1(n_53),
.B2(n_37),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_59),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_64),
.B(n_70),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_70),
.C(n_63),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_59),
.C(n_37),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_11),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_100),
.Y(n_102)
);


endmodule