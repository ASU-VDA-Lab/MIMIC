module fake_netlist_1_1057_n_11 (n_3, n_1, n_2, n_0, n_11);
input n_3;
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
OAI22xp33_ASAP7_75t_L g4 ( .A1(n_2), .A2(n_1), .B1(n_0), .B2(n_3), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_2), .B(n_0), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_1), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_5), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
NOR2x1_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .Y(n_10) );
XOR2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .Y(n_11) );
endmodule