module fake_jpeg_13005_n_132 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_12),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_67),
.B1(n_71),
.B2(n_42),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_17),
.B(n_22),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_41),
.B1(n_46),
.B2(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_11),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_12),
.B1(n_38),
.B2(n_31),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_61),
.B1(n_53),
.B2(n_63),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_5),
.B1(n_8),
.B2(n_48),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_81),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.C(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_68),
.C(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_90),
.B(n_63),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_61),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_101),
.B1(n_82),
.B2(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_51),
.B1(n_86),
.B2(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_90),
.B(n_83),
.C(n_88),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_104),
.B1(n_94),
.B2(n_102),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_123),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_112),
.B1(n_110),
.B2(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_123),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_121),
.C(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_125),
.A3(n_124),
.B1(n_110),
.B2(n_100),
.C1(n_93),
.C2(n_98),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_100),
.C(n_93),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_93),
.Y(n_132)
);


endmodule