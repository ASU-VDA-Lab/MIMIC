module fake_jpeg_31729_n_527 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_52),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_54),
.Y(n_159)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_16),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_59),
.Y(n_134)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_15),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_66),
.B(n_68),
.Y(n_166)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_15),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_89),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_28),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_103),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_28),
.B(n_14),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_29),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_45),
.B1(n_35),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_115),
.A2(n_123),
.B1(n_130),
.B2(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_80),
.B1(n_54),
.B2(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_128),
.B1(n_158),
.B2(n_38),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_52),
.A2(n_45),
.B1(n_46),
.B2(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_151),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_10),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_161),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_56),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_29),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_82),
.A2(n_42),
.B1(n_43),
.B2(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_36),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_75),
.A2(n_42),
.B1(n_17),
.B2(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_62),
.B(n_19),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_31),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_61),
.A2(n_22),
.B1(n_39),
.B2(n_17),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_22),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_170),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_106),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_110),
.B(n_38),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_192),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_78),
.B1(n_79),
.B2(n_100),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_180),
.A2(n_197),
.B1(n_209),
.B2(n_148),
.Y(n_249)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_181),
.Y(n_222)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_183),
.Y(n_225)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_188),
.B(n_205),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_18),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_193),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_106),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_18),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_155),
.B(n_95),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_109),
.A2(n_105),
.B1(n_102),
.B2(n_104),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_203),
.B1(n_213),
.B2(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_144),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_201),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_134),
.B(n_93),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_84),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_204),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_101),
.B1(n_86),
.B2(n_87),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_96),
.B1(n_92),
.B2(n_91),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_162),
.B(n_98),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_141),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_152),
.A2(n_16),
.B1(n_32),
.B2(n_24),
.Y(n_215)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_217),
.B1(n_134),
.B2(n_117),
.Y(n_247)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_113),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_229),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_114),
.C(n_120),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_215),
.C(n_77),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_138),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_212),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_214),
.B1(n_190),
.B2(n_168),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_167),
.B1(n_107),
.B2(n_131),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_112),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_253),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_189),
.B(n_147),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_193),
.B(n_122),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_212),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_182),
.B(n_196),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_275),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_183),
.B(n_181),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_286),
.B(n_230),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_172),
.B1(n_180),
.B2(n_112),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_267),
.B1(n_271),
.B2(n_273),
.Y(n_296)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_276),
.B(n_225),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_223),
.B(n_177),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_270),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_268),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_285),
.C(n_220),
.Y(n_306)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_251),
.B1(n_252),
.B2(n_249),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_253),
.B1(n_254),
.B2(n_248),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_185),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_153),
.B1(n_195),
.B2(n_164),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_252),
.B1(n_245),
.B2(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_153),
.B1(n_164),
.B2(n_149),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_216),
.B1(n_117),
.B2(n_204),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_209),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g276 ( 
.A(n_222),
.B(n_206),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_171),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_71),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_281),
.Y(n_309)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_208),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_239),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_243),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_218),
.B(n_217),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_218),
.B(n_210),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_228),
.B(n_106),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_233),
.A2(n_186),
.B1(n_187),
.B2(n_191),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_316),
.B1(n_271),
.B2(n_274),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_221),
.A3(n_248),
.B1(n_237),
.B2(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_291),
.B(n_297),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_225),
.B(n_222),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_292),
.A2(n_308),
.B(n_311),
.C(n_265),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_267),
.A2(n_221),
.B1(n_234),
.B2(n_237),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_305),
.B1(n_319),
.B2(n_275),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_261),
.A2(n_236),
.B1(n_220),
.B2(n_219),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_286),
.B1(n_224),
.B2(n_279),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_257),
.A2(n_225),
.B(n_232),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_227),
.B1(n_266),
.B2(n_175),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_268),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_236),
.B1(n_156),
.B2(n_126),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_285),
.C(n_265),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_318),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_256),
.A2(n_219),
.B(n_232),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_243),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_310),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_286),
.B(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_258),
.A2(n_236),
.B1(n_250),
.B2(n_213),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_126),
.B1(n_240),
.B2(n_231),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_279),
.B(n_264),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_320),
.A2(n_304),
.B(n_313),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_336),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_322),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_302),
.B(n_282),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_323),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_348),
.B1(n_319),
.B2(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_326),
.A2(n_335),
.B1(n_342),
.B2(n_350),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_327),
.A2(n_347),
.B1(n_291),
.B2(n_297),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_343),
.C(n_346),
.Y(n_356)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_317),
.B(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_334),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_293),
.B1(n_317),
.B2(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_338),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_259),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_339),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_259),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_285),
.C(n_262),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_283),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_351),
.B1(n_292),
.B2(n_303),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_278),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_309),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_311),
.A2(n_277),
.B1(n_275),
.B2(n_284),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_275),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_296),
.A2(n_276),
.B1(n_287),
.B2(n_280),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_293),
.A2(n_266),
.B1(n_250),
.B2(n_227),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_346),
.B(n_311),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_364),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_345),
.A2(n_290),
.B(n_317),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_358),
.A2(n_379),
.B(n_345),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_359),
.A2(n_360),
.B1(n_365),
.B2(n_370),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_317),
.B1(n_319),
.B2(n_289),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_363),
.A2(n_347),
.B1(n_324),
.B2(n_344),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_314),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_328),
.A2(n_289),
.B1(n_308),
.B2(n_301),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_288),
.B1(n_294),
.B2(n_308),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_314),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_372),
.C(n_374),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_288),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_300),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_325),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_300),
.Y(n_374)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_299),
.B(n_312),
.Y(n_375)
);

BUFx12f_ASAP7_75t_SL g399 ( 
.A(n_375),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_348),
.A2(n_316),
.B1(n_312),
.B2(n_315),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_377),
.A2(n_342),
.B1(n_322),
.B2(n_313),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_304),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_246),
.C(n_250),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_246),
.C(n_260),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_398),
.B(n_184),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_382),
.B(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_341),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AOI32xp33_ASAP7_75t_L g388 ( 
.A1(n_370),
.A2(n_358),
.A3(n_354),
.B1(n_332),
.B2(n_367),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_388),
.A2(n_399),
.B1(n_392),
.B2(n_408),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_364),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_339),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_391),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_392),
.A2(n_359),
.B1(n_365),
.B2(n_377),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_332),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_412),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_350),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_396),
.Y(n_419)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_379),
.A2(n_335),
.B(n_326),
.Y(n_398)
);

AOI32xp33_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_334),
.A3(n_330),
.B1(n_337),
.B2(n_336),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_13),
.C(n_12),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_351),
.C(n_331),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_405),
.C(n_207),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_409),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_406),
.B1(n_352),
.B2(n_378),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_224),
.C(n_240),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_360),
.A2(n_322),
.B1(n_224),
.B2(n_178),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_226),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_226),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_410),
.B(n_411),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_362),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_205),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_422),
.B1(n_423),
.B2(n_430),
.Y(n_445)
);

FAx1_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_357),
.CI(n_374),
.CON(n_417),
.SN(n_417)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_436),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_418),
.A2(n_428),
.B1(n_431),
.B2(n_406),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_435),
.Y(n_449)
);

NOR3xp33_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_369),
.C(n_353),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_433),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_397),
.A2(n_352),
.B1(n_380),
.B2(n_366),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_397),
.A2(n_380),
.B1(n_381),
.B2(n_383),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_427),
.C(n_394),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_139),
.C(n_119),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_429),
.A2(n_408),
.B(n_385),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_90),
.B1(n_108),
.B2(n_127),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_395),
.A2(n_214),
.B1(n_119),
.B2(n_10),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_71),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_407),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_437),
.B(n_438),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_440),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_404),
.B1(n_398),
.B2(n_388),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_441),
.A2(n_443),
.B1(n_454),
.B2(n_457),
.Y(n_475)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_444),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_387),
.B1(n_389),
.B2(n_384),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_448),
.B1(n_455),
.B2(n_412),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_456),
.Y(n_470)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_450),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_420),
.B(n_386),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_403),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_431),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_386),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_401),
.B1(n_394),
.B2(n_396),
.Y(n_457)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_454),
.A2(n_443),
.B(n_453),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_464),
.B(n_450),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_452),
.A2(n_421),
.B(n_427),
.Y(n_460)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_423),
.C(n_425),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_463),
.C(n_472),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g462 ( 
.A(n_453),
.B(n_425),
.CI(n_417),
.CON(n_462),
.SN(n_462)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_0),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_417),
.C(n_422),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_441),
.A2(n_413),
.B(n_409),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_465),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_430),
.B1(n_436),
.B2(n_410),
.Y(n_466)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_32),
.C(n_24),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_32),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_449),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_445),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_491),
.C(n_471),
.Y(n_493)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_459),
.B(n_440),
.CI(n_437),
.CON(n_477),
.SN(n_477)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_481),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_486),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_451),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_487),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_468),
.B(n_470),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_475),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_0),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_44),
.C(n_2),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_479),
.A2(n_469),
.B(n_464),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_492),
.B(n_494),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_496),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_478),
.A2(n_458),
.B1(n_466),
.B2(n_472),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_488),
.A2(n_475),
.B1(n_471),
.B2(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_474),
.C(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_498),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_486),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_503),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_482),
.A2(n_3),
.B(n_4),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_502),
.A2(n_3),
.B(n_4),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_44),
.Y(n_503)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_476),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_511),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_499),
.A2(n_500),
.B(n_495),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_483),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_491),
.Y(n_515)
);

OAI321xp33_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_490),
.A3(n_477),
.B1(n_503),
.B2(n_483),
.C(n_501),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_SL g519 ( 
.A1(n_513),
.A2(n_509),
.B(n_508),
.C(n_510),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_516),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_480),
.B(n_44),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_519),
.A2(n_520),
.B(n_517),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_508),
.C(n_6),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_522),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_44),
.C(n_6),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_6),
.B(n_7),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_9),
.C(n_6),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_8),
.B(n_9),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_8),
.Y(n_527)
);


endmodule