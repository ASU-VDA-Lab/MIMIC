module fake_jpeg_24661_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_16),
.Y(n_45)
);

NAND2x1_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_13),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_18),
.B1(n_24),
.B2(n_19),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_19),
.B(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_17),
.B1(n_26),
.B2(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_63),
.B1(n_51),
.B2(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_66),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_22),
.B1(n_26),
.B2(n_17),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_0),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_46),
.Y(n_77)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_27),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_39),
.B(n_50),
.C(n_27),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_87),
.B1(n_67),
.B2(n_69),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_83),
.B1(n_89),
.B2(n_55),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_82),
.B1(n_57),
.B2(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_30),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_31),
.B(n_20),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_51),
.B1(n_37),
.B2(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_32),
.C(n_50),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_66),
.C(n_30),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_78),
.B(n_71),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_25),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_70),
.B1(n_63),
.B2(n_52),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_56),
.B1(n_65),
.B2(n_55),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_87),
.C(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_66),
.B1(n_37),
.B2(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_107),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_79),
.B1(n_84),
.B2(n_82),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_118),
.C(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_126),
.B1(n_105),
.B2(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_128),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_74),
.C(n_89),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_74),
.C(n_83),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_79),
.B1(n_73),
.B2(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_97),
.B1(n_107),
.B2(n_69),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_72),
.B(n_76),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_127),
.B(n_20),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_75),
.C(n_31),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_130),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_13),
.B(n_20),
.C(n_21),
.D(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_104),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_139),
.B1(n_143),
.B2(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

OAI22x1_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_102),
.B1(n_96),
.B2(n_95),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_69),
.B1(n_21),
.B2(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_21),
.B1(n_20),
.B2(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_123),
.B(n_125),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_119),
.C(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_160),
.C(n_163),
.Y(n_173)
);

NAND4xp25_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_161),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_111),
.B1(n_117),
.B2(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_113),
.C(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_127),
.C(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_176),
.B(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_132),
.C(n_150),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_136),
.B(n_145),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_133),
.C(n_135),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_141),
.C(n_3),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_156),
.B1(n_164),
.B2(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_151),
.B(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_188),
.B(n_192),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_191),
.C(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_158),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_157),
.A3(n_159),
.B1(n_163),
.B2(n_165),
.C1(n_152),
.C2(n_7),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_193),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_178),
.C(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_210)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_176),
.B(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_173),
.C(n_8),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_190),
.B(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_211),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_201),
.B1(n_9),
.B2(n_12),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_8),
.B(n_11),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_6),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_215),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_221),
.B(n_5),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_207),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_210),
.C(n_6),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_8),
.B(n_10),
.Y(n_225)
);

AOI221xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_10),
.B1(n_11),
.B2(n_4),
.C(n_1),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_226),
.B(n_11),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_4),
.Y(n_230)
);


endmodule