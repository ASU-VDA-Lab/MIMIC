module fake_jpeg_32021_n_69 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_4),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_18),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_26),
.C(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_5),
.B(n_6),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_9),
.B(n_10),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_60),
.B(n_55),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_21),
.C(n_24),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_65),
.B(n_57),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_59),
.B(n_48),
.Y(n_69)
);


endmodule