module real_jpeg_8204_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_347, n_6, n_348, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_347;
input n_6;
input n_348;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_1),
.A2(n_35),
.B1(n_70),
.B2(n_71),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_1),
.A2(n_35),
.B1(n_49),
.B2(n_52),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_24),
.B1(n_49),
.B2(n_52),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_2),
.A2(n_24),
.B1(n_70),
.B2(n_71),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_4),
.A2(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_49),
.B1(n_52),
.B2(n_62),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_70),
.B1(n_71),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_5),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_95),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_95),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_95),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_49),
.B1(n_52),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_70),
.B1(n_71),
.B2(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_107),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_107),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_52),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_13),
.B(n_52),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_13),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_13),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_13),
.B(n_26),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_13),
.A2(n_28),
.B(n_30),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_13),
.A2(n_23),
.B1(n_25),
.B2(n_116),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_70),
.B1(n_71),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_14),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_49),
.B1(n_52),
.B2(n_100),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_100),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_14),
.A2(n_23),
.B1(n_25),
.B2(n_100),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_15),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_15),
.A2(n_49),
.B1(n_52),
.B2(n_64),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_345),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_82),
.B(n_343),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_20),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_21),
.A2(n_37),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_22),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_22),
.A2(n_26),
.B(n_36),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_27),
.B(n_32),
.C(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_32),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_23),
.A2(n_32),
.B(n_116),
.C(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_34),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_26),
.A2(n_36),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_27),
.A2(n_37),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_27),
.A2(n_37),
.B1(n_213),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_27),
.A2(n_37),
.B1(n_222),
.B2(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_27),
.A2(n_33),
.B(n_61),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_30),
.A2(n_46),
.B(n_47),
.C(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_47),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g146 ( 
.A(n_30),
.B(n_116),
.CON(n_146),
.SN(n_146)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_37),
.A2(n_79),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_40),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_76),
.C(n_80),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_41),
.A2(n_42),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_59),
.C(n_65),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_43),
.A2(n_44),
.B1(n_65),
.B2(n_318),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_45),
.A2(n_165),
.B(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_53),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_53),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_55),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_46),
.A2(n_55),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_47),
.B(n_52),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_49),
.A2(n_56),
.B1(n_146),
.B2(n_152),
.Y(n_151)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_67),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_53),
.A2(n_55),
.B(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_54),
.A2(n_132),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_55),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_58),
.B(n_132),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_59),
.A2(n_60),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_65),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_65),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_69),
.B(n_74),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_69),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_66),
.A2(n_69),
.B1(n_106),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_66),
.A2(n_69),
.B1(n_134),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_66),
.A2(n_144),
.B(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_66),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_66),
.A2(n_69),
.B1(n_228),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_66),
.A2(n_248),
.B(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_69),
.B(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_69),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_69),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_75),
.B(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_75),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_340),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_76),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_336),
.B(n_342),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_308),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_347),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_256),
.A3(n_278),
.B1(n_301),
.B2(n_307),
.C(n_348),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_215),
.C(n_252),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_186),
.B(n_214),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_159),
.B(n_185),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_139),
.B(n_158),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_127),
.B(n_138),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_113),
.B(n_126),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_96),
.B(n_156),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_119),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_108),
.B2(n_112),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_121),
.B(n_125),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_119),
.A2(n_120),
.B1(n_171),
.B2(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_119),
.A2(n_155),
.B(n_196),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_119),
.A2(n_120),
.B(n_154),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_140),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.CI(n_135),
.CON(n_130),
.SN(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_132),
.A2(n_165),
.B1(n_167),
.B2(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_136),
.B(n_172),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_150),
.B2(n_157),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_149),
.C(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_177),
.B2(n_178),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_180),
.C(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_168),
.B1(n_169),
.B2(n_176),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_165),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_181),
.B(n_229),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_188),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_200),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_199),
.C(n_200),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_210),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_207),
.C(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_205),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_234),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_216),
.B(n_234),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.C(n_232),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_220),
.C(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_233),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_231),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_245),
.C(n_249),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_239),
.C(n_243),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_244),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_257),
.A2(n_302),
.B(n_306),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_258),
.B(n_259),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_277),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_270),
.B2(n_271),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_271),
.C(n_277),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_265),
.C(n_269),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_276),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_273),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_272),
.A2(n_287),
.B(n_290),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_279),
.B(n_280),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_299),
.B2(n_300),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_291),
.B1(n_292),
.B2(n_298),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_298),
.C(n_300),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_296),
.B(n_297),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_296),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_295),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_297),
.A2(n_310),
.B1(n_320),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_322),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_322),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_320),
.C(n_321),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_312),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_318),
.C(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_324),
.C(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_315),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_338),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_339),
.Y(n_341)
);


endmodule