module fake_jpeg_26238_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_15),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_29),
.B1(n_31),
.B2(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_31),
.B1(n_15),
.B2(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_37),
.B(n_36),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_74),
.B(n_0),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_17),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_53),
.B(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_40),
.C(n_38),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_17),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_89),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_87),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_91),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_57),
.B(n_21),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_74),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_100),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_74),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_89),
.C(n_88),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_110),
.C(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_82),
.B1(n_75),
.B2(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_106),
.B1(n_97),
.B2(n_99),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_75),
.B1(n_80),
.B2(n_67),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_73),
.C(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_100),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_73),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C1(n_2),
.C2(n_3),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_1),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_7),
.C(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_119),
.B(n_110),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_116),
.B(n_104),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_126),
.B1(n_130),
.B2(n_3),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_4),
.B(n_132),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_4),
.Y(n_134)
);


endmodule