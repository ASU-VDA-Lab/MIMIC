module fake_netlist_6_1391_n_1008 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1008);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1008;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_691;
wire n_535;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_474;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_663;
wire n_361;
wire n_508;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_22),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_21),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_121),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_46),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_105),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_163),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_112),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_11),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_100),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_92),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_73),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_95),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_125),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_94),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_193),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_149),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_65),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_117),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_170),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_153),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_101),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_190),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_37),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_96),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_113),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_111),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_22),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_93),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_11),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_75),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_83),
.Y(n_266)
);

BUFx8_ASAP7_75t_SL g267 ( 
.A(n_34),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_159),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_131),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_18),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_152),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_62),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_184),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_155),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_207),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_0),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_0),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_197),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_199),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_1),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_1),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

CKINVDCx6p67_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_195),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_201),
.B(n_2),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_33),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_206),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_191),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_2),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_189),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_3),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_4),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_198),
.B(n_4),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_205),
.B(n_5),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_219),
.B(n_35),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_217),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_203),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_5),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_36),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_216),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_226),
.B(n_187),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_230),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_203),
.B(n_6),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_233),
.B(n_6),
.Y(n_323)
);

NAND2x1p5_ASAP7_75t_L g324 ( 
.A(n_235),
.B(n_7),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_204),
.B(n_7),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_204),
.B(n_277),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g328 ( 
.A(n_208),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

AO22x2_ASAP7_75t_L g332 ( 
.A1(n_286),
.A2(n_243),
.B1(n_245),
.B2(n_249),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_250),
.B1(n_252),
.B2(n_259),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_208),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_282),
.A2(n_275),
.B1(n_206),
.B2(n_210),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_283),
.A2(n_275),
.B1(n_210),
.B2(n_234),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g341 ( 
.A1(n_286),
.A2(n_256),
.B1(n_9),
.B2(n_10),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_296),
.A2(n_234),
.B1(n_273),
.B2(n_274),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_291),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_286),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g345 ( 
.A1(n_289),
.A2(n_273),
.B1(n_274),
.B2(n_277),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_209),
.Y(n_347)
);

AO22x2_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_313),
.Y(n_350)
);

OR2x6_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_209),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_238),
.B1(n_269),
.B2(n_266),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_281),
.B(n_238),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_214),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_324),
.A2(n_271),
.B1(n_263),
.B2(n_260),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_300),
.A2(n_258),
.B1(n_255),
.B2(n_253),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_232),
.B1(n_247),
.B2(n_246),
.Y(n_360)
);

AO22x2_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_231),
.B1(n_244),
.B2(n_242),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_284),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_215),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_312),
.A2(n_248),
.B1(n_239),
.B2(n_237),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_294),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_236),
.B1(n_224),
.B2(n_222),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_320),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_218),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g371 ( 
.A1(n_291),
.A2(n_221),
.B1(n_220),
.B2(n_17),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_322),
.A2(n_325),
.B1(n_304),
.B2(n_293),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_284),
.B1(n_285),
.B2(n_328),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_288),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_288),
.A2(n_293),
.B1(n_292),
.B2(n_295),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_326),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_38),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_297),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_39),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_292),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_285),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_328),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_27),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_342),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_347),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_330),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_316),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_312),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_321),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_320),
.Y(n_406)
);

NOR2x1p5_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_311),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_356),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_342),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_321),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_339),
.B(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_316),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_316),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_379),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_372),
.B(n_302),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_316),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_319),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_302),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

OR2x6_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_292),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_344),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_340),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

NAND2x1_ASAP7_75t_L g440 ( 
.A(n_351),
.B(n_308),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_351),
.B(n_319),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_351),
.B(n_319),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_360),
.B(n_319),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_309),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_362),
.B(n_359),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_366),
.B(n_292),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_343),
.B(n_309),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_339),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_335),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_295),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_295),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

BUFx4f_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_418),
.B(n_295),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_298),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_428),
.B(n_298),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_448),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_298),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_414),
.B(n_298),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_407),
.B(n_303),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_303),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_303),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_410),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_303),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_317),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_426),
.B(n_317),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_352),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_411),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_445),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_415),
.B(n_311),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_424),
.B(n_308),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_443),
.B(n_359),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_437),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_445),
.B(n_374),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_437),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_452),
.B(n_317),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_453),
.B(n_315),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_421),
.B(n_308),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_445),
.B(n_308),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_397),
.B(n_287),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_310),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_420),
.B(n_382),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_287),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_301),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_40),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_447),
.A2(n_386),
.B(n_385),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_301),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_389),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_434),
.B(n_290),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_405),
.B(n_290),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_450),
.B(n_310),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_310),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_391),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_392),
.Y(n_528)
);

AND2x2_ASAP7_75t_SL g529 ( 
.A(n_450),
.B(n_310),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_310),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_405),
.B(n_318),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_454),
.B(n_318),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_401),
.B(n_371),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_425),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_456),
.B(n_318),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_436),
.B(n_290),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_406),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_436),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_318),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_318),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_434),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_468),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_470),
.B(n_435),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_464),
.B(n_460),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

BUFx2_ASAP7_75t_SL g549 ( 
.A(n_493),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_496),
.B(n_514),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_496),
.B(n_446),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_464),
.B(n_433),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_514),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_459),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_487),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_496),
.B(n_395),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_469),
.B(n_439),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_459),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_544),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_441),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_487),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_463),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_540),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g570 ( 
.A(n_470),
.B(n_442),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_519),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_444),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_470),
.B(n_462),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_335),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_519),
.Y(n_575)
);

BUFx4_ASAP7_75t_SL g576 ( 
.A(n_501),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_455),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_462),
.B(n_451),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_451),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_471),
.B(n_28),
.Y(n_580)
);

AO21x2_ASAP7_75t_L g581 ( 
.A1(n_512),
.A2(n_461),
.B(n_455),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_471),
.B(n_30),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_463),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_516),
.B(n_461),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_297),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

BUFx4f_ASAP7_75t_SL g588 ( 
.A(n_499),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_487),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_520),
.B(n_515),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_510),
.B(n_393),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_520),
.B(n_515),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_510),
.B(n_393),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_327),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_413),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_534),
.B(n_413),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_489),
.B(n_490),
.Y(n_601)
);

AO21x2_ASAP7_75t_L g602 ( 
.A1(n_512),
.A2(n_327),
.B(n_107),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_515),
.B(n_41),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_497),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_492),
.B(n_42),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_527),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_504),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_472),
.B(n_327),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_555),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_548),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_597),
.Y(n_612)
);

BUFx2_ASAP7_75t_R g613 ( 
.A(n_549),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_551),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_576),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_548),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_594),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_596),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_599),
.Y(n_620)
);

CKINVDCx14_ASAP7_75t_R g621 ( 
.A(n_600),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_562),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_601),
.B(n_478),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_554),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_600),
.A2(n_518),
.B1(n_529),
.B2(n_525),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_557),
.B(n_502),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_546),
.A2(n_518),
.B1(n_525),
.B2(n_529),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_554),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_546),
.B(n_500),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_576),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_588),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_557),
.B(n_513),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_591),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_548),
.Y(n_639)
);

BUFx2_ASAP7_75t_SL g640 ( 
.A(n_590),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_580),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_589),
.Y(n_642)
);

BUFx4f_ASAP7_75t_SL g643 ( 
.A(n_579),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_563),
.B(n_478),
.Y(n_644)
);

BUFx4f_ASAP7_75t_SL g645 ( 
.A(n_604),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_582),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_588),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_595),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_606),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_595),
.Y(n_650)
);

BUFx12f_ASAP7_75t_L g651 ( 
.A(n_552),
.Y(n_651)
);

INVx3_ASAP7_75t_SL g652 ( 
.A(n_552),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

CKINVDCx14_ASAP7_75t_R g654 ( 
.A(n_603),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_563),
.B(n_490),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_575),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_589),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_547),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_589),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_545),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_589),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_592),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_570),
.B(n_523),
.Y(n_663)
);

INVx6_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_523),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_550),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_592),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_565),
.B(n_547),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_637),
.B(n_565),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_627),
.A2(n_529),
.B1(n_525),
.B2(n_578),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_635),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_630),
.A2(n_578),
.B1(n_573),
.B2(n_492),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_628),
.A2(n_573),
.B1(n_532),
.B2(n_605),
.Y(n_674)
);

CKINVDCx11_ASAP7_75t_R g675 ( 
.A(n_612),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_653),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_620),
.B(n_618),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_649),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_654),
.A2(n_569),
.B1(n_500),
.B2(n_466),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_616),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_620),
.B(n_497),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_656),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_658),
.A2(n_532),
.B1(n_531),
.B2(n_507),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_663),
.A2(n_531),
.B1(n_507),
.B2(n_533),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_621),
.A2(n_577),
.B1(n_585),
.B2(n_603),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_649),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_621),
.A2(n_513),
.B(n_553),
.Y(n_687)
);

BUFx8_ASAP7_75t_L g688 ( 
.A(n_651),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_669),
.A2(n_566),
.B1(n_561),
.B2(n_553),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_611),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_655),
.B(n_513),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_666),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_666),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_663),
.A2(n_533),
.B1(n_480),
.B2(n_506),
.Y(n_694)
);

INVx6_ASAP7_75t_L g695 ( 
.A(n_651),
.Y(n_695)
);

CKINVDCx11_ASAP7_75t_R g696 ( 
.A(n_612),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_610),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_624),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_635),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_665),
.A2(n_480),
.B1(n_506),
.B2(n_484),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_625),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_665),
.A2(n_484),
.B1(n_537),
.B2(n_566),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_616),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_619),
.A2(n_561),
.B1(n_466),
.B2(n_572),
.Y(n_704)
);

CKINVDCx11_ASAP7_75t_R g705 ( 
.A(n_634),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_660),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_648),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_633),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_623),
.A2(n_530),
.B1(n_479),
.B2(n_577),
.Y(n_710)
);

CKINVDCx11_ASAP7_75t_R g711 ( 
.A(n_636),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_638),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_638),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_644),
.A2(n_530),
.B1(n_479),
.B2(n_585),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_632),
.A2(n_530),
.B1(n_503),
.B2(n_482),
.Y(n_715)
);

AOI21xp33_ASAP7_75t_L g716 ( 
.A1(n_641),
.A2(n_509),
.B(n_488),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_617),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_648),
.Y(n_718)
);

BUFx12f_ASAP7_75t_L g719 ( 
.A(n_617),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_646),
.B(n_538),
.Y(n_720)
);

BUFx4_ASAP7_75t_SL g721 ( 
.A(n_636),
.Y(n_721)
);

INVx6_ASAP7_75t_SL g722 ( 
.A(n_613),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_667),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_650),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_667),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_677),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_671),
.A2(n_622),
.B1(n_643),
.B2(n_654),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_709),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_720),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_691),
.B(n_647),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_SL g731 ( 
.A1(n_687),
.A2(n_517),
.B(n_560),
.Y(n_731)
);

AOI222xp33_ASAP7_75t_L g732 ( 
.A1(n_671),
.A2(n_466),
.B1(n_614),
.B2(n_615),
.C1(n_626),
.C2(n_631),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_678),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_670),
.A2(n_530),
.B1(n_608),
.B2(n_598),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_676),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_670),
.A2(n_608),
.B1(n_598),
.B2(n_482),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_686),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_695),
.A2(n_640),
.B1(n_650),
.B2(n_615),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_685),
.A2(n_572),
.B1(n_652),
.B2(n_626),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_681),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_679),
.A2(n_539),
.B1(n_614),
.B2(n_631),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_673),
.A2(n_503),
.B1(n_517),
.B2(n_652),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_723),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_673),
.B(n_538),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_698),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_698),
.Y(n_747)
);

AOI211xp5_ASAP7_75t_L g748 ( 
.A1(n_704),
.A2(n_535),
.B(n_517),
.C(n_536),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_697),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_SL g750 ( 
.A1(n_674),
.A2(n_517),
.B(n_560),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_674),
.A2(n_524),
.B(n_521),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_689),
.A2(n_498),
.B1(n_467),
.B2(n_524),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_694),
.A2(n_491),
.B1(n_504),
.B2(n_645),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_701),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_718),
.B(n_542),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_689),
.B(n_542),
.Y(n_756)
);

CKINVDCx6p67_ASAP7_75t_R g757 ( 
.A(n_675),
.Y(n_757)
);

OAI222xp33_ASAP7_75t_L g758 ( 
.A1(n_694),
.A2(n_488),
.B1(n_498),
.B2(n_509),
.C1(n_521),
.C2(n_574),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_706),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_700),
.A2(n_467),
.B1(n_491),
.B2(n_543),
.Y(n_760)
);

OAI21xp33_ASAP7_75t_L g761 ( 
.A1(n_700),
.A2(n_543),
.B(n_508),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_SL g763 ( 
.A1(n_704),
.A2(n_509),
.B(n_488),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_715),
.A2(n_710),
.B1(n_683),
.B2(n_714),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_702),
.A2(n_684),
.B1(n_683),
.B2(n_710),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_699),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_672),
.A2(n_491),
.B1(n_488),
.B2(n_509),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_712),
.B(n_536),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_725),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_702),
.A2(n_684),
.B1(n_714),
.B2(n_716),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

BUFx2_ASAP7_75t_SL g773 ( 
.A(n_672),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_722),
.A2(n_467),
.B1(n_536),
.B2(n_475),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_699),
.B(n_708),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_708),
.B(n_467),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_722),
.A2(n_475),
.B1(n_494),
.B2(n_483),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_695),
.A2(n_574),
.B1(n_508),
.B2(n_522),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_715),
.A2(n_526),
.B(n_477),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_724),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_695),
.A2(n_504),
.B1(n_556),
.B2(n_567),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_SL g784 ( 
.A1(n_722),
.A2(n_721),
.B(n_696),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_SL g785 ( 
.A1(n_688),
.A2(n_504),
.B1(n_611),
.B2(n_602),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

BUFx8_ASAP7_75t_SL g787 ( 
.A(n_703),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_727),
.A2(n_688),
.B1(n_711),
.B2(n_705),
.Y(n_788)
);

OAI222xp33_ASAP7_75t_L g789 ( 
.A1(n_727),
.A2(n_574),
.B1(n_690),
.B2(n_568),
.C1(n_583),
.C2(n_587),
.Y(n_789)
);

OAI221xp5_ASAP7_75t_SL g790 ( 
.A1(n_763),
.A2(n_475),
.B1(n_477),
.B2(n_483),
.C(n_485),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_765),
.A2(n_494),
.B1(n_477),
.B2(n_483),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_764),
.A2(n_680),
.B1(n_713),
.B2(n_504),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_747),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_765),
.A2(n_485),
.B1(n_494),
.B2(n_713),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_747),
.B(n_746),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_741),
.A2(n_485),
.B1(n_680),
.B2(n_527),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_762),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_726),
.B(n_717),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_771),
.A2(n_528),
.B1(n_527),
.B2(n_504),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_730),
.B(n_717),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_771),
.A2(n_528),
.B1(n_522),
.B2(n_581),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_SL g802 ( 
.A1(n_748),
.A2(n_707),
.B1(n_690),
.B2(n_642),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_743),
.B(n_752),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_761),
.A2(n_528),
.B1(n_522),
.B2(n_581),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_732),
.A2(n_522),
.B1(n_602),
.B2(n_526),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_SL g806 ( 
.A(n_778),
.B(n_586),
.C(n_584),
.Y(n_806)
);

OAI222xp33_ASAP7_75t_L g807 ( 
.A1(n_743),
.A2(n_593),
.B1(n_609),
.B2(n_639),
.C1(n_661),
.C2(n_586),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_751),
.A2(n_729),
.B1(n_745),
.B2(n_740),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_766),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_733),
.B(n_639),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_752),
.A2(n_522),
.B1(n_558),
.B2(n_511),
.Y(n_811)
);

OAI222xp33_ASAP7_75t_L g812 ( 
.A1(n_778),
.A2(n_609),
.B1(n_661),
.B2(n_639),
.C1(n_558),
.C2(n_511),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_774),
.A2(n_707),
.B1(n_607),
.B2(n_592),
.Y(n_813)
);

AOI222xp33_ASAP7_75t_L g814 ( 
.A1(n_750),
.A2(n_522),
.B1(n_327),
.B2(n_32),
.C1(n_31),
.C2(n_30),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_774),
.B(n_327),
.C(n_657),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_753),
.A2(n_522),
.B1(n_511),
.B2(n_607),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_767),
.A2(n_522),
.B1(n_661),
.B2(n_664),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_731),
.A2(n_784),
.B(n_758),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_733),
.B(n_617),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_738),
.A2(n_707),
.B1(n_611),
.B2(n_567),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_773),
.A2(n_611),
.B1(n_668),
.B2(n_662),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_769),
.B(n_617),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_737),
.B(n_617),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_735),
.B(n_629),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_742),
.A2(n_556),
.B1(n_567),
.B2(n_664),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_776),
.B(n_756),
.C(n_775),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_757),
.A2(n_664),
.B1(n_474),
.B2(n_476),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_781),
.A2(n_668),
.B1(n_662),
.B2(n_659),
.Y(n_828)
);

AOI222xp33_ASAP7_75t_L g829 ( 
.A1(n_736),
.A2(n_755),
.B1(n_749),
.B2(n_739),
.C1(n_754),
.C2(n_759),
.Y(n_829)
);

OA222x2_ASAP7_75t_L g830 ( 
.A1(n_770),
.A2(n_31),
.B1(n_32),
.B2(n_473),
.C1(n_465),
.C2(n_474),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_737),
.B(n_629),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_744),
.B(n_629),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_728),
.A2(n_664),
.B1(n_474),
.B2(n_476),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_736),
.A2(n_474),
.B1(n_476),
.B2(n_486),
.Y(n_834)
);

OAI222xp33_ASAP7_75t_L g835 ( 
.A1(n_779),
.A2(n_473),
.B1(n_465),
.B2(n_486),
.C1(n_476),
.C2(n_567),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_760),
.A2(n_486),
.B1(n_473),
.B2(n_659),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_772),
.B(n_629),
.Y(n_837)
);

AOI221xp5_ASAP7_75t_L g838 ( 
.A1(n_734),
.A2(n_473),
.B1(n_486),
.B2(n_297),
.C(n_657),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_768),
.B(n_629),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_782),
.B(n_657),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_734),
.B(n_772),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_760),
.A2(n_668),
.B1(n_662),
.B2(n_659),
.Y(n_842)
);

OAI221xp5_ASAP7_75t_L g843 ( 
.A1(n_818),
.A2(n_785),
.B1(n_786),
.B2(n_780),
.C(n_783),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_809),
.B(n_777),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_826),
.B(n_787),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_SL g846 ( 
.A1(n_814),
.A2(n_787),
.B(n_668),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_788),
.A2(n_792),
.B1(n_808),
.B2(n_796),
.C(n_802),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_809),
.B(n_657),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_824),
.B(n_657),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_800),
.B(n_659),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_803),
.A2(n_668),
.B1(n_662),
.B2(n_659),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_798),
.B(n_662),
.Y(n_852)
);

OA21x2_ASAP7_75t_L g853 ( 
.A1(n_792),
.A2(n_556),
.B(n_297),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_829),
.B(n_43),
.Y(n_854)
);

OAI221xp5_ASAP7_75t_SL g855 ( 
.A1(n_805),
.A2(n_830),
.B1(n_794),
.B2(n_842),
.C(n_801),
.Y(n_855)
);

OAI221xp5_ASAP7_75t_SL g856 ( 
.A1(n_830),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.C(n_49),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_795),
.B(n_50),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_SL g858 ( 
.A1(n_789),
.A2(n_51),
.B(n_53),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_795),
.B(n_54),
.Y(n_859)
);

NAND4xp25_ASAP7_75t_L g860 ( 
.A(n_841),
.B(n_56),
.C(n_57),
.D(n_58),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_797),
.B(n_59),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_SL g862 ( 
.A1(n_811),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.C(n_64),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_802),
.B(n_66),
.Y(n_863)
);

OAI221xp5_ASAP7_75t_SL g864 ( 
.A1(n_804),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.C(n_71),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_797),
.B(n_72),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_L g866 ( 
.A(n_790),
.B(n_815),
.C(n_820),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_803),
.A2(n_815),
.B1(n_827),
.B2(n_817),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_791),
.B(n_833),
.C(n_799),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_824),
.B(n_74),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_832),
.B(n_76),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_840),
.B(n_556),
.C(n_79),
.Y(n_871)
);

NAND4xp25_ASAP7_75t_SL g872 ( 
.A(n_838),
.B(n_78),
.C(n_80),
.D(n_81),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_825),
.A2(n_185),
.B1(n_84),
.B2(n_85),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_822),
.B(n_82),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_806),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_816),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_793),
.B(n_102),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_822),
.B(n_103),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_836),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_L g880 ( 
.A(n_828),
.B(n_109),
.C(n_114),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_821),
.B(n_116),
.C(n_119),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_807),
.A2(n_120),
.B(n_122),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_813),
.A2(n_123),
.B(n_124),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_793),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_884),
.B(n_837),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_844),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_858),
.A2(n_872),
.B(n_875),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_852),
.B(n_831),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_853),
.B(n_839),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_853),
.B(n_837),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_850),
.B(n_823),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_860),
.A2(n_834),
.B1(n_831),
.B2(n_810),
.Y(n_892)
);

NOR2x1_ASAP7_75t_SL g893 ( 
.A(n_851),
.B(n_819),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_849),
.B(n_126),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_845),
.B(n_848),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_849),
.B(n_127),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_856),
.B(n_835),
.C(n_812),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_882),
.B(n_874),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_845),
.B(n_128),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_866),
.A2(n_129),
.B(n_130),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_882),
.B(n_132),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_878),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_857),
.B(n_859),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_854),
.B(n_135),
.C(n_136),
.Y(n_904)
);

NAND4xp75_ASAP7_75t_L g905 ( 
.A(n_863),
.B(n_138),
.C(n_139),
.D(n_140),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_869),
.B(n_142),
.Y(n_906)
);

NAND4xp75_ASAP7_75t_L g907 ( 
.A(n_863),
.B(n_144),
.C(n_145),
.D(n_148),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_866),
.B(n_150),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_861),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_865),
.B(n_156),
.Y(n_910)
);

OAI211xp5_ASAP7_75t_SL g911 ( 
.A1(n_846),
.A2(n_157),
.B(n_158),
.C(n_160),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_885),
.Y(n_912)
);

XNOR2xp5_ASAP7_75t_L g913 ( 
.A(n_902),
.B(n_847),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_885),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_895),
.B(n_843),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_885),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_885),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_909),
.B(n_867),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_886),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_893),
.Y(n_921)
);

XOR2xp5_ASAP7_75t_L g922 ( 
.A(n_902),
.B(n_870),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_886),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_909),
.B(n_877),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_894),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_888),
.B(n_875),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_891),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_904),
.B(n_864),
.C(n_862),
.Y(n_928)
);

NOR2x1_ASAP7_75t_R g929 ( 
.A(n_899),
.B(n_855),
.Y(n_929)
);

NOR4xp75_ASAP7_75t_L g930 ( 
.A(n_905),
.B(n_883),
.C(n_881),
.D(n_880),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_920),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_927),
.B(n_891),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_925),
.Y(n_933)
);

XOR2xp5_ASAP7_75t_L g934 ( 
.A(n_913),
.B(n_887),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_925),
.Y(n_935)
);

OA22x2_ASAP7_75t_L g936 ( 
.A1(n_921),
.A2(n_908),
.B1(n_898),
.B2(n_894),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_914),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_915),
.B(n_903),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_912),
.Y(n_940)
);

XOR2x2_ASAP7_75t_L g941 ( 
.A(n_922),
.B(n_907),
.Y(n_941)
);

XOR2xp5_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_903),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_934),
.A2(n_917),
.B1(n_915),
.B2(n_928),
.Y(n_943)
);

OA22x2_ASAP7_75t_L g944 ( 
.A1(n_934),
.A2(n_921),
.B1(n_919),
.B2(n_923),
.Y(n_944)
);

XNOR2x1_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_930),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_932),
.Y(n_946)
);

XOR2xp5_ASAP7_75t_L g947 ( 
.A(n_942),
.B(n_936),
.Y(n_947)
);

OA22x2_ASAP7_75t_L g948 ( 
.A1(n_942),
.A2(n_918),
.B1(n_916),
.B2(n_908),
.Y(n_948)
);

AO22x1_ASAP7_75t_L g949 ( 
.A1(n_939),
.A2(n_917),
.B1(n_928),
.B2(n_901),
.Y(n_949)
);

XOR2x2_ASAP7_75t_L g950 ( 
.A(n_933),
.B(n_905),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_935),
.B(n_929),
.Y(n_951)
);

AOI22x1_ASAP7_75t_L g952 ( 
.A1(n_935),
.A2(n_898),
.B1(n_894),
.B2(n_906),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_931),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_944),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_953),
.Y(n_955)
);

OAI322xp33_ASAP7_75t_L g956 ( 
.A1(n_945),
.A2(n_926),
.A3(n_924),
.B1(n_938),
.B2(n_904),
.C1(n_889),
.C2(n_940),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_946),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_950),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_948),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_954),
.A2(n_943),
.B1(n_947),
.B2(n_951),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_954),
.A2(n_947),
.B1(n_949),
.B2(n_900),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_954),
.A2(n_900),
.B1(n_911),
.B2(n_917),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_955),
.Y(n_963)
);

OAI31xp33_ASAP7_75t_L g964 ( 
.A1(n_961),
.A2(n_959),
.A3(n_958),
.B(n_957),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_963),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_960),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_962),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_966),
.A2(n_917),
.B1(n_900),
.B2(n_937),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_964),
.B(n_952),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_965),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_966),
.B(n_956),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_889),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

OA22x2_ASAP7_75t_L g974 ( 
.A1(n_966),
.A2(n_894),
.B1(n_896),
.B2(n_873),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_970),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_973),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_972),
.Y(n_978)
);

NOR2x2_ASAP7_75t_L g979 ( 
.A(n_971),
.B(n_907),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_969),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_980),
.B(n_968),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_978),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_975),
.Y(n_983)
);

NAND2x1_ASAP7_75t_L g984 ( 
.A(n_976),
.B(n_896),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_979),
.A2(n_906),
.B1(n_897),
.B2(n_910),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_982),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_985),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_981),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_986),
.B(n_893),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_990),
.A2(n_984),
.B1(n_979),
.B2(n_871),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_988),
.A2(n_890),
.B1(n_892),
.B2(n_876),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_SL g994 ( 
.A1(n_987),
.A2(n_879),
.B1(n_876),
.B2(n_868),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_989),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_995),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_992),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_994),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_997),
.A2(n_991),
.B1(n_993),
.B2(n_890),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_998),
.A2(n_991),
.B1(n_879),
.B2(n_164),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_999),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_1000),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_1001),
.A2(n_996),
.B1(n_162),
.B2(n_165),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_1002),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1003),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1004),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_1006),
.A2(n_168),
.B1(n_171),
.B2(n_173),
.C(n_175),
.Y(n_1007)
);

AOI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_1007),
.A2(n_1005),
.B(n_179),
.C(n_183),
.Y(n_1008)
);


endmodule