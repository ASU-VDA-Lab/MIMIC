module fake_jpeg_18373_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_45),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_9),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_60),
.Y(n_110)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_77),
.Y(n_118)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_64),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_35),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_73),
.B(n_74),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_19),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_22),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_30),
.B1(n_37),
.B2(n_35),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_33),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_17),
.B(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_23),
.C(n_28),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_62),
.C(n_80),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_28),
.B(n_23),
.C(n_37),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_62),
.B(n_64),
.C(n_79),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_28),
.B1(n_36),
.B2(n_32),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_107),
.B1(n_112),
.B2(n_92),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_36),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_131),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_109),
.Y(n_142)
);

NOR2x1_ASAP7_75t_R g147 ( 
.A(n_105),
.B(n_85),
.Y(n_147)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_31),
.B1(n_30),
.B2(n_17),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_37),
.A3(n_35),
.B1(n_10),
.B2(n_12),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_119),
.Y(n_163)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_90),
.B1(n_8),
.B2(n_10),
.Y(n_164)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_8),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_145),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_152),
.B1(n_159),
.B2(n_160),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_65),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_146),
.A2(n_147),
.B(n_160),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_103),
.C(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_72),
.B1(n_89),
.B2(n_58),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_164),
.B1(n_113),
.B2(n_95),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_75),
.B1(n_67),
.B2(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_96),
.A2(n_78),
.B1(n_75),
.B2(n_67),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_111),
.B1(n_95),
.B2(n_100),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_111),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_123),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_147),
.B(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_169),
.B1(n_191),
.B2(n_137),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_171),
.Y(n_209)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_181),
.B(n_13),
.Y(n_210)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

NAND2x1_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_108),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_180),
.B(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_128),
.B(n_118),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_109),
.B(n_124),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_141),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_125),
.B(n_107),
.C(n_97),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_144),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_99),
.B(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_197),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_116),
.C(n_132),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_151),
.C(n_165),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_199),
.B(n_226),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_212),
.C(n_192),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_142),
.A3(n_136),
.B1(n_133),
.B2(n_137),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_183),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_133),
.B1(n_144),
.B2(n_134),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_207),
.B1(n_227),
.B2(n_167),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_227),
.B1(n_202),
.B2(n_213),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_210),
.B(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_149),
.C(n_135),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_157),
.B(n_145),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_214),
.B(n_221),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_175),
.B(n_7),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_223),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_1),
.B(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_6),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_188),
.B1(n_195),
.B2(n_177),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_6),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_235),
.B1(n_241),
.B2(n_244),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_179),
.C(n_170),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_233),
.A2(n_240),
.B(n_242),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_201),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_234),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_187),
.B1(n_186),
.B2(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_201),
.C(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_189),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_172),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_210),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_172),
.B1(n_171),
.B2(n_185),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_217),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_184),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_252),
.B(n_250),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_223),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_176),
.B1(n_196),
.B2(n_198),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_255),
.B1(n_245),
.B2(n_241),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_229),
.A2(n_202),
.B1(n_218),
.B2(n_214),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_215),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_211),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_211),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_205),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_205),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_204),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_238),
.C(n_236),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_273),
.B1(n_242),
.B2(n_240),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_239),
.B1(n_230),
.B2(n_237),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_281),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_257),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_232),
.C(n_230),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_277),
.C(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_232),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_204),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_293),
.Y(n_302)
);

OAI221xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_258),
.B1(n_260),
.B2(n_268),
.C(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_267),
.C(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_255),
.B1(n_264),
.B2(n_265),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_294),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_274),
.B(n_275),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_238),
.C(n_271),
.Y(n_296)
);

NAND4xp25_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_190),
.C(n_196),
.D(n_224),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_305),
.Y(n_312)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_277),
.B(n_274),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_290),
.B1(n_288),
.B2(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_287),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_190),
.B(n_4),
.C(n_5),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_3),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_297),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_314),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_312),
.B(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_3),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_302),
.C(n_299),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_312),
.B1(n_296),
.B2(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_319),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_323),
.B(n_322),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_316),
.C(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_315),
.C(n_11),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_11),
.B(n_14),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_16),
.Y(n_329)
);


endmodule