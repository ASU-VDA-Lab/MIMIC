module fake_jpeg_8870_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_11),
.B1(n_16),
.B2(n_14),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_22),
.B1(n_9),
.B2(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_2),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_35),
.B(n_26),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_23),
.B(n_21),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_21),
.C(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_45),
.B1(n_40),
.B2(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_37),
.CI(n_45),
.CON(n_53),
.SN(n_53)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_50),
.C(n_7),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_51),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_53),
.B1(n_30),
.B2(n_19),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule