module real_jpeg_14497_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_84),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_84),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_57),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_26),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_51),
.C(n_90),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_72),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_47),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_11),
.B(n_124),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_12),
.A2(n_27),
.B1(n_69),
.B2(n_70),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_97),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_97),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_59),
.B2(n_60),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_46),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_23),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_25),
.A2(n_30),
.B1(n_113),
.B2(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_28),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_26),
.A2(n_44),
.B(n_68),
.C(n_73),
.Y(n_67)
);

HAxp5_ASAP7_75t_SL g113 ( 
.A(n_26),
.B(n_72),
.CON(n_113),
.SN(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_45),
.C(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x4_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_35),
.B(n_113),
.C(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_35),
.A2(n_37),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_35),
.B(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_68),
.B1(n_76),
.B2(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_45),
.B1(n_69),
.B2(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_54),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_56),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_47),
.B(n_72),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_47),
.A2(n_147),
.B1(n_155),
.B2(n_156),
.Y(n_159)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_48),
.A2(n_58),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_48),
.B(n_110),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_51),
.B1(n_88),
.B2(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_50),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.CON(n_68),
.SN(n_68)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_72),
.B(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_96),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_94),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_86),
.A2(n_127),
.B1(n_143),
.B2(n_144),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g90 ( 
.A(n_88),
.Y(n_90)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_103),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.C(n_106),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_132),
.B(n_179),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_129),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_121),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_125),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_173),
.B(n_178),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_162),
.B(n_172),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_150),
.B(n_161),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_145),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_156),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_157),
.B(n_160),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);


endmodule