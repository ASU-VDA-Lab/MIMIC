module fake_jpeg_13985_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_22),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_9),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_53),
.CI(n_80),
.CON(n_94),
.SN(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_79),
.B(n_56),
.C(n_57),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_73),
.B1(n_60),
.B2(n_65),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_107),
.B1(n_66),
.B2(n_58),
.Y(n_112)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_81),
.B1(n_68),
.B2(n_69),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_72),
.C(n_63),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_65),
.B1(n_69),
.B2(n_66),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_78),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_114),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_99),
.B1(n_106),
.B2(n_64),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_113),
.B(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_123),
.B1(n_124),
.B2(n_11),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_61),
.B(n_67),
.C(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_125),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_96),
.B1(n_102),
.B2(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_21),
.C(n_44),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_13),
.B1(n_17),
.B2(n_19),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_143),
.B1(n_48),
.B2(n_25),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_32),
.B(n_34),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_23),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_10),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_142),
.B(n_145),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_155),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_154),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_156),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_26),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_158),
.C(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_28),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_42),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_141),
.C(n_136),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.C(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_163),
.B1(n_162),
.B2(n_150),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_164),
.B(n_168),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_164),
.B(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_157),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_147),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_137),
.Y(n_176)
);


endmodule