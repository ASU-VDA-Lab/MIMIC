module fake_jpeg_2940_n_65 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_65);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_23),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_17),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_31),
.B1(n_0),
.B2(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_18),
.B1(n_19),
.B2(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_19),
.C(n_27),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_32),
.C(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_50),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_12),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.C(n_7),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_4),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_13),
.C(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_45),
.CI(n_6),
.CON(n_54),
.SN(n_54)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_8),
.C(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_62),
.B(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

AOI221xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_61),
.B1(n_60),
.B2(n_16),
.C(n_14),
.Y(n_65)
);


endmodule