module fake_jpeg_29443_n_382 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_57),
.Y(n_89)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_16),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_63),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_75),
.Y(n_83)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_77),
.B1(n_79),
.B2(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_78),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_39),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_30),
.B1(n_19),
.B2(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_91),
.B1(n_107),
.B2(n_109),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_82),
.A2(n_90),
.B1(n_104),
.B2(n_120),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_86),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_25),
.B(n_37),
.C(n_26),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_87),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_43),
.B1(n_34),
.B2(n_24),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_8),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_26),
.B1(n_41),
.B2(n_36),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_56),
.B1(n_62),
.B2(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_40),
.B1(n_31),
.B2(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_97),
.B1(n_108),
.B2(n_114),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_31),
.B1(n_40),
.B2(n_18),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_43),
.B1(n_24),
.B2(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_37),
.B1(n_31),
.B2(n_38),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_18),
.B1(n_38),
.B2(n_36),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_18),
.B1(n_33),
.B2(n_41),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_39),
.B1(n_9),
.B2(n_10),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_113),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_47),
.A2(n_39),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_39),
.B1(n_9),
.B2(n_11),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_0),
.C(n_2),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_73),
.C(n_3),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_80),
.B(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_126),
.B(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_76),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_12),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_106),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_59),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_73),
.B1(n_12),
.B2(n_50),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_59),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_64),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_88),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_145),
.B(n_156),
.Y(n_202)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_111),
.C(n_84),
.Y(n_175)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx6p67_ASAP7_75t_R g152 ( 
.A(n_93),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_91),
.A2(n_55),
.B1(n_49),
.B2(n_50),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_166),
.B1(n_124),
.B2(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_50),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_12),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_159),
.B1(n_90),
.B2(n_82),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_83),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_163),
.B1(n_125),
.B2(n_5),
.Y(n_197)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_103),
.B1(n_99),
.B2(n_117),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_102),
.B(n_92),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_173),
.B1(n_199),
.B2(n_128),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_115),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_175),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_87),
.B1(n_122),
.B2(n_116),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_99),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_177),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_125),
.B1(n_117),
.B2(n_92),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_138),
.B1(n_152),
.B2(n_149),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_117),
.B(n_124),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_198),
.B(n_166),
.Y(n_211)
);

OR2x2_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_121),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_152),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_130),
.B(n_116),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_122),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_163),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_137),
.A2(n_124),
.B(n_121),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_129),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_142),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_212),
.B1(n_215),
.B2(n_220),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_211),
.B(n_174),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_208),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_152),
.B(n_140),
.C(n_139),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_210),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_128),
.B1(n_139),
.B2(n_157),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_131),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_150),
.B1(n_161),
.B2(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_182),
.A2(n_147),
.B1(n_134),
.B2(n_158),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_236),
.B1(n_198),
.B2(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_146),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_226),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_148),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_229),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_151),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_230),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_141),
.B(n_158),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_207),
.B(n_209),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_235),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_194),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_175),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_177),
.B1(n_167),
.B2(n_186),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_237),
.B(n_220),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_167),
.C(n_189),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_245),
.C(n_261),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_180),
.B1(n_168),
.B2(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_244),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_180),
.B1(n_193),
.B2(n_187),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_170),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_185),
.B(n_187),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_218),
.A2(n_185),
.B(n_195),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_257),
.B(n_264),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_205),
.A2(n_195),
.B(n_176),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_225),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_234),
.C(n_217),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_208),
.A2(n_176),
.B(n_181),
.Y(n_264)
);

BUFx12_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_238),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_222),
.C(n_232),
.D(n_210),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_267),
.B(n_256),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_231),
.B1(n_204),
.B2(n_215),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_276),
.B1(n_278),
.B2(n_243),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_275),
.B(n_279),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_209),
.B1(n_212),
.B2(n_228),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_260),
.B1(n_239),
.B2(n_246),
.Y(n_296)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_228),
.B(n_236),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_223),
.B1(n_221),
.B2(n_213),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_227),
.B1(n_229),
.B2(n_214),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_219),
.B(n_230),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_288),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_189),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_241),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_233),
.C(n_181),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_249),
.C(n_237),
.Y(n_303)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_274),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_294),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_261),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_302),
.B1(n_270),
.B2(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_301),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_282),
.B1(n_285),
.B2(n_288),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_239),
.B1(n_240),
.B2(n_238),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_255),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_249),
.C(n_257),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_303),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_310),
.B(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_276),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_285),
.C(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_313),
.B(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_317),
.A2(n_292),
.B1(n_305),
.B2(n_270),
.Y(n_332)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_286),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_309),
.C(n_295),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_268),
.B1(n_280),
.B2(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_323),
.Y(n_333)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_325),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_283),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_262),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_329),
.C(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_249),
.C(n_291),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_317),
.A2(n_305),
.B1(n_292),
.B2(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_321),
.A2(n_285),
.B(n_275),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g350 ( 
.A(n_335),
.B(n_265),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_291),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_339),
.B(n_319),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_266),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_323),
.Y(n_342)
);

OAI221xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_316),
.B1(n_304),
.B2(n_313),
.C(n_318),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_341),
.B(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_345),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_339),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_315),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_327),
.B(n_324),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_348),
.B(n_352),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_333),
.A2(n_338),
.B1(n_336),
.B2(n_293),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_349),
.A2(n_343),
.B(n_334),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_265),
.Y(n_360)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_328),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_353),
.A2(n_356),
.B(n_325),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_293),
.B1(n_300),
.B2(n_289),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_332),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_359),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_346),
.A2(n_329),
.B(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_360),
.B(n_347),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_330),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_282),
.C(n_244),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_350),
.C(n_351),
.Y(n_363)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_363),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_365),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_188),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_262),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_259),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_355),
.A3(n_360),
.B1(n_266),
.B2(n_259),
.C1(n_263),
.C2(n_361),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_371),
.B(n_372),
.Y(n_377)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_365),
.A2(n_188),
.A3(n_201),
.B1(n_263),
.B2(n_266),
.C1(n_359),
.C2(n_366),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_188),
.C(n_201),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

AOI21x1_ASAP7_75t_SL g379 ( 
.A1(n_377),
.A2(n_375),
.B(n_376),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_375),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_380),
.Y(n_382)
);


endmodule