module real_jpeg_26208_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_354, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_354;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_0),
.A2(n_47),
.B1(n_61),
.B2(n_64),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_0),
.A2(n_47),
.B1(n_76),
.B2(n_85),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_5),
.B(n_87),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_30),
.C(n_42),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_70),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_27),
.B1(n_169),
.B2(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_SL g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_7),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_7),
.A2(n_35),
.B1(n_61),
.B2(n_64),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_7),
.A2(n_35),
.B1(n_258),
.B2(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_57),
.B1(n_61),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_57),
.B1(n_85),
.B2(n_258),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_10),
.A2(n_38),
.B1(n_61),
.B2(n_64),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_10),
.A2(n_38),
.B1(n_75),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_11),
.A2(n_61),
.B1(n_64),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_72),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_11),
.A2(n_72),
.B1(n_84),
.B2(n_85),
.Y(n_234)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_12),
.B(n_64),
.C(n_82),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_84),
.B1(n_85),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_13),
.A2(n_61),
.B1(n_64),
.B2(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_90),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_90),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_346),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_333),
.B(n_345),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_296),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_354),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_269),
.B(n_295),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_240),
.B(n_268),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_131),
.B(n_219),
.C(n_239),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_115),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_23),
.B(n_115),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_91),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_25),
.B(n_54),
.C(n_91),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_26),
.B(n_39),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_27),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_27),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_27),
.A2(n_36),
.B(n_151),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_27),
.A2(n_151),
.B(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_28),
.A2(n_34),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_28),
.B(n_37),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_123),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_31),
.Y(n_170)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_48),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_40),
.A2(n_50),
.B1(n_144),
.B2(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_40),
.B(n_77),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_40),
.A2(n_50),
.B(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_43),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_44),
.A2(n_68),
.B(n_185),
.C(n_187),
.Y(n_184)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_45),
.B(n_139),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_64),
.C(n_67),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_48),
.B(n_209),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_56),
.B(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_49),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_49),
.A2(n_142),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_49),
.A2(n_142),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_50),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_50),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_73),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_56),
.B(n_142),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_56),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_59)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_64),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_74),
.B(n_80),
.C(n_113),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_61),
.B(n_77),
.CON(n_186),
.SN(n_186)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_65),
.A2(n_70),
.B1(n_129),
.B2(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_65),
.A2(n_102),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_65),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_65),
.A2(n_70),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_65),
.A2(n_236),
.B(n_276),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_65),
.A2(n_70),
.B(n_102),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_69),
.A2(n_100),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_69),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_69),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_78),
.B1(n_87),
.B2(n_88),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.CON(n_74),
.SN(n_74)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_75),
.Y(n_258)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_76),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_77),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_78),
.A2(n_87),
.B1(n_97),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_78),
.B(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_78),
.A2(n_87),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_78),
.A2(n_321),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_89),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_79),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_86),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_87),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_87),
.B(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_103),
.B2(n_114),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_94),
.B(n_98),
.C(n_114),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_95),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_95),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_101),
.B(n_262),
.Y(n_318)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_105),
.B1(n_112),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_116),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_120),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_127),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_124),
.B(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_218),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_213),
.B(n_217),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_197),
.B(n_212),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_180),
.B(n_196),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_158),
.B(n_179),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_140),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_153),
.C(n_156),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_165),
.B(n_178),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_171),
.B(n_177),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_191),
.C(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.C(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_230),
.C(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_242),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_267),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_251),
.B1(n_265),
.B2(n_266),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_266),
.C(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_250),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_246),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_245),
.A2(n_280),
.B(n_284),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_259),
.C(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B1(n_260),
.B2(n_264),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_256),
.B(n_302),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_271),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_279),
.B1(n_290),
.B2(n_291),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_277),
.B(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_278),
.A2(n_298),
.B1(n_310),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_290),
.C(n_294),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_289),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_312),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_312),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_310),
.C(n_311),
.Y(n_297)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_300),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_305),
.C(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_315),
.C(n_325),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_317),
.C(n_319),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_325),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_341),
.C(n_343),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_352),
.Y(n_351)
);


endmodule