module fake_jpeg_24773_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_15),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_20),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_36),
.B(n_13),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_17),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_12),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_23),
.B1(n_19),
.B2(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_53),
.B1(n_40),
.B2(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_32),
.Y(n_54)
);

OA21x2_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_43),
.B(n_39),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_41),
.C(n_38),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_60),
.C(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_45),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_30),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_40),
.B(n_28),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_49),
.C(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_44),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_30),
.B(n_33),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_65),
.B1(n_55),
.B2(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_60),
.B1(n_33),
.B2(n_29),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_70),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.C(n_29),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_69),
.B(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_17),
.B1(n_16),
.B2(n_3),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B1(n_14),
.B2(n_73),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_71),
.C(n_4),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.C(n_76),
.Y(n_78)
);


endmodule