module fake_jpeg_31076_n_519 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_60),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_73),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_2),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_32),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_93),
.Y(n_129)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_87),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_18),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_18),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_32),
.B(n_3),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_18),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_26),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_23),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_29),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_49),
.Y(n_145)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_42),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_145),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_146),
.Y(n_171)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_154),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_95),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_42),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_60),
.B(n_52),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_160),
.Y(n_201)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_81),
.B(n_49),
.Y(n_160)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_45),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_175),
.B(n_178),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_45),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_48),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_183),
.Y(n_237)
);

CKINVDCx12_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_48),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_29),
.B1(n_74),
.B2(n_85),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_194),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_56),
.B1(n_77),
.B2(n_101),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_190),
.B1(n_195),
.B2(n_210),
.Y(n_223)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_197),
.Y(n_234)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_62),
.B1(n_102),
.B2(n_65),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_29),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_216),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_41),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_100),
.B1(n_92),
.B2(n_78),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_34),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

CKINVDCx9p33_ASAP7_75t_R g202 ( 
.A(n_130),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_129),
.B(n_34),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_33),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_33),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_50),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_131),
.A2(n_68),
.B1(n_43),
.B2(n_36),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_211),
.B(n_166),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_165),
.A2(n_53),
.B1(n_104),
.B2(n_79),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_215),
.B1(n_131),
.B2(n_128),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_133),
.A2(n_64),
.B1(n_43),
.B2(n_39),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_121),
.A2(n_23),
.B(n_51),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

CKINVDCx9p33_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_219),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_21),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_222),
.B(n_50),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_21),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_228),
.C(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_128),
.C(n_139),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_206),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_243),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_174),
.B(n_127),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_246),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_192),
.A2(n_133),
.B1(n_162),
.B2(n_151),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_168),
.B1(n_162),
.B2(n_107),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_214),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_204),
.C(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_255),
.B(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_188),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_260),
.Y(n_321)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_216),
.B1(n_121),
.B2(n_219),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_199),
.B1(n_245),
.B2(n_143),
.Y(n_303)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_273),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_283),
.B1(n_247),
.B2(n_231),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_198),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_282),
.C(n_286),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_253),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_224),
.A2(n_218),
.B(n_217),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_288),
.B(n_248),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_282),
.Y(n_305)
);

OR2x2_ASAP7_75t_SL g276 ( 
.A(n_224),
.B(n_172),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_284),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_182),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_172),
.C(n_139),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_132),
.C(n_123),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_257),
.Y(n_318)
);

NAND2x1_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_202),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_182),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_291),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g350 ( 
.A1(n_294),
.A2(n_270),
.B1(n_280),
.B2(n_269),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_226),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_297),
.B(n_322),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_298),
.A2(n_312),
.B(n_288),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_229),
.B1(n_223),
.B2(n_193),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_301),
.A2(n_314),
.B1(n_268),
.B2(n_263),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_242),
.C(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_306),
.C(n_310),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_286),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_232),
.C(n_256),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_223),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_245),
.B1(n_168),
.B2(n_220),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_320),
.B1(n_287),
.B2(n_250),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_256),
.B(n_227),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_276),
.A2(n_148),
.B1(n_111),
.B2(n_108),
.Y(n_314)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_257),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_285),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_200),
.B1(n_177),
.B2(n_170),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_289),
.B(n_51),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_335),
.C(n_343),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_330),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_313),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_328),
.Y(n_356)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

A2O1A1O1Ixp25_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_307),
.B(n_319),
.C(n_308),
.D(n_312),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_51),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_336),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_301),
.A2(n_310),
.B1(n_298),
.B2(n_295),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_342),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_274),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_259),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_261),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_346),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_338),
.A2(n_347),
.B(n_304),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_262),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_339),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_262),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_340),
.B(n_339),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_265),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_350),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_309),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_307),
.A2(n_294),
.B(n_300),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_266),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_351),
.Y(n_378)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_353),
.A2(n_213),
.B(n_24),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_349),
.A2(n_315),
.B1(n_264),
.B2(n_299),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_370),
.B1(n_250),
.B2(n_196),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_332),
.A2(n_293),
.B1(n_316),
.B2(n_311),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_359),
.A2(n_324),
.B1(n_332),
.B2(n_325),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_351),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_364),
.Y(n_384)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_340),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_322),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_367),
.B(n_383),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_342),
.B(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_352),
.A2(n_315),
.B1(n_302),
.B2(n_125),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_382),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_345),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_350),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_278),
.Y(n_379)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_338),
.A2(n_334),
.B(n_339),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_381),
.A2(n_161),
.B(n_209),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_213),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_385),
.A2(n_394),
.B1(n_395),
.B2(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_360),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_388),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_343),
.C(n_344),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_390),
.C(n_396),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_344),
.C(n_335),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_375),
.A2(n_353),
.B(n_364),
.C(n_381),
.Y(n_391)
);

AO21x1_ASAP7_75t_L g420 ( 
.A1(n_391),
.A2(n_397),
.B(n_405),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_347),
.B1(n_331),
.B2(n_348),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_254),
.C(n_279),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_213),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_406),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_401),
.A2(n_403),
.B(n_357),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_378),
.A2(n_365),
.B(n_369),
.Y(n_403)
);

AO22x1_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_284),
.B1(n_251),
.B2(n_241),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_254),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_408),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_380),
.A2(n_170),
.B1(n_251),
.B2(n_148),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_191),
.C(n_161),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_362),
.C(n_361),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_363),
.B1(n_378),
.B2(n_375),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_412),
.A2(n_417),
.B1(n_421),
.B2(n_196),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_367),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_415),
.B(n_418),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_376),
.B1(n_356),
.B2(n_373),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_384),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_405),
.A2(n_371),
.B1(n_383),
.B2(n_357),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_398),
.B(n_369),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_434),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_433),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_393),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_5),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g429 ( 
.A(n_398),
.B(n_358),
.CI(n_354),
.CON(n_429),
.SN(n_429)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_429),
.B(n_410),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_358),
.C(n_354),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_396),
.C(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_24),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_372),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_406),
.B(n_372),
.Y(n_434)
);

AO32x1_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_391),
.A3(n_399),
.B1(n_400),
.B2(n_387),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_437),
.Y(n_455)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

INVx13_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_443),
.C(n_449),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_409),
.B1(n_411),
.B2(n_391),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_425),
.B1(n_419),
.B2(n_432),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_391),
.C(n_372),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_397),
.B(n_6),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_445),
.A2(n_412),
.B(n_421),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_447),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_23),
.Y(n_448)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_111),
.C(n_140),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_417),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_450),
.B(n_451),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_24),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_420),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_461),
.A2(n_466),
.B1(n_31),
.B2(n_138),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_468),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_444),
.B(n_433),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_467),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_416),
.C(n_424),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_470),
.C(n_449),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_429),
.B1(n_422),
.B2(n_434),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_443),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_173),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_439),
.A2(n_196),
.B(n_137),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_469),
.A2(n_445),
.B(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_97),
.C(n_173),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_456),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_472),
.B(n_474),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_454),
.A2(n_435),
.B1(n_438),
.B2(n_437),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_39),
.C(n_114),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_465),
.B(n_452),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_475),
.B(n_478),
.Y(n_496)
);

AOI21xp33_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_447),
.B(n_453),
.Y(n_477)
);

AOI31xp67_ASAP7_75t_L g492 ( 
.A1(n_477),
.A2(n_480),
.A3(n_483),
.B(n_485),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_459),
.B(n_39),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_479),
.A2(n_480),
.B1(n_482),
.B2(n_464),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_459),
.A2(n_137),
.B(n_138),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_5),
.B(n_8),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_457),
.A2(n_158),
.B(n_122),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_485),
.A2(n_30),
.B(n_9),
.Y(n_495)
);

OA21x2_ASAP7_75t_SL g486 ( 
.A1(n_476),
.A2(n_467),
.B(n_468),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_492),
.B(n_493),
.Y(n_502)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_487),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_495),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_479),
.A2(n_458),
.B1(n_470),
.B2(n_122),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_490),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_39),
.C(n_108),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_497),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_481),
.B(n_9),
.C(n_10),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_SL g508 ( 
.A(n_500),
.B(n_495),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_114),
.C(n_31),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_504),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_497),
.A2(n_46),
.B1(n_30),
.B2(n_11),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_505),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_509),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_508),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_498),
.A2(n_503),
.B(n_496),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_46),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_504),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_513),
.B(n_506),
.C(n_46),
.Y(n_515)
);

AO21x1_ASAP7_75t_SL g514 ( 
.A1(n_512),
.A2(n_502),
.B(n_511),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g516 ( 
.A1(n_514),
.A2(n_515),
.A3(n_8),
.B1(n_10),
.B2(n_12),
.C(n_31),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_516),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_10),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_12),
.B(n_500),
.Y(n_519)
);


endmodule