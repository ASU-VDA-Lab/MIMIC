module fake_jpeg_28425_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_13),
.Y(n_19)
);

OR2x2_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_13),
.B1(n_12),
.B2(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_16),
.B1(n_15),
.B2(n_9),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_28),
.B1(n_15),
.B2(n_9),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_33),
.Y(n_44)
);

OAI31xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_32),
.A3(n_21),
.B(n_14),
.Y(n_41)
);

AOI32xp33_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_21),
.A3(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_30),
.B1(n_32),
.B2(n_18),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_20),
.C(n_26),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.C(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_11),
.B1(n_26),
.B2(n_3),
.Y(n_54)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_14),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_54),
.B1(n_46),
.B2(n_41),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_34),
.B(n_2),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_51),
.B(n_44),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_39),
.C(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_11),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_46),
.C(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_44),
.B1(n_39),
.B2(n_40),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_45),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_53),
.B(n_26),
.Y(n_67)
);

OAI322xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_11),
.A3(n_53),
.B1(n_8),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_61),
.B1(n_3),
.B2(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_2),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_61),
.Y(n_71)
);

OAI211xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B(n_70),
.C(n_3),
.Y(n_73)
);

NAND4xp25_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_71),
.C(n_5),
.D(n_6),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_2),
.Y(n_75)
);


endmodule