module fake_jpeg_4547_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_27),
.B1(n_17),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_60),
.B1(n_42),
.B2(n_39),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_26),
.B(n_30),
.C(n_18),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_24),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_22),
.C(n_34),
.Y(n_73)
);

NAND2x1_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_60),
.B1(n_52),
.B2(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_91),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_40),
.B1(n_43),
.B2(n_22),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_87),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_40),
.C(n_37),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_53),
.C(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_43),
.B1(n_33),
.B2(n_34),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_66),
.B1(n_61),
.B2(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_52),
.Y(n_111)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_64),
.B1(n_66),
.B2(n_58),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_113),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_104),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_45),
.B1(n_51),
.B2(n_49),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_92),
.B(n_45),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_109),
.B(n_116),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_47),
.B1(n_56),
.B2(n_55),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_46),
.B1(n_43),
.B2(n_48),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_81),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_73),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_52),
.B(n_48),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_70),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_81),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_123),
.B(n_35),
.C(n_34),
.Y(n_179)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_126),
.Y(n_158)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_98),
.CI(n_105),
.CON(n_127),
.SN(n_127)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_149),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_74),
.B1(n_75),
.B2(n_88),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_50),
.B1(n_70),
.B2(n_87),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_94),
.B1(n_74),
.B2(n_93),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_144),
.B1(n_119),
.B2(n_87),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_88),
.B1(n_82),
.B2(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_148),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_113),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_71),
.B1(n_95),
.B2(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_103),
.B(n_50),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_101),
.B1(n_106),
.B2(n_108),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_137),
.B1(n_144),
.B2(n_150),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_149),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_164),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_139),
.CI(n_143),
.CON(n_156),
.SN(n_156)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_157),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_104),
.Y(n_163)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_37),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_35),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_178),
.B(n_179),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_35),
.CI(n_86),
.CON(n_168),
.SN(n_168)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_181),
.B(n_178),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_103),
.B1(n_21),
.B2(n_29),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_76),
.B(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_183),
.B1(n_129),
.B2(n_124),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_128),
.A2(n_25),
.B(n_31),
.C(n_29),
.D(n_50),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_160),
.B1(n_168),
.B2(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_130),
.B(n_135),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_196),
.B(n_198),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_205),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_130),
.B(n_147),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_209),
.B(n_183),
.C(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_201),
.B1(n_181),
.B2(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_126),
.B1(n_21),
.B2(n_31),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_161),
.B(n_175),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_225),
.B(n_229),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_166),
.B(n_156),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_164),
.B1(n_156),
.B2(n_166),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_216),
.B1(n_224),
.B2(n_8),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_220),
.B1(n_233),
.B2(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_155),
.C(n_168),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_200),
.C(n_184),
.Y(n_236)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_221),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_31),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_29),
.B(n_25),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_31),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_29),
.B1(n_25),
.B2(n_31),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_25),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_190),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_238),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_254),
.B1(n_233),
.B2(n_226),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_198),
.C(n_196),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_244),
.C(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_202),
.C(n_187),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_193),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_210),
.B1(n_204),
.B2(n_203),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_246),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_0),
.C(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_10),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_8),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_11),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_215),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_231),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_215),
.B1(n_222),
.B2(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_215),
.B1(n_225),
.B2(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

AOI221xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_242),
.B1(n_240),
.B2(n_250),
.C(n_253),
.Y(n_279)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_266),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_225),
.B1(n_228),
.B2(n_231),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_217),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_7),
.B(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_0),
.C(n_1),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_7),
.C(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_238),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_280),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_240),
.Y(n_280)
);

OAI322xp33_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_243),
.A3(n_11),
.B1(n_4),
.B2(n_6),
.C1(n_7),
.C2(n_16),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_269),
.C(n_271),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_287),
.B1(n_268),
.B2(n_283),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_275),
.B(n_284),
.C(n_264),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_277),
.B1(n_257),
.B2(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_4),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_268),
.C(n_276),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_297),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_302),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_4),
.B1(n_6),
.B2(n_12),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_0),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_293),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_289),
.B1(n_291),
.B2(n_13),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_309),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

AOI32xp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_305),
.A3(n_311),
.B1(n_13),
.B2(n_16),
.Y(n_315)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_2),
.A3(n_12),
.B1(n_295),
.B2(n_309),
.C(n_282),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_12),
.CI(n_2),
.CON(n_317),
.SN(n_317)
);


endmodule