module real_aes_7804_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_363;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_756;
wire n_288;
wire n_598;
wire n_404;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_385;
wire n_275;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_0), .A2(n_149), .B1(n_619), .B2(n_621), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_1), .A2(n_38), .B1(n_382), .B2(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_2), .A2(n_228), .B1(n_531), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_3), .A2(n_177), .B1(n_775), .B2(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_4), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_5), .A2(n_235), .B1(n_378), .B2(n_380), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_6), .A2(n_27), .B1(n_104), .B2(n_366), .C1(n_492), .C2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_7), .A2(n_29), .B1(n_426), .B2(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_8), .A2(n_106), .B1(n_375), .B2(n_382), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_9), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_10), .A2(n_111), .B1(n_417), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_11), .A2(n_183), .B1(n_324), .B2(n_330), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_12), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_13), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_14), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_15), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_16), .B(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_17), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_18), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_19), .A2(n_191), .B1(n_569), .B2(n_571), .C(n_572), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_20), .A2(n_37), .B1(n_589), .B2(n_591), .C(n_592), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_21), .A2(n_128), .B1(n_623), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_22), .A2(n_182), .B1(n_346), .B2(n_402), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_23), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_24), .Y(n_694) );
AO22x2_ASAP7_75t_L g263 ( .A1(n_25), .A2(n_73), .B1(n_264), .B2(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g750 ( .A(n_25), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_26), .A2(n_63), .B1(n_335), .B2(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_28), .A2(n_61), .B1(n_339), .B2(n_579), .C(n_582), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_30), .A2(n_229), .B1(n_344), .B2(n_426), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_31), .A2(n_136), .B1(n_319), .B2(n_439), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_32), .A2(n_202), .B1(n_319), .B2(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_33), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_34), .A2(n_754), .B1(n_778), .B2(n_779), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_34), .Y(n_778) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_35), .A2(n_166), .B1(n_474), .B2(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_36), .Y(n_715) );
AO22x2_ASAP7_75t_L g267 ( .A1(n_39), .A2(n_78), .B1(n_264), .B2(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g751 ( .A(n_39), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_40), .A2(n_84), .B1(n_382), .B2(n_680), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_41), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_42), .A2(n_216), .B1(n_680), .B2(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_43), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_44), .A2(n_167), .B1(n_346), .B2(n_373), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_45), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_46), .A2(n_181), .B1(n_429), .B2(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_47), .A2(n_70), .B1(n_337), .B2(n_346), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_48), .A2(n_133), .B1(n_140), .B2(n_284), .C1(n_405), .C2(n_623), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_49), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_50), .A2(n_137), .B1(n_366), .B2(n_655), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_51), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_52), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_53), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_54), .A2(n_68), .B1(n_289), .B2(n_296), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_55), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_56), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_57), .A2(n_109), .B1(n_424), .B2(n_425), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_58), .A2(n_116), .B1(n_367), .B2(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_59), .Y(n_642) );
XNOR2x2_ASAP7_75t_L g601 ( .A(n_60), .B(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_62), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_64), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_65), .A2(n_194), .B1(n_296), .B2(n_405), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_66), .A2(n_72), .B1(n_335), .B2(n_346), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_67), .A2(n_163), .B1(n_373), .B2(n_375), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_69), .A2(n_131), .B1(n_450), .B2(n_452), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_71), .A2(n_134), .B1(n_342), .B2(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_74), .Y(n_305) );
AOI222xp33_ASAP7_75t_L g733 ( .A1(n_75), .A2(n_77), .B1(n_108), .B2(n_284), .C1(n_452), .C2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_76), .A2(n_123), .B1(n_590), .B2(n_765), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_79), .A2(n_567), .B1(n_599), .B2(n_600), .Y(n_566) );
INVx1_ASAP7_75t_L g599 ( .A(n_79), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_80), .A2(n_224), .B1(n_290), .B2(n_545), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_81), .Y(n_696) );
INVx1_ASAP7_75t_L g247 ( .A(n_82), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_83), .A2(n_165), .B1(n_470), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_85), .A2(n_222), .B1(n_428), .B2(n_474), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_86), .A2(n_237), .B1(n_528), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_87), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_88), .A2(n_461), .B1(n_503), .B2(n_504), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_88), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_89), .Y(n_685) );
INVx1_ASAP7_75t_L g245 ( .A(n_90), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_91), .A2(n_208), .B1(n_611), .B2(n_612), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_92), .A2(n_114), .B1(n_297), .B2(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_93), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_94), .A2(n_232), .B1(n_297), .B2(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_95), .A2(n_203), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_96), .A2(n_164), .B1(n_611), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_97), .A2(n_209), .B1(n_659), .B2(n_660), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_98), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_99), .A2(n_103), .B1(n_361), .B2(n_523), .Y(n_522) );
OA22x2_ASAP7_75t_L g506 ( .A1(n_100), .A2(n_507), .B1(n_508), .B2(n_533), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_100), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_101), .B(n_408), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_102), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_105), .B(n_519), .Y(n_518) );
OA22x2_ASAP7_75t_L g534 ( .A1(n_107), .A2(n_535), .B1(n_536), .B2(n_557), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_107), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_110), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_112), .A2(n_121), .B1(n_659), .B2(n_660), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_113), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_115), .A2(n_141), .B1(n_683), .B2(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_117), .A2(n_221), .B1(n_470), .B2(n_614), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_118), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_119), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_120), .B(n_671), .Y(n_670) );
XNOR2x2_ASAP7_75t_L g630 ( .A(n_122), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g248 ( .A(n_124), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_125), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_126), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_127), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_129), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_130), .B(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_132), .A2(n_135), .B1(n_607), .B2(n_608), .Y(n_606) );
AND2x6_ASAP7_75t_L g244 ( .A(n_138), .B(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_138), .Y(n_744) );
AO22x2_ASAP7_75t_L g273 ( .A1(n_139), .A2(n_192), .B1(n_264), .B2(n_268), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_142), .A2(n_162), .B1(n_335), .B2(n_339), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_143), .A2(n_171), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_144), .A2(n_196), .B1(n_485), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_145), .A2(n_204), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_146), .A2(n_219), .B1(n_373), .B2(n_429), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_147), .A2(n_234), .B1(n_771), .B2(n_772), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_148), .A2(n_180), .B1(n_344), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g348 ( .A(n_150), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_151), .A2(n_195), .B1(n_362), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_152), .A2(n_206), .B1(n_428), .B2(n_430), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_153), .A2(n_225), .B1(n_342), .B2(n_375), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_154), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_155), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_156), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_157), .B(n_656), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_158), .A2(n_213), .B1(n_440), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_159), .A2(n_186), .B1(n_468), .B2(n_470), .Y(n_467) );
AO22x2_ASAP7_75t_L g271 ( .A1(n_160), .A2(n_210), .B1(n_264), .B2(n_265), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_161), .Y(n_300) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_168), .A2(n_193), .B1(n_326), .B2(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_169), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_170), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_172), .A2(n_212), .B1(n_405), .B2(n_458), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_173), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_174), .A2(n_205), .B1(n_316), .B2(n_635), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_175), .A2(n_178), .B1(n_637), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_176), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_179), .Y(n_480) );
INVx1_ASAP7_75t_L g616 ( .A(n_184), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_185), .A2(n_218), .B1(n_316), .B2(n_319), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_187), .A2(n_223), .B1(n_296), .B2(n_361), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g239 ( .A1(n_188), .A2(n_240), .B(n_249), .C(n_752), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_189), .B(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_190), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_192), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g788 ( .A(n_197), .Y(n_788) );
OA22x2_ASAP7_75t_L g789 ( .A1(n_197), .A2(n_755), .B1(n_756), .B2(n_788), .Y(n_789) );
INVx1_ASAP7_75t_L g435 ( .A(n_198), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_199), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_200), .B(n_519), .Y(n_617) );
INVx1_ASAP7_75t_L g385 ( .A(n_201), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_207), .Y(n_573) );
INVx1_ASAP7_75t_L g747 ( .A(n_210), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_211), .A2(n_230), .B1(n_344), .B2(n_346), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_214), .A2(n_220), .B1(n_382), .B2(n_485), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_215), .Y(n_667) );
XNOR2x2_ASAP7_75t_L g717 ( .A(n_217), .B(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_226), .Y(n_403) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_227), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_231), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_233), .Y(n_281) );
AOI22x1_ASAP7_75t_L g393 ( .A1(n_236), .A2(n_394), .B1(n_431), .B2(n_432), .Y(n_393) );
INVx1_ASAP7_75t_L g431 ( .A(n_236), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_238), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_245), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_246), .A2(n_742), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_561), .B1(n_737), .B2(n_738), .C(n_739), .Y(n_249) );
INVx1_ASAP7_75t_L g737 ( .A(n_250), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B1(n_386), .B2(n_387), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
XNOR2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_349), .Y(n_252) );
XOR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_348), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_313), .Y(n_254) );
NOR3xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_280), .C(n_299), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B1(n_274), .B2(n_275), .Y(n_256) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g398 ( .A(n_259), .Y(n_398) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g354 ( .A(n_260), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_260), .A2(n_277), .B1(n_447), .B2(n_448), .C(n_449), .Y(n_446) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_260), .Y(n_500) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
INVx2_ASAP7_75t_L g338 ( .A(n_261), .Y(n_338) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
AND2x2_ASAP7_75t_L g279 ( .A(n_262), .B(n_267), .Y(n_279) );
AND2x2_ASAP7_75t_L g318 ( .A(n_262), .B(n_294), .Y(n_318) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g285 ( .A(n_263), .B(n_267), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_263), .B(n_273), .Y(n_295) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g268 ( .A(n_266), .Y(n_268) );
INVx2_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
INVx1_ASAP7_75t_L g332 ( .A(n_267), .Y(n_332) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_270), .B(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g342 ( .A(n_270), .B(n_318), .Y(n_342) );
AND2x6_ASAP7_75t_L g517 ( .A(n_270), .B(n_279), .Y(n_517) );
AND2x4_ASAP7_75t_L g521 ( .A(n_270), .B(n_338), .Y(n_521) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g287 ( .A(n_271), .Y(n_287) );
INVx1_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
INVx1_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_271), .B(n_273), .Y(n_322) );
AND2x2_ASAP7_75t_L g286 ( .A(n_272), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g329 ( .A(n_273), .B(n_312), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_275), .A2(n_699), .B1(n_700), .B2(n_702), .Y(n_698) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g357 ( .A(n_278), .Y(n_357) );
AND2x2_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g345 ( .A(n_279), .B(n_286), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_279), .B(n_329), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_288), .Y(n_280) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_283), .A2(n_359), .B(n_360), .Y(n_358) );
INVx4_ASAP7_75t_L g492 ( .A(n_283), .Y(n_492) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
BUFx3_ASAP7_75t_L g455 ( .A(n_284), .Y(n_455) );
INVx2_ASAP7_75t_L g648 ( .A(n_284), .Y(n_648) );
INVx2_ASAP7_75t_L g666 ( .A(n_284), .Y(n_666) );
AND2x6_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
AND2x4_ASAP7_75t_L g362 ( .A(n_285), .B(n_311), .Y(n_362) );
AND2x2_ASAP7_75t_L g317 ( .A(n_286), .B(n_318), .Y(n_317) );
AND2x6_ASAP7_75t_L g337 ( .A(n_286), .B(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx4_ASAP7_75t_L g652 ( .A(n_290), .Y(n_652) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_291), .Y(n_367) );
BUFx4f_ASAP7_75t_SL g405 ( .A(n_291), .Y(n_405) );
BUFx2_ASAP7_75t_L g553 ( .A(n_291), .Y(n_553) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
INVx1_ASAP7_75t_L g304 ( .A(n_294), .Y(n_304) );
AND2x4_ASAP7_75t_L g297 ( .A(n_295), .B(n_298), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g450 ( .A(n_295), .B(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g497 ( .A(n_296), .Y(n_497) );
INVx2_ASAP7_75t_L g735 ( .A(n_296), .Y(n_735) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_297), .Y(n_408) );
BUFx12f_ASAP7_75t_L g458 ( .A(n_297), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_305), .B2(n_306), .Y(n_299) );
INVx3_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g594 ( .A(n_302), .Y(n_594) );
INVx4_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_303), .A2(n_364), .B1(n_365), .B2(n_368), .Y(n_363) );
BUFx3_ASAP7_75t_L g411 ( .A(n_303), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_303), .A2(n_306), .B1(n_488), .B2(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_L g442 ( .A(n_304), .B(n_321), .Y(n_442) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g596 ( .A(n_307), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g413 ( .A(n_308), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_308), .A2(n_331), .B1(n_547), .B2(n_548), .Y(n_546) );
OR2x6_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_333), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_323), .Y(n_314) );
BUFx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_317), .Y(n_732) );
AND2x4_ASAP7_75t_L g320 ( .A(n_318), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g347 ( .A(n_318), .B(n_329), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_318), .B(n_329), .Y(n_478) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g375 ( .A(n_320), .Y(n_375) );
BUFx3_ASAP7_75t_L g421 ( .A(n_320), .Y(n_421) );
BUFx3_ASAP7_75t_L g485 ( .A(n_320), .Y(n_485) );
BUFx3_ASAP7_75t_L g571 ( .A(n_320), .Y(n_571) );
BUFx3_ASAP7_75t_L g608 ( .A(n_320), .Y(n_608) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_320), .Y(n_635) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x6_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_326), .Y(n_637) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g380 ( .A(n_327), .Y(n_380) );
INVx5_ASAP7_75t_L g429 ( .A(n_327), .Y(n_429) );
INVx1_ASAP7_75t_L g469 ( .A(n_327), .Y(n_469) );
INVx2_ASAP7_75t_L g614 ( .A(n_327), .Y(n_614) );
BUFx3_ASAP7_75t_L g678 ( .A(n_327), .Y(n_678) );
INVx8_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx6_ASAP7_75t_SL g384 ( .A(n_331), .Y(n_384) );
INVx1_ASAP7_75t_SL g528 ( .A(n_331), .Y(n_528) );
INVx1_ASAP7_75t_L g451 ( .A(n_332), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_343), .Y(n_333) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx4_ASAP7_75t_L g440 ( .A(n_336), .Y(n_440) );
OAI21xp33_ASAP7_75t_SL g542 ( .A1(n_336), .A2(n_543), .B(n_544), .Y(n_542) );
INVx4_ASAP7_75t_L g683 ( .A(n_336), .Y(n_683) );
INVx11_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx11_ASAP7_75t_L g466 ( .A(n_337), .Y(n_466) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g607 ( .A(n_340), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_340), .A2(n_639), .B1(n_640), .B2(n_642), .Y(n_638) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
BUFx3_ASAP7_75t_L g482 ( .A(n_342), .Y(n_482) );
BUFx3_ASAP7_75t_L g714 ( .A(n_342), .Y(n_714) );
INVx2_ASAP7_75t_L g724 ( .A(n_342), .Y(n_724) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx6_ASAP7_75t_L g379 ( .A(n_345), .Y(n_379) );
BUFx3_ASAP7_75t_L g424 ( .A(n_345), .Y(n_424) );
BUFx3_ASAP7_75t_L g585 ( .A(n_345), .Y(n_585) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g426 ( .A(n_347), .Y(n_426) );
BUFx3_ASAP7_75t_L g612 ( .A(n_347), .Y(n_612) );
BUFx3_ASAP7_75t_L g730 ( .A(n_347), .Y(n_730) );
XOR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_385), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_369), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_358), .C(n_363), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_355), .B2(n_356), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_354), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_356), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_396) );
OA211x2_ASAP7_75t_L g615 ( .A1(n_356), .A2(n_616), .B(n_617), .C(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g502 ( .A(n_357), .Y(n_502) );
INVx1_ASAP7_75t_SL g541 ( .A(n_357), .Y(n_541) );
BUFx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_362), .Y(n_452) );
BUFx2_ASAP7_75t_SL g621 ( .A(n_362), .Y(n_621) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g494 ( .A(n_366), .Y(n_494) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g705 ( .A(n_367), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_376), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g439 ( .A(n_374), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g474 ( .A(n_379), .Y(n_474) );
INVx3_ASAP7_75t_L g531 ( .A(n_379), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_379), .A2(n_587), .B1(n_644), .B2(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g721 ( .A(n_379), .Y(n_721) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx4f_ASAP7_75t_SL g430 ( .A(n_384), .Y(n_430) );
BUFx2_ASAP7_75t_L g470 ( .A(n_384), .Y(n_470) );
BUFx2_ASAP7_75t_L g680 ( .A(n_384), .Y(n_680) );
BUFx2_ASAP7_75t_L g772 ( .A(n_384), .Y(n_772) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_459), .B2(n_560), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_433), .B2(n_434), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g432 ( .A(n_394), .Y(n_432) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_414), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .C(n_409), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B1(n_404), .B2(n_406), .C(n_407), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g693 ( .A(n_402), .Y(n_693) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx4f_ASAP7_75t_L g623 ( .A(n_408), .Y(n_623) );
INVx1_ASAP7_75t_L g695 ( .A(n_408), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_411), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_422), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g570 ( .A(n_418), .Y(n_570) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_418), .Y(n_611) );
BUFx3_ASAP7_75t_L g775 ( .A(n_418), .Y(n_775) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
XNOR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NOR4xp75_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .C(n_446), .D(n_453), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_441), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_444), .B(n_445), .Y(n_443) );
BUFx3_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
BUFx2_ASAP7_75t_L g545 ( .A(n_450), .Y(n_545) );
INVx1_ASAP7_75t_L g620 ( .A(n_450), .Y(n_620) );
BUFx2_ASAP7_75t_L g763 ( .A(n_450), .Y(n_763) );
INVx1_ASAP7_75t_SL g657 ( .A(n_452), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_456), .B(n_457), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_454), .A2(n_511), .B(n_512), .Y(n_510) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx4f_ASAP7_75t_SL g598 ( .A(n_458), .Y(n_598) );
INVx2_ASAP7_75t_SL g560 ( .A(n_459), .Y(n_560) );
OA22x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_505), .B1(n_558), .B2(n_559), .Y(n_459) );
INVx1_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
INVx1_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_462), .B(n_486), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .C(n_479), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g581 ( .A(n_466), .Y(n_581) );
INVx2_ASAP7_75t_L g605 ( .A(n_466), .Y(n_605) );
INVx5_ASAP7_75t_SL g641 ( .A(n_466), .Y(n_641) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_466), .Y(n_769) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g577 ( .A(n_470), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_475), .B2(n_476), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g587 ( .A(n_477), .Y(n_587) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_483), .B2(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g776 ( .A(n_481), .Y(n_776) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR3xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_490), .C(n_498), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B1(n_494), .B2(n_495), .C(n_496), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g701 ( .A(n_500), .Y(n_701) );
INVx1_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
XOR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_534), .Y(n_505) );
INVx1_ASAP7_75t_L g533 ( .A(n_508), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_524), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .C(n_522), .Y(n_513) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_SL g765 ( .A(n_516), .Y(n_765) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
BUFx2_ASAP7_75t_L g660 ( .A(n_517), .Y(n_660) );
BUFx2_ASAP7_75t_L g671 ( .A(n_517), .Y(n_671) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_519), .Y(n_673) );
INVx5_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
INVx2_ASAP7_75t_L g659 ( .A(n_520), .Y(n_659) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g557 ( .A(n_536), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_549), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .C(n_546), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g738 ( .A(n_561), .Y(n_738) );
AOI22xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_686), .B1(n_687), .B2(n_736), .Y(n_561) );
INVx1_ASAP7_75t_L g736 ( .A(n_562), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B1(n_625), .B2(n_626), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B1(n_601), .B2(n_624), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g600 ( .A(n_567), .Y(n_600) );
AND4x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_578), .C(n_588), .D(n_597), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_576), .B2(n_577), .Y(n_572) );
BUFx2_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g624 ( .A(n_601), .Y(n_624) );
NAND4xp75_ASAP7_75t_L g602 ( .A(n_603), .B(n_609), .C(n_615), .D(n_622), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_614), .Y(n_771) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g655 ( .A(n_620), .Y(n_655) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_661), .B2(n_662), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_632), .B(n_646), .Y(n_631) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_638), .C(n_643), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_653), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B(n_650), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g758 ( .A1(n_648), .A2(n_759), .B(n_760), .Y(n_758) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_658), .Y(n_653) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
XOR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_685), .Y(n_662) );
NAND3x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_675), .C(n_681), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_669), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B(n_668), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .C(n_674), .Y(n_669) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B1(n_716), .B2(n_717), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
XOR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_715), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_707), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_698), .C(n_703), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_695), .B2(n_696), .C(n_697), .Y(n_692) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND4xp75_ASAP7_75t_L g718 ( .A(n_719), .B(n_725), .C(n_728), .D(n_733), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_726), .B(n_727), .Y(n_725) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
OR2x2_ASAP7_75t_SL g792 ( .A(n_741), .B(n_746), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_742), .Y(n_781) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_743), .B(n_784), .Y(n_787) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_744), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
OAI322xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_780), .A3(n_782), .B1(n_785), .B2(n_788), .C1(n_789), .C2(n_790), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_754), .Y(n_779) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
NAND3x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_766), .C(n_773), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
CKINVDCx16_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
endmodule