module fake_jpeg_10029_n_274 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_28),
.B(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_52),
.B1(n_33),
.B2(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_24),
.B1(n_25),
.B2(n_16),
.Y(n_52)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_24),
.B1(n_13),
.B2(n_33),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_13),
.B1(n_33),
.B2(n_15),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_30),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_29),
.C(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_51),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_23),
.B(n_15),
.C(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_29),
.B(n_30),
.C(n_35),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_35),
.B1(n_44),
.B2(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_59),
.B1(n_13),
.B2(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_38),
.B1(n_52),
.B2(n_75),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_30),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_82),
.C(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_89),
.Y(n_100)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_53),
.B1(n_39),
.B2(n_55),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_107),
.B1(n_108),
.B2(n_39),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_117),
.B1(n_84),
.B2(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_116),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_31),
.B1(n_37),
.B2(n_53),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_82),
.B1(n_79),
.B2(n_95),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_26),
.B(n_19),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_20),
.B(n_19),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_74),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_29),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_78),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_12),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_20),
.B(n_19),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_131),
.B(n_137),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_34),
.C(n_36),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_36),
.C(n_34),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_136),
.B1(n_114),
.B2(n_37),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_87),
.B1(n_65),
.B2(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_101),
.B1(n_103),
.B2(n_111),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_87),
.B1(n_94),
.B2(n_65),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_15),
.B(n_56),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_139),
.B1(n_98),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_99),
.B1(n_100),
.B2(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_151),
.B1(n_21),
.B2(n_16),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_145),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_150),
.B1(n_121),
.B2(n_122),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_148),
.B(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_134),
.B1(n_129),
.B2(n_132),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_127),
.B1(n_130),
.B2(n_124),
.Y(n_150)
);

NOR2x1_ASAP7_75t_R g151 ( 
.A(n_137),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_156),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_27),
.B(n_21),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_63),
.C(n_36),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_164),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_36),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_176),
.B1(n_178),
.B2(n_154),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_177),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_119),
.B1(n_126),
.B2(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_37),
.B1(n_31),
.B2(n_16),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_181),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_162),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_14),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_149),
.B1(n_145),
.B2(n_162),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_194),
.B1(n_198),
.B2(n_202),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_165),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_187),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_146),
.B1(n_160),
.B2(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_161),
.B1(n_157),
.B2(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_161),
.C(n_63),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_165),
.C(n_170),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_18),
.B1(n_9),
.B2(n_12),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_205),
.B1(n_177),
.B2(n_173),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_37),
.B1(n_31),
.B2(n_18),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_217),
.C(n_219),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_186),
.B1(n_166),
.B2(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_199),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_167),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_7),
.B(n_11),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_193),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_184),
.B1(n_178),
.B2(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_185),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_220),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_34),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_8),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_8),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_187),
.B(n_7),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_199),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_213),
.B(n_217),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_189),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_4),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_205),
.C(n_198),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_233),
.C(n_27),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_31),
.C(n_27),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_234),
.B(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_241),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_243),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_247),
.B1(n_10),
.B2(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_18),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_246),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_0),
.C(n_1),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_223),
.C(n_2),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_5),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_232),
.B1(n_228),
.B2(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_254),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_1),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_1),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_261),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_251),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_266),
.B(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_251),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_258),
.B(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_267),
.C(n_2),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_2),
.B(n_3),
.C(n_199),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_3),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_273),
.B(n_3),
.Y(n_274)
);


endmodule