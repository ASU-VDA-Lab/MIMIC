module fake_jpeg_28230_n_279 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_28),
.B1(n_18),
.B2(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_27),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_18),
.B(n_23),
.C(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_38),
.B1(n_51),
.B2(n_50),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_16),
.A3(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_68),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_42),
.B1(n_46),
.B2(n_41),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_31),
.A3(n_30),
.B1(n_26),
.B2(n_21),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_16),
.B1(n_26),
.B2(n_12),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_83),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_30),
.C(n_31),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_30),
.C(n_31),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_87),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_84),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_41),
.B1(n_48),
.B2(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_69),
.B1(n_53),
.B2(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_24),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_71),
.B1(n_55),
.B2(n_63),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_41),
.B1(n_48),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_87),
.B1(n_90),
.B2(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_97),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_92),
.B1(n_37),
.B2(n_22),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_85),
.B1(n_88),
.B2(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_105),
.B1(n_93),
.B2(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_72),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_84),
.B1(n_77),
.B2(n_83),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_63),
.B(n_55),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_109),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_115),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_78),
.C(n_94),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_63),
.B(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_26),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_26),
.A3(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_14),
.B(n_71),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_82),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_14),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_78),
.B(n_74),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_124),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_143),
.B1(n_106),
.B2(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_142),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_138),
.B1(n_144),
.B2(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_146),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_137),
.B(n_139),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_84),
.B1(n_74),
.B2(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_14),
.B(n_25),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_25),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_25),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_92),
.B1(n_37),
.B2(n_22),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_22),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_37),
.C(n_17),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_111),
.C(n_120),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_119),
.B1(n_99),
.B2(n_102),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_17),
.B1(n_13),
.B2(n_3),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_151),
.B1(n_105),
.B2(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_17),
.B1(n_13),
.B2(n_3),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_160),
.C(n_176),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_120),
.B(n_112),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_155),
.B1(n_165),
.B2(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_156),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_135),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_115),
.C(n_108),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_113),
.B(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_113),
.C(n_109),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_118),
.B(n_2),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_141),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_183),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_140),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_133),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_191),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_199),
.B1(n_201),
.B2(n_165),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_147),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_110),
.B1(n_13),
.B2(n_4),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_1),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_159),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_154),
.B1(n_157),
.B2(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_220),
.B1(n_189),
.B2(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_170),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_161),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_219),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_177),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_216),
.B1(n_3),
.B2(n_5),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_160),
.C(n_152),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_185),
.C(n_181),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_186),
.B(n_166),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_157),
.B1(n_155),
.B2(n_167),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_190),
.B1(n_199),
.B2(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_153),
.B1(n_166),
.B2(n_5),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_229),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_183),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_217),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_210),
.C(n_212),
.Y(n_242)
);

BUFx12f_ASAP7_75t_SL g226 ( 
.A(n_220),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_205),
.B(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_184),
.B1(n_194),
.B2(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_231),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_198),
.B1(n_4),
.B2(n_5),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_6),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_219),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_224),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_215),
.C(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_221),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_246),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_240),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_232),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_229),
.B1(n_232),
.B2(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_222),
.C(n_7),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_10),
.C(n_7),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_6),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_261),
.Y(n_265)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_251),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_260),
.B(n_262),
.Y(n_267)
);

NAND4xp25_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_256),
.C(n_255),
.D(n_249),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_267),
.A2(n_268),
.B1(n_6),
.B2(n_8),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_253),
.B(n_7),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_6),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.C(n_265),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.C(n_8),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_261),
.B(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_10),
.B(n_8),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_9),
.B(n_226),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_9),
.Y(n_279)
);


endmodule