module fake_netlist_1_12613_n_464 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_464);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_464;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g66 ( .A(n_11), .Y(n_66) );
CKINVDCx20_ASAP7_75t_R g67 ( .A(n_52), .Y(n_67) );
INVxp67_ASAP7_75t_SL g68 ( .A(n_18), .Y(n_68) );
CKINVDCx5p33_ASAP7_75t_R g69 ( .A(n_11), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_49), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_22), .Y(n_71) );
CKINVDCx16_ASAP7_75t_R g72 ( .A(n_57), .Y(n_72) );
INVxp67_ASAP7_75t_SL g73 ( .A(n_2), .Y(n_73) );
INVxp67_ASAP7_75t_L g74 ( .A(n_26), .Y(n_74) );
INVxp67_ASAP7_75t_L g75 ( .A(n_1), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_12), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_31), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_1), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_34), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_23), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_38), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_51), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_50), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_15), .B(n_24), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_35), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_14), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_55), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_54), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_14), .Y(n_96) );
INVx4_ASAP7_75t_R g97 ( .A(n_25), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_20), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_47), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_19), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_44), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_37), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_80), .B(n_0), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_72), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
NAND2xp33_ASAP7_75t_R g107 ( .A(n_80), .B(n_0), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
NOR2xp67_ASAP7_75t_L g111 ( .A(n_74), .B(n_3), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_96), .B(n_3), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_74), .B(n_4), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_86), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_86), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_103), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_96), .B(n_4), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_98), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_69), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_71), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_98), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_78), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_117), .B(n_66), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_114), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_114), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_117), .B(n_70), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_122), .A2(n_68), .B1(n_73), .B2(n_94), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_104), .B(n_79), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_117), .B(n_104), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_123), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_119), .A2(n_66), .B1(n_76), .B2(n_100), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_119), .B(n_79), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_114), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_108), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_116), .Y(n_152) );
OAI221xp5_ASAP7_75t_L g153 ( .A1(n_112), .A2(n_68), .B1(n_73), .B2(n_84), .C(n_75), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g154 ( .A1(n_132), .A2(n_104), .B(n_112), .C(n_101), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_131), .B(n_121), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_131), .B(n_116), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_149), .B(n_124), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_149), .B(n_131), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_136), .B(n_105), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_151), .A2(n_110), .B(n_101), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_151), .A2(n_110), .B(n_92), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_148), .A2(n_92), .B(n_89), .Y(n_162) );
NOR2xp33_ASAP7_75t_R g163 ( .A(n_152), .B(n_122), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_134), .B(n_125), .Y(n_164) );
OR2x2_ASAP7_75t_L g165 ( .A(n_133), .B(n_120), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_148), .A2(n_92), .B(n_93), .Y(n_166) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_142), .A2(n_82), .B(n_90), .Y(n_167) );
OR2x6_ASAP7_75t_SL g168 ( .A(n_152), .B(n_120), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_145), .A2(n_93), .B(n_89), .C(n_82), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_136), .B(n_132), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_128), .B(n_111), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_142), .A2(n_87), .B(n_99), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_142), .A2(n_90), .B(n_87), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_134), .A2(n_107), .B1(n_127), .B2(n_106), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_153), .A2(n_107), .B1(n_115), .B2(n_126), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_145), .A2(n_111), .B(n_113), .C(n_99), .Y(n_180) );
NOR2x1_ASAP7_75t_R g181 ( .A(n_128), .B(n_118), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_137), .A2(n_113), .B(n_76), .C(n_102), .Y(n_182) );
NOR3xp33_ASAP7_75t_SL g183 ( .A(n_133), .B(n_88), .C(n_102), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_142), .A2(n_88), .B(n_81), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_140), .B(n_85), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_165), .B(n_128), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_173), .A2(n_153), .B1(n_83), .B2(n_95), .Y(n_187) );
NAND2xp33_ASAP7_75t_L g188 ( .A(n_178), .B(n_150), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_163), .Y(n_189) );
AOI21x1_ASAP7_75t_L g190 ( .A1(n_167), .A2(n_138), .B(n_129), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_147), .B(n_130), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_171), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
AOI221xp5_ASAP7_75t_L g196 ( .A1(n_172), .A2(n_139), .B1(n_83), .B2(n_95), .C(n_100), .Y(n_196) );
BUFx2_ASAP7_75t_SL g197 ( .A(n_164), .Y(n_197) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_161), .A2(n_135), .B(n_147), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_164), .B(n_150), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
OAI21x1_ASAP7_75t_L g201 ( .A1(n_162), .A2(n_135), .B(n_147), .Y(n_201) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_170), .A2(n_138), .B(n_129), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_185), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_154), .A2(n_150), .B(n_137), .Y(n_204) );
OAI21x1_ASAP7_75t_L g205 ( .A1(n_166), .A2(n_130), .B(n_147), .Y(n_205) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_175), .A2(n_135), .B(n_130), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_174), .B(n_150), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_163), .Y(n_208) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_184), .A2(n_139), .B(n_138), .Y(n_209) );
INVx1_ASAP7_75t_SL g210 ( .A(n_169), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_158), .B(n_150), .Y(n_211) );
OAI21xp33_ASAP7_75t_SL g212 ( .A1(n_158), .A2(n_143), .B(n_141), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_155), .B(n_141), .Y(n_214) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_170), .A2(n_129), .B(n_144), .Y(n_215) );
OAI21x1_ASAP7_75t_SL g216 ( .A1(n_177), .A2(n_143), .B(n_135), .Y(n_216) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_185), .A2(n_130), .B(n_144), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_214), .B(n_159), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_213), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_186), .A2(n_174), .B1(n_157), .B2(n_156), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_212), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
NAND2xp33_ASAP7_75t_R g224 ( .A(n_208), .B(n_183), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_214), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_214), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_186), .B(n_157), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_204), .Y(n_228) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_217), .A2(n_180), .B(n_182), .Y(n_229) );
NOR2xp33_ASAP7_75t_R g230 ( .A(n_189), .B(n_126), .Y(n_230) );
NAND2xp33_ASAP7_75t_R g231 ( .A(n_186), .B(n_168), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_204), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_212), .B(n_179), .Y(n_233) );
INVx4_ASAP7_75t_SL g234 ( .A(n_193), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_140), .B(n_84), .C(n_75), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_210), .B(n_140), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_189), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_210), .B(n_140), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_197), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_207), .B(n_181), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_243), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_243), .Y(n_246) );
AND4x1_ASAP7_75t_L g247 ( .A(n_233), .B(n_196), .C(n_211), .D(n_197), .Y(n_247) );
OR2x6_ASAP7_75t_L g248 ( .A(n_221), .B(n_216), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_219), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_243), .A2(n_217), .B(n_216), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_225), .B(n_200), .Y(n_253) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_221), .A2(n_216), .B(n_217), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_243), .A2(n_198), .B(n_205), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_196), .B1(n_200), .B2(n_203), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_241), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_223), .Y(n_258) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_228), .A2(n_198), .B(n_201), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_222), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_236), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_231), .A2(n_200), .B1(n_203), .B2(n_187), .Y(n_263) );
AOI21xp5_ASAP7_75t_SL g264 ( .A1(n_240), .A2(n_191), .B(n_195), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_228), .A2(n_201), .B(n_205), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_233), .A2(n_202), .B(n_215), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_258), .B(n_227), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_249), .B(n_226), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_249), .B(n_226), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_245), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_247), .B(n_218), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_258), .B(n_234), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_258), .B(n_234), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_227), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_245), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_266), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_245), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_266), .B(n_232), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_266), .B(n_227), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_266), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_245), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_251), .B(n_234), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_251), .B(n_234), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_249), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_272), .B(n_246), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_288), .B(n_253), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_272), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_275), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_281), .B(n_246), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_279), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_280), .B(n_246), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_286), .B(n_263), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_275), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_275), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_284), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_274), .B(n_247), .C(n_231), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_288), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_285), .B(n_246), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_278), .B(n_248), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_273), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_270), .B(n_253), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_281), .B(n_248), .Y(n_311) );
AOI22x1_ASAP7_75t_L g312 ( .A1(n_287), .A2(n_240), .B1(n_237), .B2(n_257), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_289), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g316 ( .A(n_301), .B(n_230), .C(n_247), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_290), .B(n_250), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_303), .B(n_256), .Y(n_318) );
AOI221x1_ASAP7_75t_L g319 ( .A1(n_291), .A2(n_264), .B1(n_256), .B2(n_250), .C(n_276), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_297), .A2(n_224), .B1(n_242), .B2(n_218), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_304), .B(n_278), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_294), .A2(n_264), .B(n_275), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_294), .B(n_278), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_303), .B(n_270), .Y(n_325) );
NOR3xp33_ASAP7_75t_L g326 ( .A(n_295), .B(n_237), .C(n_187), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_312), .A2(n_235), .B(n_220), .Y(n_327) );
AOI31xp33_ASAP7_75t_L g328 ( .A1(n_293), .A2(n_287), .A3(n_286), .B(n_276), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_310), .B(n_269), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_311), .A2(n_248), .B1(n_287), .B2(n_286), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_296), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_296), .B(n_269), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_304), .B(n_285), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_311), .A2(n_248), .B1(n_283), .B2(n_277), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_302), .B(n_277), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_293), .A2(n_248), .B1(n_251), .B2(n_283), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_302), .B(n_282), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_298), .B(n_271), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_299), .Y(n_341) );
INVxp33_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_305), .A2(n_248), .B1(n_251), .B2(n_262), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_305), .A2(n_248), .B1(n_276), .B2(n_251), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_307), .A2(n_238), .B(n_236), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_333), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_308), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_331), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_331), .B(n_309), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_325), .B(n_313), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_321), .B(n_305), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_325), .B(n_282), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_316), .B(n_5), .Y(n_354) );
OAI22x1_ASAP7_75t_L g355 ( .A1(n_341), .A2(n_292), .B1(n_314), .B2(n_254), .Y(n_355) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_337), .B(n_314), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_320), .B(n_5), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_318), .B(n_282), .Y(n_358) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_327), .B(n_254), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_321), .B(n_334), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_324), .Y(n_361) );
NAND2xp33_ASAP7_75t_L g362 ( .A(n_326), .B(n_257), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_322), .B(n_257), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_324), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_334), .B(n_254), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_344), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_329), .B(n_261), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_343), .A2(n_262), .B1(n_203), .B2(n_267), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_254), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_254), .B1(n_260), .B2(n_232), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_319), .B(n_255), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_317), .B(n_267), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_342), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_345), .B(n_6), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_323), .B(n_254), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_323), .B(n_254), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_323), .B(n_267), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_362), .A2(n_239), .B(n_188), .C(n_8), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_260), .B(n_252), .C(n_238), .Y(n_384) );
OA211x2_ASAP7_75t_L g385 ( .A1(n_365), .A2(n_6), .B(n_7), .C(n_8), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_371), .B(n_7), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_361), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_188), .B(n_199), .C(n_207), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_356), .B(n_259), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_200), .B1(n_199), .B2(n_207), .C1(n_234), .C2(n_241), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_365), .B(n_259), .Y(n_392) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_369), .A2(n_244), .B1(n_222), .B2(n_10), .C(n_13), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_355), .A2(n_200), .B1(n_199), .B2(n_207), .C(n_146), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_367), .Y(n_395) );
NAND4xp75_ASAP7_75t_L g396 ( .A(n_359), .B(n_229), .C(n_259), .D(n_209), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_355), .A2(n_199), .B1(n_146), .B2(n_244), .C(n_16), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g398 ( .A1(n_378), .A2(n_229), .B(n_222), .C(n_202), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_348), .A2(n_229), .B(n_222), .C(n_259), .Y(n_399) );
AOI311xp33_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_9), .A3(n_16), .B(n_17), .C(n_18), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_352), .A2(n_259), .B1(n_191), .B2(n_195), .Y(n_401) );
NOR2xp33_ASAP7_75t_R g402 ( .A(n_349), .B(n_27), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_376), .A2(n_202), .B(n_259), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_379), .B(n_259), .Y(n_404) );
NAND4xp25_ASAP7_75t_SL g405 ( .A(n_372), .B(n_234), .C(n_252), .D(n_255), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_215), .B(n_209), .C(n_194), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_382), .A2(n_209), .B1(n_194), .B2(n_190), .C(n_97), .Y(n_408) );
AOI221xp5_ASAP7_75t_SL g409 ( .A1(n_374), .A2(n_97), .B1(n_194), .B2(n_30), .C(n_32), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_373), .A2(n_215), .B1(n_252), .B2(n_209), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_374), .A2(n_255), .B(n_265), .C(n_205), .Y(n_411) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_379), .B(n_215), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_363), .B(n_255), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_370), .B(n_28), .C(n_29), .D(n_33), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_350), .A2(n_215), .B1(n_39), .B2(n_40), .C(n_42), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g416 ( .A1(n_377), .A2(n_36), .B(n_43), .C(n_45), .Y(n_416) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_360), .A3(n_380), .B1(n_381), .B2(n_358), .C1(n_368), .C2(n_351), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_388), .B(n_375), .Y(n_418) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_405), .B(n_375), .Y(n_419) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_416), .B(n_353), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_400), .A2(n_265), .B(n_190), .C(n_201), .Y(n_421) );
NAND2xp33_ASAP7_75t_SL g422 ( .A(n_402), .B(n_46), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_407), .B(n_56), .Y(n_423) );
OR3x1_ASAP7_75t_L g424 ( .A(n_414), .B(n_58), .C(n_59), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_387), .B(n_60), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_413), .B(n_206), .Y(n_426) );
OAI321xp33_ASAP7_75t_L g427 ( .A1(n_393), .A2(n_62), .A3(n_63), .B1(n_64), .B2(n_65), .C(n_192), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_390), .B(n_404), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_394), .B(n_397), .C(n_392), .Y(n_429) );
AOI222xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_384), .B1(n_401), .B2(n_399), .C1(n_415), .C2(n_408), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_389), .B(n_416), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_409), .B(n_398), .C(n_406), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_411), .A2(n_391), .B1(n_410), .B2(n_403), .C(n_385), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_395), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_404), .B(n_390), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_388), .A2(n_369), .B1(n_328), .B2(n_393), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_437), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_435), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_428), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_422), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_424), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_418), .B(n_436), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_431), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_417), .B(n_433), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_436), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_426), .B(n_432), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_425), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_420), .A2(n_421), .B(n_429), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_423), .Y(n_450) );
CKINVDCx6p67_ASAP7_75t_R g451 ( .A(n_427), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_438), .A2(n_419), .B1(n_434), .B2(n_421), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_445), .B(n_430), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_440), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_447), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_449), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_452), .A2(n_439), .B1(n_443), .B2(n_444), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_455), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_456), .A2(n_439), .B1(n_443), .B2(n_446), .Y(n_459) );
OAI22x1_ASAP7_75t_L g460 ( .A1(n_453), .A2(n_441), .B1(n_442), .B2(n_450), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_458), .Y(n_461) );
XOR2xp5_ASAP7_75t_L g462 ( .A(n_460), .B(n_448), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_461), .A2(n_457), .B1(n_459), .B2(n_451), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_463), .A2(n_462), .B(n_454), .Y(n_464) );
endmodule