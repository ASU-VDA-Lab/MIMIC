module fake_jpeg_23418_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_45),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_24),
.Y(n_64)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_49),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_25),
.B1(n_15),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_70),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_16),
.B1(n_23),
.B2(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_58),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_18),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_23),
.C(n_19),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_26),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_44),
.B(n_41),
.C(n_42),
.D(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_77),
.B1(n_80),
.B2(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_86),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_29),
.B(n_26),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_24),
.B(n_41),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_94),
.B1(n_63),
.B2(n_67),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_3),
.B(n_4),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_92),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_68),
.B1(n_5),
.B2(n_10),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_68),
.B1(n_51),
.B2(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_60),
.B1(n_48),
.B2(n_12),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_79),
.B(n_77),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_122),
.B(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_103),
.B1(n_97),
.B2(n_95),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_105),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_83),
.B(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_74),
.C(n_78),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.C(n_99),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_133),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_98),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_80),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_106),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_147),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_121),
.A3(n_115),
.B1(n_114),
.B2(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_131),
.C(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_151),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_134),
.C(n_122),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_115),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_146),
.B(n_145),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_158),
.B(n_91),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_148),
.B1(n_141),
.B2(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_104),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_141),
.B(n_138),
.Y(n_158)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_157),
.B(n_89),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_104),
.C(n_154),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_161),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_87),
.Y(n_165)
);


endmodule