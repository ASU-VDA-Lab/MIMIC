module fake_jpeg_23348_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_14),
.B1(n_17),
.B2(n_13),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_39),
.C(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_15),
.B1(n_23),
.B2(n_24),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_30),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_7),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_71),
.C(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_31),
.B1(n_26),
.B2(n_41),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_67),
.B1(n_12),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_26),
.B1(n_37),
.B2(n_25),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_27),
.C(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_11),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_54),
.B(n_49),
.C(n_58),
.D(n_60),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_81),
.C(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_49),
.B(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_56),
.B1(n_52),
.B2(n_47),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_12),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_5),
.C(n_6),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_65),
.C(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_89),
.C(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_64),
.B1(n_61),
.B2(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_67),
.C(n_66),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_83),
.C(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_63),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_2),
.B(n_7),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_88),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_93),
.B(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_88),
.B1(n_9),
.B2(n_11),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_101),
.Y(n_108)
);

OAI321xp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_106),
.A3(n_107),
.B1(n_105),
.B2(n_9),
.C(n_2),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_2),
.Y(n_110)
);


endmodule