module fake_jpeg_20103_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_0),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_73),
.B1(n_79),
.B2(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_106),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_67),
.B1(n_62),
.B2(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_54),
.B1(n_78),
.B2(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_92),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_69),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_70),
.B1(n_75),
.B2(n_61),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_118),
.B1(n_120),
.B2(n_126),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_54),
.B1(n_72),
.B2(n_60),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_124),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_68),
.C(n_58),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_33),
.C(n_46),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_68),
.B1(n_58),
.B2(n_56),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_56),
.B1(n_52),
.B2(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_2),
.B(n_3),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_63),
.A3(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_35),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_134),
.B(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_119),
.C(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_142),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_2),
.B(n_4),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_141),
.B(n_5),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_5),
.B(n_6),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_150),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_149),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_36),
.B(n_47),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_154),
.B1(n_147),
.B2(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_144),
.B(n_145),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_153),
.C(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_123),
.Y(n_160)
);

AOI21x1_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_140),
.B(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_23),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_43),
.CI(n_45),
.CON(n_166),
.SN(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_10),
.Y(n_167)
);


endmodule