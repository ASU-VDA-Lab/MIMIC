module fake_aes_6630_n_25 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
BUFx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_0), .B(n_1), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_2), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_1), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_3), .B(n_5), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_16), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
OAI21xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_15), .B(n_18), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_6), .B(n_7), .Y(n_23) );
AOI21xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_8), .B(n_9), .Y(n_24) );
AOI22xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_25) );
endmodule