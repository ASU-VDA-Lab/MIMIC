module real_jpeg_25170_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_216;
wire n_213;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_71),
.B1(n_84),
.B2(n_88),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_71),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_88),
.B(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_79),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_4),
.B(n_26),
.C(n_27),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_69),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_41),
.B1(n_194),
.B2(n_199),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_5),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_73),
.Y(n_177)
);

INVx8_ASAP7_75t_SL g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_83),
.B1(n_84),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_7),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_7),
.A2(n_66),
.B1(n_68),
.B2(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_96),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_49)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_58),
.B1(n_66),
.B2(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_142)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_115),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_54),
.B1(n_97),
.B2(n_98),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_22),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_24),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_24),
.B(n_92),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_25),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_31),
.A2(n_32),
.B1(n_64),
.B2(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_31),
.B(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_32),
.A2(n_65),
.A3(n_68),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_32),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_57),
.B(n_59),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_35),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_35),
.A2(n_147),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_35),
.A2(n_146),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_35),
.A2(n_145),
.B1(n_146),
.B2(n_167),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_41),
.A2(n_48),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_41),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_41),
.A2(n_185),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_42),
.A2(n_46),
.B1(n_52),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_42),
.B(n_49),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_42),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_53),
.Y(n_203)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_75),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_72),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_61),
.A2(n_70),
.B1(n_74),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_62),
.A2(n_69),
.B1(n_129),
.B2(n_138),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_81),
.B(n_91),
.C(n_110),
.Y(n_109)
);

HAxp5_ASAP7_75t_SL g138 ( 
.A(n_66),
.B(n_92),
.CON(n_138),
.SN(n_138)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_80),
.C(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_87),
.B2(n_94),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_79),
.B1(n_95),
.B2(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_86),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.C(n_121),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_116),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_119),
.B(n_121),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_127),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_213),
.B(n_217),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_161),
.B(n_212),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_148),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_135),
.B(n_148),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.C(n_144),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_143),
.B(n_144),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_156),
.C(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_207),
.B(n_211),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_181),
.B(n_206),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_164),
.B(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_168),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_190),
.B(n_205),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_189),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_197),
.B(n_204),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);


endmodule