module fake_jpeg_10604_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_19),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_25),
.B1(n_34),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_51),
.B1(n_57),
.B2(n_68),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_26),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_52),
.B(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_34),
.B1(n_18),
.B2(n_17),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_20),
.CON(n_52),
.SN(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_34),
.B1(n_25),
.B2(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_45),
.C(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_30),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_33),
.B1(n_22),
.B2(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_54),
.B1(n_42),
.B2(n_58),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_96),
.Y(n_124)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_89),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_36),
.B1(n_30),
.B2(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_14),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_67),
.C(n_27),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_36),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_47),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_71),
.B(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_47),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_41),
.B1(n_27),
.B2(n_43),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_32),
.B1(n_24),
.B2(n_27),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_56),
.B1(n_67),
.B2(n_32),
.Y(n_106)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_32),
.B1(n_24),
.B2(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_126),
.B1(n_127),
.B2(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_14),
.C(n_16),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_119),
.C(n_130),
.Y(n_153)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_121),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_43),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_102),
.Y(n_144)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_103),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_1),
.C(n_2),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_140),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_96),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_138),
.B(n_5),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_139),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_149),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_73),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_6),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_84),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_148),
.C(n_112),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_87),
.B1(n_72),
.B2(n_83),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_150),
.B1(n_117),
.B2(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_76),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_100),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_94),
.B1(n_2),
.B2(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_16),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_93),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_129),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_1),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_108),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.C(n_144),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_180),
.B(n_155),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_139),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_6),
.B(n_7),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_138),
.B(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_184),
.B(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.C(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_132),
.C(n_149),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_176),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_199),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_134),
.C(n_150),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_178),
.B1(n_166),
.B2(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_162),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_173),
.C(n_177),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_173),
.B(n_169),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_192),
.B1(n_193),
.B2(n_158),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_180),
.C(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_163),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_182),
.B(n_197),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_163),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_188),
.B1(n_136),
.B2(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

OAI322xp33_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_199),
.A3(n_181),
.B1(n_196),
.B2(n_195),
.C1(n_184),
.C2(n_187),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_165),
.B1(n_159),
.B2(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_225),
.B1(n_203),
.B2(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_191),
.B1(n_203),
.B2(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_230),
.Y(n_235)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_171),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_171),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_223),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_228),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_216),
.B1(n_214),
.B2(n_223),
.C(n_218),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_240),
.B(n_7),
.Y(n_245)
);

OAI221xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_216),
.B1(n_218),
.B2(n_174),
.C(n_10),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_226),
.C(n_233),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_244),
.C(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_12),
.C(n_15),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.C(n_8),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_245),
.B(n_8),
.C(n_9),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_250),
.B(n_7),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_9),
.Y(n_253)
);


endmodule