module fake_jpeg_582_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_0),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_48),
.B1(n_42),
.B2(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_72),
.B1(n_56),
.B2(n_60),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_40),
.B1(n_49),
.B2(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_46),
.B1(n_38),
.B2(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_49),
.B1(n_46),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_61),
.B1(n_39),
.B2(n_41),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_79),
.B1(n_61),
.B2(n_69),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_85),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_44),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_69),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_45),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_65),
.B1(n_67),
.B2(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_67),
.B1(n_71),
.B2(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_95),
.B1(n_84),
.B2(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_51),
.B1(n_47),
.B2(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_51),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_100),
.C(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_19),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_82),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_113),
.B(n_18),
.Y(n_125)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_31),
.B(n_30),
.C(n_28),
.D(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_25),
.B(n_23),
.C(n_21),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_3),
.B(n_4),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_120),
.B(n_11),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_134),
.Y(n_142)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_109),
.C(n_111),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_113),
.C(n_15),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_117),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_14),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_135),
.B1(n_132),
.B2(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_131),
.B1(n_135),
.B2(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_148),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_136),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_149),
.A3(n_140),
.B1(n_139),
.B2(n_145),
.C1(n_148),
.C2(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_138),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_122),
.B(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_15),
.C(n_16),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_16),
.B(n_17),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_17),
.Y(n_156)
);


endmodule