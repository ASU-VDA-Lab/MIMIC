module fake_jpeg_19892_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_73),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_84),
.Y(n_87)
);

INVx2_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_52),
.B1(n_41),
.B2(n_57),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_86),
.B1(n_82),
.B2(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_41),
.B1(n_57),
.B2(n_55),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_50),
.B(n_66),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_45),
.B(n_65),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_98),
.B1(n_46),
.B2(n_58),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_62),
.B(n_44),
.C(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_59),
.B1(n_54),
.B2(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_40),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_109),
.B(n_1),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_49),
.B1(n_56),
.B2(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_0),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_120),
.B1(n_101),
.B2(n_106),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_126),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_132),
.B(n_124),
.C(n_121),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_116),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_131),
.C(n_127),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_117),
.C(n_135),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_130),
.B(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_14),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_15),
.C(n_18),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_19),
.Y(n_147)
);


endmodule