module real_aes_12127_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_698, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_698;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_92;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g158 ( .A(n_0), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g511 ( .A(n_1), .Y(n_511) );
AND2x2_ASAP7_75t_L g515 ( .A(n_1), .B(n_510), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_1), .B(n_61), .Y(n_526) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_1), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_2), .Y(n_164) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_3), .A2(n_62), .B1(n_496), .B2(n_501), .C(n_506), .Y(n_495) );
INVx1_ASAP7_75t_L g562 ( .A(n_3), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_4), .B(n_157), .Y(n_156) );
OR2x2_ASAP7_75t_L g573 ( .A(n_5), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g605 ( .A(n_5), .Y(n_605) );
BUFx2_ASAP7_75t_L g559 ( .A(n_6), .Y(n_559) );
INVx1_ASAP7_75t_L g575 ( .A(n_6), .Y(n_575) );
BUFx2_ASAP7_75t_L g600 ( .A(n_6), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_7), .B(n_165), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_8), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_9), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_10), .B(n_139), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_11), .A2(n_15), .B1(n_538), .B2(n_539), .C(n_540), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_11), .A2(n_15), .B1(n_647), .B2(n_651), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_12), .B(n_155), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_13), .B(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_13), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_14), .B(n_155), .Y(n_226) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_16), .Y(n_465) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g460 ( .A(n_18), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_19), .B(n_165), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_20), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_21), .B(n_124), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_22), .A2(n_44), .B1(n_519), .B2(n_527), .Y(n_518) );
INVx1_ASAP7_75t_L g628 ( .A(n_22), .Y(n_628) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_24), .B(n_139), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_25), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g574 ( .A(n_26), .Y(n_574) );
INVx1_ASAP7_75t_L g640 ( .A(n_26), .Y(n_640) );
NAND2xp33_ASAP7_75t_SL g122 ( .A(n_27), .B(n_90), .Y(n_122) );
INVx2_ASAP7_75t_SL g476 ( .A(n_28), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_29), .B(n_202), .Y(n_227) );
INVx1_ASAP7_75t_L g531 ( .A(n_30), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_30), .A2(n_31), .B1(n_656), .B2(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g535 ( .A(n_31), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_32), .A2(n_68), .B1(n_483), .B2(n_490), .Y(n_482) );
INVx1_ASAP7_75t_L g583 ( .A(n_32), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_33), .B(n_118), .Y(n_245) );
OAI21x1_ASAP7_75t_L g112 ( .A1(n_34), .A2(n_54), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_35), .B(n_202), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_36), .Y(n_471) );
INVx1_ASAP7_75t_L g517 ( .A(n_37), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_37), .A2(n_74), .B1(n_647), .B2(n_654), .Y(n_653) );
AND2x6_ASAP7_75t_L g84 ( .A(n_38), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_38), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_38), .B(n_666), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_39), .B(n_109), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_40), .B(n_109), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_41), .B(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_42), .A2(n_478), .B1(n_681), .B2(n_682), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_42), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_L g629 ( .A(n_44), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_45), .Y(n_151) );
INVx1_ASAP7_75t_L g85 ( .A(n_46), .Y(n_85) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_46), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_47), .B(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_48), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g119 ( .A(n_49), .B(n_90), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_124), .Y(n_199) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_50), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_51), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_52), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g489 ( .A(n_53), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_55), .B(n_139), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_56), .A2(n_59), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_56), .A2(n_59), .B1(n_642), .B2(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_57), .B(n_183), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_58), .B(n_202), .Y(n_247) );
BUFx10_ASAP7_75t_L g675 ( .A(n_60), .Y(n_675) );
INVx2_ASAP7_75t_L g510 ( .A(n_61), .Y(n_510) );
INVx1_ASAP7_75t_L g589 ( .A(n_62), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_63), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_64), .B(n_221), .Y(n_220) );
INVxp33_ASAP7_75t_SL g474 ( .A(n_64), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_65), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_66), .B(n_155), .Y(n_195) );
INVx2_ASAP7_75t_L g113 ( .A(n_67), .Y(n_113) );
INVx1_ASAP7_75t_L g576 ( .A(n_68), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_69), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_70), .B(n_137), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_71), .B(n_165), .Y(n_173) );
INVx2_ASAP7_75t_L g486 ( .A(n_72), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_73), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g549 ( .A(n_74), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_75), .Y(n_224) );
BUFx3_ASAP7_75t_L g568 ( .A(n_76), .Y(n_568) );
INVx1_ASAP7_75t_L g588 ( .A(n_76), .Y(n_588) );
BUFx3_ASAP7_75t_L g570 ( .A(n_77), .Y(n_570) );
INVx1_ASAP7_75t_L g581 ( .A(n_77), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_95), .B(n_453), .Y(n_78) );
BUFx2_ASAP7_75t_SL g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx2_ASAP7_75t_SL g127 ( .A(n_83), .Y(n_127) );
INVx8_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_84), .A2(n_126), .B(n_150), .C(n_153), .Y(n_149) );
OAI21x1_ASAP7_75t_SL g162 ( .A1(n_84), .A2(n_163), .B(n_170), .Y(n_162) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_84), .A2(n_194), .B(n_197), .Y(n_193) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g694 ( .A1(n_87), .A2(n_695), .B(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g172 ( .A(n_90), .Y(n_172) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_91), .Y(n_155) );
INVx1_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_93), .Y(n_92) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_93), .A2(n_154), .B(n_156), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_93), .A2(n_171), .B(n_173), .Y(n_170) );
BUFx12f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx5_ASAP7_75t_L g120 ( .A(n_94), .Y(n_120) );
INVx5_ASAP7_75t_L g169 ( .A(n_94), .Y(n_169) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NAND2x1p5_ASAP7_75t_L g98 ( .A(n_99), .B(n_374), .Y(n_98) );
NOR2x1_ASAP7_75t_L g99 ( .A(n_100), .B(n_298), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_101), .B(n_268), .Y(n_100) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_176), .B1(n_204), .B2(n_235), .C(n_248), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_129), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g327 ( .A(n_105), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_105), .B(n_326), .Y(n_392) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g276 ( .A(n_106), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g349 ( .A(n_106), .B(n_215), .Y(n_349) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g251 ( .A(n_107), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_107), .B(n_215), .Y(n_313) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_107), .Y(n_354) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g236 ( .A(n_108), .B(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_108), .Y(n_321) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_128), .Y(n_108) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_109), .A2(n_193), .B(n_201), .Y(n_192) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g175 ( .A(n_110), .Y(n_175) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx5_ASAP7_75t_L g133 ( .A(n_111), .Y(n_133) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g160 ( .A(n_112), .Y(n_160) );
OAI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B(n_127), .Y(n_114) );
O2A1O1Ixp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_119), .C(n_120), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g150 ( .A1(n_118), .A2(n_139), .B1(n_151), .B2(n_152), .Y(n_150) );
INVx2_ASAP7_75t_SL g126 ( .A(n_120), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_120), .A2(n_136), .B(n_138), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_120), .A2(n_182), .B(n_184), .Y(n_181) );
INVx2_ASAP7_75t_SL g200 ( .A(n_120), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B(n_126), .Y(n_121) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g137 ( .A(n_125), .Y(n_137) );
INVx2_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx2_ASAP7_75t_L g221 ( .A(n_125), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_126), .A2(n_141), .B(n_143), .Y(n_140) );
AOI21x1_ASAP7_75t_L g185 ( .A1(n_126), .A2(n_186), .B(n_187), .Y(n_185) );
OAI21x1_ASAP7_75t_L g180 ( .A1(n_127), .A2(n_181), .B(n_185), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_127), .A2(n_219), .B(n_223), .Y(n_218) );
INVx1_ASAP7_75t_SL g451 ( .A(n_129), .Y(n_451) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_147), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_130), .B(n_296), .Y(n_330) );
BUFx2_ASAP7_75t_L g352 ( .A(n_130), .Y(n_352) );
AND2x2_ASAP7_75t_L g367 ( .A(n_130), .B(n_210), .Y(n_367) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx3_ASAP7_75t_L g261 ( .A(n_131), .Y(n_261) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_145), .Y(n_132) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_133), .A2(n_149), .B(n_158), .Y(n_148) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_133), .A2(n_218), .B(n_227), .Y(n_217) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_133), .A2(n_240), .B(n_247), .Y(n_239) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_140), .B(n_144), .Y(n_134) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_144), .A2(n_241), .B(n_244), .Y(n_240) );
AND2x2_ASAP7_75t_L g372 ( .A(n_147), .B(n_178), .Y(n_372) );
AND2x2_ASAP7_75t_L g448 ( .A(n_147), .B(n_274), .Y(n_448) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_161), .Y(n_147) );
INVx3_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx2_ASAP7_75t_L g272 ( .A(n_148), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_148), .B(n_233), .Y(n_287) );
INVx5_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_159), .A2(n_162), .B(n_174), .Y(n_161) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
INVx3_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_167), .C(n_169), .Y(n_163) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g168 ( .A(n_166), .Y(n_168) );
INVx2_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_169), .A2(n_195), .B(n_196), .Y(n_194) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_169), .A2(n_224), .B(n_225), .C(n_226), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_169), .A2(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x6_ASAP7_75t_L g406 ( .A(n_177), .B(n_407), .Y(n_406) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_177), .A2(n_272), .A3(n_276), .B1(n_450), .B2(n_451), .B3(n_452), .Y(n_449) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_178), .B(n_343), .Y(n_396) );
INVx1_ASAP7_75t_L g419 ( .A(n_178), .Y(n_419) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
AND2x2_ASAP7_75t_L g206 ( .A(n_179), .B(n_192), .Y(n_206) );
BUFx2_ASAP7_75t_L g342 ( .A(n_179), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_189), .B(n_190), .Y(n_179) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_189), .B(n_190), .Y(n_234) );
AND2x2_ASAP7_75t_L g229 ( .A(n_191), .B(n_209), .Y(n_229) );
INVx1_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_191), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g323 ( .A(n_191), .B(n_264), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_191), .Y(n_340) );
INVx1_ASAP7_75t_L g369 ( .A(n_191), .Y(n_369) );
AND2x2_ASAP7_75t_L g380 ( .A(n_191), .B(n_333), .Y(n_380) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_200), .A2(n_220), .B(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_242), .B(n_243), .Y(n_241) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B1(n_216), .B2(n_228), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_206), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g303 ( .A(n_206), .Y(n_303) );
AND2x2_ASAP7_75t_L g331 ( .A(n_206), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_206), .B(n_290), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_206), .B(n_305), .Y(n_394) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_208), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_209), .Y(n_290) );
AND2x2_ASAP7_75t_L g305 ( .A(n_209), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_SL g333 ( .A(n_209), .Y(n_333) );
INVx1_ASAP7_75t_L g343 ( .A(n_209), .Y(n_343) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_209), .Y(n_385) );
AND2x2_ASAP7_75t_L g232 ( .A(n_210), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g306 ( .A(n_210), .Y(n_306) );
AND2x2_ASAP7_75t_L g332 ( .A(n_210), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x4_ASAP7_75t_L g316 ( .A(n_212), .B(n_297), .Y(n_316) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g422 ( .A(n_213), .B(n_250), .Y(n_422) );
INVx1_ASAP7_75t_L g435 ( .A(n_213), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
INVx2_ASAP7_75t_L g359 ( .A(n_214), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_214), .B(n_251), .Y(n_404) );
BUFx2_ASAP7_75t_L g429 ( .A(n_214), .Y(n_429) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g326 ( .A(n_216), .Y(n_326) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AND2x4_ASAP7_75t_L g273 ( .A(n_229), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g280 ( .A(n_229), .Y(n_280) );
AND2x2_ASAP7_75t_L g421 ( .A(n_229), .B(n_386), .Y(n_421) );
AND2x2_ASAP7_75t_L g443 ( .A(n_229), .B(n_271), .Y(n_443) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x6_ASAP7_75t_L g425 ( .A(n_231), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g322 ( .A(n_232), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g416 ( .A(n_232), .B(n_380), .Y(n_416) );
AND2x4_ASAP7_75t_L g266 ( .A(n_233), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g274 ( .A(n_233), .Y(n_274) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_R g386 ( .A(n_234), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_235), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g446 ( .A(n_235), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_236), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_236), .B(n_294), .Y(n_363) );
AOI322xp5_ASAP7_75t_L g364 ( .A1(n_236), .A2(n_318), .A3(n_365), .B1(n_368), .B2(n_370), .C1(n_372), .C2(n_373), .Y(n_364) );
INVx1_ASAP7_75t_L g277 ( .A(n_237), .Y(n_277) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g256 ( .A(n_238), .Y(n_256) );
AND2x2_ASAP7_75t_L g283 ( .A(n_238), .B(n_254), .Y(n_283) );
INVx1_ASAP7_75t_L g320 ( .A(n_238), .Y(n_320) );
AND2x2_ASAP7_75t_L g337 ( .A(n_238), .B(n_255), .Y(n_337) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI21xp33_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_257), .B(n_262), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_249), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
OR2x2_ASAP7_75t_L g329 ( .A(n_250), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g415 ( .A(n_250), .B(n_337), .Y(n_415) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g302 ( .A(n_251), .B(n_277), .Y(n_302) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g258 ( .A(n_253), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g408 ( .A(n_253), .B(n_352), .Y(n_408) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_254), .Y(n_311) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g296 ( .A(n_255), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_256), .Y(n_297) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g281 ( .A(n_260), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g301 ( .A(n_260), .B(n_302), .Y(n_301) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_260), .B(n_336), .Y(n_335) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_260), .B(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g294 ( .A(n_261), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g373 ( .A(n_261), .B(n_326), .Y(n_373) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
OR2x2_ASAP7_75t_L g399 ( .A(n_263), .B(n_285), .Y(n_399) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g450 ( .A(n_266), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B(n_278), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g279 ( .A(n_271), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g418 ( .A(n_271), .B(n_419), .Y(n_418) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_272), .B(n_340), .Y(n_371) );
INVx2_ASAP7_75t_L g362 ( .A(n_274), .Y(n_362) );
BUFx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g401 ( .A(n_276), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_276), .B(n_429), .Y(n_428) );
NAND2xp67_ASAP7_75t_SL g452 ( .A(n_276), .B(n_359), .Y(n_452) );
OAI222xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B1(n_281), .B2(n_284), .C1(n_291), .C2(n_293), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_281), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g393 ( .A(n_282), .Y(n_393) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g353 ( .A(n_283), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
BUFx3_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
NAND2x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g379 ( .A(n_287), .B(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2x1_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_294), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g439 ( .A(n_294), .B(n_388), .Y(n_439) );
INVx1_ASAP7_75t_L g445 ( .A(n_294), .Y(n_445) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_324), .C(n_344), .Y(n_298) );
AOI322xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .A3(n_304), .B1(n_307), .B2(n_309), .C1(n_314), .C2(n_322), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_301), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g388 ( .A(n_302), .Y(n_388) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
BUFx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g414 ( .A(n_305), .B(n_366), .Y(n_414) );
AND2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_308), .A2(n_425), .B1(n_428), .B2(n_430), .Y(n_427) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_316), .A2(n_377), .B1(n_379), .B2(n_381), .C1(n_383), .C2(n_387), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_318), .B(n_359), .Y(n_382) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g358 ( .A(n_319), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_322), .A2(n_325), .B1(n_328), .B2(n_331), .C(n_334), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g413 ( .A(n_327), .B(n_337), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_330), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g447 ( .A(n_330), .Y(n_447) );
INVx2_ASAP7_75t_L g407 ( .A(n_332), .Y(n_407) );
AND2x2_ASAP7_75t_L g432 ( .A(n_332), .B(n_386), .Y(n_432) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g348 ( .A(n_337), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g440 ( .A(n_337), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_339), .Y(n_345) );
AND2x4_ASAP7_75t_L g383 ( .A(n_339), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g366 ( .A(n_342), .Y(n_366) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_342), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B(n_355), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B1(n_360), .B2(n_363), .C(n_364), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_359), .A2(n_424), .B(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_385), .Y(n_426) );
INVx1_ASAP7_75t_L g378 ( .A(n_372), .Y(n_378) );
INVxp67_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_375), .B(n_411), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_389), .C(n_397), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_388), .B(n_435), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B(n_394), .C(n_395), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_396), .B(n_410), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_405), .B2(n_408), .C(n_409), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .C(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g411 ( .A(n_412), .B(n_423), .C(n_431), .D(n_442), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_436), .B2(n_439), .C1(n_440), .C2(n_698), .Y(n_431) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_446), .B2(n_448), .C(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI221xp5_ASAP7_75t_R g453 ( .A1(n_454), .A2(n_663), .B1(n_680), .B2(n_683), .C(n_687), .Y(n_453) );
XOR2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_478), .Y(n_454) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_469), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_462), .B1(n_467), .B2(n_468), .Y(n_456) );
INVx1_ASAP7_75t_L g467 ( .A(n_457), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_460), .Y(n_461) );
INVx1_ASAP7_75t_L g468 ( .A(n_462), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_465), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_473) );
INVx1_ASAP7_75t_SL g477 ( .A(n_474), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g682 ( .A(n_478), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_478), .A2(n_682), .B1(n_691), .B2(n_692), .Y(n_690) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR4xp75_ASAP7_75t_L g479 ( .A(n_480), .B(n_560), .C(n_596), .D(n_611), .Y(n_479) );
AOI31xp33_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_529), .A3(n_536), .B(n_556), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_495), .B1(n_512), .B2(n_517), .C(n_518), .Y(n_481) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g530 ( .A(n_484), .B(n_515), .Y(n_530) );
BUFx2_ASAP7_75t_L g544 ( .A(n_484), .Y(n_544) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g528 ( .A(n_485), .Y(n_528) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g493 ( .A(n_486), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g500 ( .A(n_486), .B(n_489), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_486), .Y(n_505) );
INVx1_ASAP7_75t_L g555 ( .A(n_486), .Y(n_555) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g494 ( .A(n_489), .Y(n_494) );
INVx1_ASAP7_75t_L g522 ( .A(n_489), .Y(n_522) );
INVx1_ASAP7_75t_L g554 ( .A(n_489), .Y(n_554) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AND2x4_ASAP7_75t_L g504 ( .A(n_494), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g610 ( .A(n_499), .Y(n_610) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_500), .Y(n_548) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g516 ( .A(n_504), .Y(n_516) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g542 ( .A(n_510), .Y(n_542) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
AND2x4_ASAP7_75t_L g532 ( .A(n_513), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g547 ( .A(n_515), .B(n_548), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OR2x6_ASAP7_75t_L g527 ( .A(n_524), .B(n_528), .Y(n_527) );
OR2x6_ASAP7_75t_L g551 ( .A(n_524), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_535), .Y(n_529) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_543), .B1(n_547), .B2(n_549), .C(n_550), .Y(n_536) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
CKINVDCx8_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g607 ( .A(n_558), .Y(n_607) );
OR2x6_ASAP7_75t_L g637 ( .A(n_558), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_582), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_576), .B2(n_577), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g601 ( .A(n_566), .B(n_602), .Y(n_601) );
INVx6_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g634 ( .A(n_567), .Y(n_634) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g580 ( .A(n_568), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g617 ( .A(n_568), .B(n_570), .Y(n_617) );
INVx1_ASAP7_75t_L g626 ( .A(n_569), .Y(n_626) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g587 ( .A(n_570), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g577 ( .A(n_571), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x6_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
OR2x6_ASAP7_75t_L g591 ( .A(n_572), .B(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_580), .Y(n_643) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_580), .Y(n_657) );
INVx1_ASAP7_75t_L g595 ( .A(n_581), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_589), .B2(n_590), .Y(n_582) );
CKINVDCx6p67_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
INVx1_ASAP7_75t_L g659 ( .A(n_587), .Y(n_659) );
INVx1_ASAP7_75t_L g594 ( .A(n_588), .Y(n_594) );
CKINVDCx6p67_ASAP7_75t_R g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_599), .B(n_606), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x4_ASAP7_75t_L g661 ( .A(n_600), .B(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_602), .B(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g678 ( .A(n_602), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x4_ASAP7_75t_L g662 ( .A(n_604), .B(n_640), .Y(n_662) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g639 ( .A(n_605), .B(n_640), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_621), .C(n_635), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_615), .Y(n_654) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g652 ( .A(n_616), .Y(n_652) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g627 ( .A(n_619), .Y(n_627) );
OR2x6_ASAP7_75t_L g631 ( .A(n_619), .B(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g673 ( .A(n_624), .Y(n_673) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g679 ( .A(n_625), .Y(n_679) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI33xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_641), .A3(n_646), .B1(n_653), .B2(n_655), .B3(n_660), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_SL g671 ( .A(n_639), .Y(n_671) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx4f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x6_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
OR2x4_ASAP7_75t_L g689 ( .A(n_665), .B(n_669), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_666), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g695 ( .A(n_666), .Y(n_695) );
INVx1_ASAP7_75t_L g686 ( .A(n_667), .Y(n_686) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI31xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .A3(n_674), .B(n_676), .Y(n_669) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx6_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_691), .B2(n_693), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_691), .Y(n_692) );
BUFx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
endmodule