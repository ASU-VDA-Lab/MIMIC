module fake_jpeg_27544_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_42),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_45),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_26),
.B1(n_16),
.B2(n_18),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_26),
.B1(n_16),
.B2(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_60),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_16),
.B1(n_26),
.B2(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_42),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_28),
.B(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_38),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_34),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_80),
.B1(n_63),
.B2(n_43),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_65),
.B1(n_86),
.B2(n_82),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_40),
.B1(n_39),
.B2(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_41),
.B1(n_21),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_22),
.B(n_32),
.C(n_29),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_114),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_20),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_51),
.B(n_37),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_48),
.C(n_29),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_27),
.C(n_17),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_94),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_138)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_32),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_104),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_88),
.B1(n_66),
.B2(n_41),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_102),
.B1(n_65),
.B2(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_41),
.B1(n_59),
.B2(n_61),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_38),
.Y(n_141)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_110),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_51),
.B1(n_28),
.B2(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_75),
.B1(n_87),
.B2(n_81),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_142),
.B(n_116),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_65),
.B1(n_70),
.B2(n_89),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_89),
.B1(n_74),
.B2(n_21),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_128),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_140),
.B1(n_97),
.B2(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_115),
.B1(n_98),
.B2(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_89),
.B1(n_74),
.B2(n_21),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_132),
.B1(n_90),
.B2(n_38),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_74),
.B1(n_38),
.B2(n_37),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_37),
.B(n_38),
.C(n_20),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_110),
.B(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.C(n_96),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_27),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_38),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_149),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_99),
.B(n_104),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_146),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_155),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_152),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_158),
.A2(n_163),
.B1(n_168),
.B2(n_31),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_25),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_166),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_90),
.B(n_108),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_165),
.B(n_169),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_20),
.B(n_17),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_20),
.B(n_17),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_20),
.B(n_27),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_1),
.Y(n_197)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_137),
.B1(n_124),
.B2(n_133),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_135),
.B1(n_133),
.B2(n_136),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_184),
.B1(n_188),
.B2(n_192),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_133),
.B(n_19),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_169),
.B(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_27),
.C(n_19),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_179),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_27),
.C(n_19),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_18),
.C(n_25),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_182),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_25),
.B1(n_31),
.B2(n_8),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

NAND4xp25_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_31),
.C(n_2),
.D(n_3),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_8),
.A3(n_14),
.B1(n_12),
.B2(n_10),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_200),
.B1(n_156),
.B2(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_157),
.B(n_146),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_219),
.B1(n_225),
.B2(n_186),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_210),
.B1(n_222),
.B2(n_191),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_148),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_149),
.B1(n_160),
.B2(n_171),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_145),
.B1(n_165),
.B2(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_4),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_5),
.Y(n_224)
);

OAI21x1_ASAP7_75t_SL g228 ( 
.A1(n_224),
.A2(n_222),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_208),
.B(n_174),
.CI(n_181),
.CON(n_226),
.SN(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_182),
.C(n_178),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_209),
.C(n_220),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_179),
.C(n_187),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_207),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_184),
.B1(n_199),
.B2(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_176),
.B1(n_180),
.B2(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_210),
.B1(n_203),
.B2(n_214),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_176),
.B(n_180),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_215),
.B1(n_224),
.B2(n_211),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_202),
.B(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_204),
.B(n_9),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_259),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_230),
.B1(n_240),
.B2(n_234),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_232),
.C(n_226),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_216),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_254),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_213),
.C(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_261),
.Y(n_274)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g262 ( 
.A(n_255),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_7),
.C(n_8),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_236),
.B1(n_231),
.B2(n_233),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_260),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_275),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_256),
.B(n_255),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_237),
.B(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_234),
.B1(n_226),
.B2(n_244),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_286),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_258),
.C(n_248),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_205),
.C(n_238),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_9),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_6),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_265),
.B(n_262),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_263),
.B(n_274),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_293),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_267),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_15),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_12),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_14),
.B(n_15),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_5),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_276),
.Y(n_298)
);

OAI21x1_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_303),
.B(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_280),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_276),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_299),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_296),
.B(n_303),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.C(n_288),
.Y(n_311)
);

NAND2x1_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_305),
.Y(n_312)
);


endmodule