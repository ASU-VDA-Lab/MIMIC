module fake_netlist_1_11657_n_623 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_623, n_193);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_623;
output n_193;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_69), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_61), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_70), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_22), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_57), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_73), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_56), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_32), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_36), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_27), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_14), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_62), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_53), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_39), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_51), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_1), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_13), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_30), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_18), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_45), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_50), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_58), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_66), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_10), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_7), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_9), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_41), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_68), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_115), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_78), .Y(n_121) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_79), .A2(n_23), .B(n_71), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_114), .Y(n_123) );
NAND2x1_ASAP7_75t_L g124 ( .A(n_81), .B(n_0), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_111), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_102), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_80), .A2(n_72), .B(n_67), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_86), .B(n_2), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_86), .B(n_2), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_105), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_105), .B(n_3), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_102), .Y(n_134) );
NAND2x1_ASAP7_75t_L g135 ( .A(n_81), .B(n_3), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_100), .B(n_4), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_115), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_116), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_104), .B(n_5), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_88), .B(n_5), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_88), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_99), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_104), .B(n_6), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_117), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_107), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_87), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_90), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_90), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_91), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_127), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_131), .A2(n_89), .B1(n_103), .B2(n_77), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_127), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_132), .B(n_74), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_126), .B(n_119), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_131), .A2(n_118), .B1(n_112), .B2(n_91), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_132), .B(n_75), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_131), .B(n_89), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_134), .B(n_98), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_131), .B(n_133), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_127), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_144), .B(n_97), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_144), .B(n_101), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_136), .Y(n_178) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_122), .A2(n_118), .B(n_93), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
INVx4_ASAP7_75t_SL g181 ( .A(n_133), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
AO22x2_ASAP7_75t_L g183 ( .A1(n_133), .A2(n_93), .B1(n_112), .B2(n_94), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_147), .B(n_109), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_147), .B(n_106), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_136), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_133), .B(n_94), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_136), .B(n_92), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_141), .B(n_113), .Y(n_192) );
UNKNOWN g193 ( );
INVx1_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_139), .B(n_110), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_130), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_120), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_141), .B(n_108), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_122), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_128), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_148), .B(n_96), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_128), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_156), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_128), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_152), .B(n_95), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_138), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_156), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_156), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_200), .Y(n_217) );
BUFx12f_ASAP7_75t_L g218 ( .A(n_214), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_200), .Y(n_219) );
AND3x2_ASAP7_75t_SL g220 ( .A(n_167), .B(n_157), .C(n_122), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_203), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_211), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_181), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_181), .B(n_129), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_199), .B(n_129), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_199), .B(n_159), .Y(n_227) );
BUFx4f_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_191), .B(n_149), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_176), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_211), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_201), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
AND3x1_ASAP7_75t_SL g235 ( .A(n_193), .B(n_125), .C(n_158), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_191), .B(n_159), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_214), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_202), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_197), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_167), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_181), .B(n_149), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_167), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_178), .B(n_158), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_178), .B(n_140), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_188), .B(n_189), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_188), .B(n_140), .Y(n_248) );
AOI22x1_ASAP7_75t_L g249 ( .A1(n_212), .A2(n_157), .B1(n_155), .B2(n_153), .Y(n_249) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_161), .A2(n_146), .B(n_155), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_189), .B(n_153), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_205), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_181), .B(n_124), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
NOR3xp33_ASAP7_75t_SL g255 ( .A(n_165), .B(n_121), .C(n_123), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_189), .B(n_142), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_175), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_189), .B(n_142), .Y(n_259) );
INVx5_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_210), .Y(n_261) );
NAND3xp33_ASAP7_75t_SL g262 ( .A(n_173), .B(n_135), .C(n_124), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_171), .B(n_150), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_175), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_162), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_167), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_172), .B(n_146), .C(n_143), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_171), .B(n_135), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_171), .B(n_150), .Y(n_272) );
BUFx8_ASAP7_75t_L g273 ( .A(n_171), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_185), .B(n_143), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_216), .Y(n_275) );
NOR3xp33_ASAP7_75t_SL g276 ( .A(n_208), .B(n_76), .C(n_8), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_232), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_224), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_222), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_229), .B(n_185), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
BUFx4_ASAP7_75t_SL g282 ( .A(n_240), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_273), .A2(n_183), .B1(n_173), .B2(n_213), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_183), .B1(n_190), .B2(n_204), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_229), .B(n_187), .Y(n_285) );
INVx5_ASAP7_75t_L g286 ( .A(n_224), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_218), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_241), .A2(n_183), .B1(n_204), .B2(n_192), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_266), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_243), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_273), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_228), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_227), .A2(n_206), .B(n_176), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_221), .Y(n_295) );
NAND2x1_ASAP7_75t_L g296 ( .A(n_243), .B(n_176), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_226), .A2(n_206), .B(n_192), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_218), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_250), .A2(n_261), .B(n_259), .C(n_256), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_274), .B(n_187), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_271), .B(n_183), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_264), .B(n_195), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_271), .B(n_195), .Y(n_303) );
INVx3_ASAP7_75t_SL g304 ( .A(n_240), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_251), .A2(n_206), .B(n_192), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_263), .A2(n_204), .B(n_192), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_222), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_261), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_273), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_231), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_233), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_233), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_234), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_244), .Y(n_318) );
INVx8_ASAP7_75t_L g319 ( .A(n_242), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_271), .B(n_169), .Y(n_320) );
NAND3x1_ASAP7_75t_L g321 ( .A(n_245), .B(n_177), .C(n_164), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_237), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_244), .A2(n_204), .B1(n_212), .B2(n_215), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_322), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_303), .B(n_257), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_282), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_319), .B(n_269), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_318), .A2(n_269), .B1(n_228), .B2(n_225), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_322), .B(n_236), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_295), .B(n_228), .Y(n_331) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_299), .A2(n_179), .B(n_220), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_303), .B(n_225), .Y(n_333) );
INVx8_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
AOI221x1_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_212), .B1(n_162), .B2(n_209), .C(n_207), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_303), .B(n_246), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_318), .A2(n_225), .B1(n_242), .B2(n_262), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_288), .A2(n_284), .B1(n_283), .B2(n_321), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_285), .A2(n_248), .B1(n_255), .B2(n_270), .C(n_276), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_321), .A2(n_272), .B1(n_238), .B2(n_268), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_302), .B(n_242), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_301), .A2(n_253), .B1(n_267), .B2(n_234), .Y(n_343) );
BUFx10_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_302), .B(n_217), .Y(n_345) );
INVx6_ASAP7_75t_L g346 ( .A(n_281), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_304), .A2(n_235), .B1(n_253), .B2(n_234), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_292), .B(n_253), .Y(n_349) );
INVx8_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_313), .B(n_219), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_339), .A2(n_304), .B1(n_291), .B2(n_320), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_327), .B(n_319), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_330), .A2(n_310), .B1(n_291), .B2(n_287), .Y(n_356) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_332), .A2(n_305), .B(n_179), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_346), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_325), .B(n_287), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_324), .A2(n_298), .B1(n_292), .B2(n_294), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_323), .B1(n_306), .B2(n_292), .C(n_309), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_341), .A2(n_277), .B1(n_294), .B2(n_309), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_327), .A2(n_277), .B1(n_311), .B2(n_315), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_298), .B1(n_267), .B2(n_317), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_352), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_311), .B1(n_315), .B2(n_316), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_317), .B1(n_230), .B2(n_260), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_345), .B(n_279), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_342), .A2(n_297), .B1(n_157), .B2(n_223), .C(n_239), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_333), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_337), .B(n_331), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_349), .B(n_281), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
BUFx5_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
AO21x1_ASAP7_75t_SL g379 ( .A1(n_354), .A2(n_347), .B(n_338), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_356), .A2(n_328), .B(n_343), .C(n_216), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
OAI31xp33_ASAP7_75t_L g382 ( .A1(n_365), .A2(n_349), .A3(n_329), .B(n_252), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_378), .Y(n_383) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_357), .A2(n_332), .B(n_179), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_367), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_369), .B(n_332), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_369), .B(n_327), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_372), .Y(n_388) );
OAI33xp33_ASAP7_75t_L g389 ( .A1(n_362), .A2(n_174), .A3(n_163), .B1(n_166), .B2(n_168), .B3(n_180), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_378), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_360), .A2(n_198), .B(n_258), .C(n_265), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_376), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
NAND5xp2_ASAP7_75t_SL g396 ( .A(n_364), .B(n_344), .C(n_8), .D(n_9), .E(n_11), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_363), .A2(n_349), .B(n_279), .C(n_312), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_374), .A2(n_373), .B1(n_375), .B2(n_361), .C(n_359), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_373), .B(n_308), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_375), .A2(n_249), .B1(n_316), .B2(n_312), .C(n_308), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_370), .B(n_344), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
BUFx10_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_355), .A2(n_350), .B1(n_334), .B2(n_317), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_198), .A3(n_254), .B(n_275), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_355), .A2(n_350), .B1(n_334), .B2(n_344), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_357), .B(n_335), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_355), .A2(n_350), .B1(n_334), .B2(n_346), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_368), .A2(n_163), .B(n_166), .C(n_168), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_378), .A2(n_350), .B1(n_334), .B2(n_346), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_403), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_386), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_386), .B(n_378), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_398), .A2(n_371), .B1(n_378), .B2(n_358), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_398), .A2(n_7), .A3(n_11), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_392), .B(n_358), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_395), .B(n_378), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g422 ( .A1(n_391), .A2(n_275), .A3(n_254), .B(n_220), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_403), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_385), .B(n_378), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_384), .B(n_377), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_401), .B(n_12), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_384), .B(n_377), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_391), .B(n_15), .C(n_16), .D(n_17), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_384), .B(n_377), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_384), .B(n_377), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_399), .B(n_17), .Y(n_434) );
AOI322xp5_ASAP7_75t_L g435 ( .A1(n_407), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_21), .C1(n_22), .C2(n_220), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_399), .B(n_19), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_394), .B(n_377), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_405), .B(n_21), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_394), .B(n_128), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_408), .B(n_212), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_408), .B(n_348), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_383), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_383), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_393), .B(n_348), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_383), .B(n_348), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g448 ( .A(n_409), .B(n_24), .C(n_25), .D(n_28), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_402), .B(n_209), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_390), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_387), .B(n_207), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_390), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_387), .B(n_207), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_382), .B(n_162), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_425), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_413), .B(n_382), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_425), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_420), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_413), .B(n_397), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_414), .B(n_406), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_416), .B(n_403), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_414), .B(n_379), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_427), .B(n_380), .Y(n_467) );
OR2x6_ASAP7_75t_L g468 ( .A(n_412), .B(n_406), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_421), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_417), .A2(n_404), .B(n_411), .C(n_396), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_418), .B(n_400), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_429), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_426), .B(n_379), .Y(n_474) );
NOR4xp25_ASAP7_75t_SL g475 ( .A(n_456), .B(n_400), .C(n_380), .D(n_410), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_424), .B(n_209), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_445), .B(n_29), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_434), .B(n_207), .Y(n_478) );
OAI33xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_410), .A3(n_182), .B1(n_180), .B2(n_194), .B3(n_186), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_419), .B(n_296), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_429), .Y(n_481) );
AOI22x1_ASAP7_75t_L g482 ( .A1(n_412), .A2(n_196), .B1(n_160), .B2(n_170), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g483 ( .A(n_423), .B(n_314), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_412), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_438), .B(n_389), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_435), .A2(n_182), .B(n_194), .C(n_186), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_443), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_430), .A2(n_174), .B(n_160), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_444), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_445), .B(n_34), .Y(n_496) );
NAND2xp33_ASAP7_75t_L g497 ( .A(n_423), .B(n_314), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_426), .B(n_196), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_446), .B(n_296), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_451), .B(n_162), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_428), .B(n_196), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_451), .B(n_162), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_446), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_441), .B(n_37), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_447), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_454), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_432), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_468), .A2(n_415), .B1(n_457), .B2(n_452), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_459), .Y(n_510) );
NAND2x1_ASAP7_75t_L g511 ( .A(n_485), .B(n_468), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_504), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_490), .B(n_433), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_461), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_469), .Y(n_515) );
AOI21xp33_ASAP7_75t_SL g516 ( .A1(n_468), .A2(n_422), .B(n_452), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_472), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_506), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_492), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_468), .A2(n_452), .B1(n_453), .B2(n_450), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_467), .A2(n_448), .B1(n_428), .B2(n_455), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_467), .A2(n_455), .B1(n_450), .B2(n_437), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g523 ( .A1(n_489), .A2(n_442), .B(n_449), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_506), .B(n_437), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_489), .B(n_447), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_470), .B(n_449), .C(n_439), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_493), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_460), .A2(n_207), .B1(n_162), .B2(n_209), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_495), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_491), .A2(n_170), .B(n_160), .C(n_290), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_474), .A2(n_209), .B(n_207), .Y(n_531) );
AOI211xp5_ASAP7_75t_L g532 ( .A1(n_466), .A2(n_483), .B(n_497), .C(n_471), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_466), .B(n_38), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_508), .B(n_209), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_500), .Y(n_535) );
OAI21xp5_ASAP7_75t_SL g536 ( .A1(n_477), .A2(n_290), .B(n_278), .Y(n_536) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_483), .Y(n_537) );
OAI32xp33_ASAP7_75t_L g538 ( .A1(n_505), .A2(n_278), .A3(n_290), .B1(n_44), .B2(n_46), .Y(n_538) );
OAI322xp33_ASAP7_75t_L g539 ( .A1(n_463), .A2(n_249), .A3(n_278), .B1(n_266), .B2(n_52), .C1(n_54), .C2(n_63), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_494), .A2(n_42), .B(n_43), .C(n_47), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_508), .B(n_65), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_480), .A2(n_281), .B1(n_307), .B2(n_286), .C1(n_230), .C2(n_260), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_498), .B(n_184), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_481), .B(n_184), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_465), .B(n_184), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_479), .A2(n_266), .B1(n_230), .B2(n_260), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_486), .B(n_184), .Y(n_547) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_497), .B(n_314), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_487), .B(n_184), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_499), .B(n_184), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_507), .B(n_230), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_539), .B(n_478), .C(n_502), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_513), .B(n_484), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_536), .A2(n_477), .B(n_496), .Y(n_554) );
NAND2xp33_ASAP7_75t_SL g555 ( .A(n_511), .B(n_477), .Y(n_555) );
INVx3_ASAP7_75t_SL g556 ( .A(n_518), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_532), .B(n_496), .Y(n_557) );
AND2x4_ASAP7_75t_SL g558 ( .A(n_524), .B(n_496), .Y(n_558) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_525), .A2(n_498), .B1(n_502), .B2(n_473), .C1(n_488), .C2(n_484), .Y(n_559) );
XNOR2xp5_ASAP7_75t_L g560 ( .A(n_512), .B(n_464), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_514), .Y(n_562) );
NOR3xp33_ASAP7_75t_SL g563 ( .A(n_509), .B(n_476), .C(n_501), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_537), .A2(n_482), .B(n_462), .Y(n_566) );
NAND2x1_ASAP7_75t_L g567 ( .A(n_548), .B(n_462), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_519), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_527), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_523), .A2(n_458), .B1(n_503), .B2(n_475), .C(n_230), .Y(n_570) );
NOR3xp33_ASAP7_75t_SL g571 ( .A(n_520), .B(n_286), .C(n_307), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_543), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_535), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_523), .B(n_260), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_526), .Y(n_576) );
OAI211xp5_ASAP7_75t_L g577 ( .A1(n_516), .A2(n_286), .B(n_307), .C(n_260), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_533), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_576), .A2(n_521), .B(n_540), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_562), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_562), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_564), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_563), .B(n_522), .C(n_550), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_555), .A2(n_542), .A3(n_531), .B(n_545), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_556), .A2(n_541), .B1(n_549), .B2(n_547), .Y(n_586) );
XOR2x2_ASAP7_75t_L g587 ( .A(n_556), .B(n_549), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_554), .B(n_547), .Y(n_588) );
XNOR2x2_ASAP7_75t_SL g589 ( .A(n_560), .B(n_528), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_563), .A2(n_544), .B(n_538), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_559), .B(n_534), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_567), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_579), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_578), .B(n_568), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_561), .Y(n_595) );
NOR2x1p5_ASAP7_75t_L g596 ( .A(n_557), .B(n_551), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_566), .B(n_530), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_570), .A2(n_546), .B(n_289), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_589), .A2(n_558), .B(n_577), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_580), .A2(n_571), .B(n_552), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_585), .A2(n_571), .B(n_573), .C(n_552), .Y(n_601) );
NOR2xp33_ASAP7_75t_R g602 ( .A(n_593), .B(n_575), .Y(n_602) );
BUFx12f_ASAP7_75t_L g603 ( .A(n_596), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_584), .A2(n_574), .B1(n_572), .B2(n_569), .Y(n_604) );
INVxp33_ASAP7_75t_L g605 ( .A(n_587), .Y(n_605) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_597), .B(n_565), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_591), .B(n_553), .Y(n_607) );
OAI322xp33_ASAP7_75t_L g608 ( .A1(n_588), .A2(n_594), .A3(n_582), .B1(n_595), .B2(n_581), .C1(n_592), .C2(n_583), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_598), .A2(n_581), .B(n_586), .C(n_583), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_585), .A2(n_576), .B1(n_589), .B2(n_590), .C(n_584), .Y(n_610) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_580), .A2(n_585), .B(n_576), .C(n_584), .Y(n_611) );
OA22x2_ASAP7_75t_L g612 ( .A1(n_611), .A2(n_600), .B1(n_610), .B2(n_607), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_603), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_599), .B(n_601), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_602), .Y(n_615) );
NOR3xp33_ASAP7_75t_SL g616 ( .A(n_613), .B(n_608), .C(n_609), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_614), .B(n_604), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_615), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_618), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_617), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_619), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_621), .A2(n_612), .B1(n_614), .B2(n_620), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_622), .A2(n_616), .B(n_605), .C(n_606), .Y(n_623) );
endmodule