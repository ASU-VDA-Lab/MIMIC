module fake_netlist_1_2797_n_826 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_191, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_826);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_826;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_132), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_40), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_120), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_17), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_177), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_1), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_167), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_63), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_188), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_192), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_66), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_195), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_151), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_92), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_164), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_24), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_112), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_178), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_157), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_11), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_84), .B(n_124), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_62), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_182), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_180), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_133), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_146), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_115), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_51), .B(n_15), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_107), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_27), .Y(n_234) );
NOR2xp67_ASAP7_75t_L g235 ( .A(n_125), .B(n_24), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_2), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_29), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_88), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_97), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_136), .Y(n_240) );
INVxp33_ASAP7_75t_SL g241 ( .A(n_109), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_121), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_35), .Y(n_243) );
CKINVDCx14_ASAP7_75t_R g244 ( .A(n_18), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_134), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_174), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_48), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_93), .Y(n_248) );
BUFx2_ASAP7_75t_SL g249 ( .A(n_172), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_75), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_29), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_82), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_131), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_19), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_49), .Y(n_255) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_26), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_80), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_40), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_98), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_42), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_83), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_90), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_30), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_50), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_34), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_5), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_61), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_169), .B(n_59), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_95), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_49), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_18), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_12), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_73), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_41), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_162), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_173), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_61), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_60), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_38), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_189), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_161), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_103), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_39), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_47), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_56), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_171), .Y(n_287) );
CKINVDCx14_ASAP7_75t_R g288 ( .A(n_21), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_152), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_187), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_22), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_78), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_2), .Y(n_293) );
INVx2_ASAP7_75t_SL g294 ( .A(n_156), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_1), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_13), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_119), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_79), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_110), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_105), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_135), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_160), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_81), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_13), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_106), .Y(n_305) );
INVxp33_ASAP7_75t_SL g306 ( .A(n_154), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_223), .B(n_0), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_245), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_212), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_223), .B(n_0), .Y(n_311) );
BUFx8_ASAP7_75t_L g312 ( .A(n_225), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_245), .Y(n_313) );
INVx5_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_212), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_251), .B(n_3), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_205), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_258), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_222), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_205), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_222), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_244), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_323) );
OAI22xp5_ASAP7_75t_SL g324 ( .A1(n_219), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_200), .B(n_7), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_236), .B(n_8), .Y(n_326) );
OAI22x1_ASAP7_75t_SL g327 ( .A1(n_219), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_258), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_264), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_264), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_198), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_199), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_244), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_333) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_269), .B(n_197), .Y(n_334) );
BUFx8_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_287), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_14), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_288), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_334), .B(n_215), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_335), .B(n_220), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_334), .A2(n_288), .B1(n_252), .B2(n_221), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_331), .B(n_297), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_326), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_326), .Y(n_346) );
AND3x4_ASAP7_75t_L g347 ( .A(n_326), .B(n_235), .C(n_227), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_326), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_307), .B(n_285), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_332), .B(n_282), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_333), .B(n_291), .C(n_259), .Y(n_353) );
AND2x6_ASAP7_75t_L g354 ( .A(n_307), .B(n_218), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_308), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_307), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_307), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_338), .B(n_206), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_311), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_332), .B(n_287), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_334), .A2(n_252), .B1(n_221), .B2(n_284), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_311), .A2(n_203), .B1(n_243), .B2(n_234), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_311), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_311), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_320), .B(n_298), .Y(n_370) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_325), .B(n_202), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_314), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_316), .B(n_284), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_319), .B(n_208), .C(n_207), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_310), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_314), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_321), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_321), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_344), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_359), .B(n_312), .Y(n_383) );
NOR2xp33_ASAP7_75t_SL g384 ( .A(n_369), .B(n_312), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_346), .A2(n_337), .B1(n_322), .B2(n_329), .Y(n_385) );
INVx5_ASAP7_75t_L g386 ( .A(n_354), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_346), .A2(n_337), .B1(n_322), .B2(n_329), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_378), .Y(n_390) );
NOR2x2_ASAP7_75t_L g391 ( .A(n_364), .B(n_327), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_350), .B(n_250), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_348), .A2(n_317), .B(n_330), .C(n_232), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_350), .B(n_250), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_374), .B(n_276), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_374), .B(n_286), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_349), .B(n_281), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_342), .B(n_241), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_369), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_371), .B(n_306), .Y(n_403) );
AND2x6_ASAP7_75t_SL g404 ( .A(n_370), .B(n_327), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_368), .B(n_283), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_351), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_351), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_362), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_368), .B(n_290), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_357), .A2(n_330), .B(n_317), .C(n_323), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_354), .B(n_290), .Y(n_412) );
OR2x6_ASAP7_75t_L g413 ( .A(n_362), .B(n_324), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_352), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_364), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_366), .B(n_292), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_354), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_347), .B(n_320), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_354), .B(n_292), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_366), .B(n_302), .Y(n_420) );
O2A1O1Ixp5_ASAP7_75t_L g421 ( .A1(n_357), .A2(n_270), .B(n_217), .C(n_209), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_354), .B(n_302), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_354), .B(n_320), .Y(n_423) );
INVx8_ASAP7_75t_L g424 ( .A(n_354), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_341), .B(n_204), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_348), .B(n_228), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_345), .B(n_339), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_341), .A2(n_278), .B1(n_296), .B2(n_267), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_345), .B(n_231), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_357), .B(n_238), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_361), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_367), .B(n_242), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_358), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_343), .B(n_286), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_367), .B(n_248), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_367), .B(n_253), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_361), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_358), .B(n_303), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_365), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_358), .B(n_256), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_363), .B(n_263), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_343), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_365), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_380), .B(n_274), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_375), .A2(n_211), .B(n_210), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_380), .B(n_300), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_353), .B(n_247), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_347), .A2(n_226), .B1(n_237), .B2(n_201), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_433), .A2(n_347), .B(n_372), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_417), .B(n_296), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_381), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_433), .A2(n_377), .B(n_372), .Y(n_452) );
BUFx8_ASAP7_75t_SL g453 ( .A(n_413), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_421), .A2(n_379), .B(n_378), .C(n_255), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_382), .B(n_379), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_381), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_392), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_429), .A2(n_377), .B(n_379), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_440), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_387), .B(n_379), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_261), .B1(n_265), .B2(n_254), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_387), .B(n_397), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
AND2x2_ASAP7_75t_SL g465 ( .A(n_417), .B(n_266), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_421), .A2(n_272), .B(n_273), .C(n_271), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_399), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_418), .A2(n_279), .B1(n_280), .B2(n_275), .Y(n_469) );
NAND2xp33_ASAP7_75t_L g470 ( .A(n_424), .B(n_258), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_424), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_411), .A2(n_295), .B(n_304), .C(n_293), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_445), .A2(n_214), .B(n_213), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_434), .A2(n_447), .B1(n_383), .B2(n_420), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_401), .B(n_249), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g478 ( .A1(n_425), .A2(n_216), .B(n_229), .C(n_224), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_440), .B(n_268), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_426), .A2(n_233), .B(n_230), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_393), .B(n_239), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_427), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_386), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_423), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_410), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_407), .Y(n_487) );
OR2x6_ASAP7_75t_L g488 ( .A(n_447), .B(n_240), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_441), .B(n_246), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_406), .A2(n_400), .B(n_444), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_405), .Y(n_492) );
BUFx8_ASAP7_75t_L g493 ( .A(n_391), .Y(n_493) );
BUFx12f_ASAP7_75t_L g494 ( .A(n_404), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_395), .A2(n_260), .B(n_262), .C(n_257), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_408), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_386), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_409), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_394), .B(n_396), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_414), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_409), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_432), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_385), .B(n_299), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_439), .A2(n_305), .B(n_301), .C(n_218), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_443), .B(n_20), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_409), .B(n_227), .Y(n_507) );
INVx6_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_389), .A2(n_277), .B1(n_289), .B2(n_314), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_435), .B(n_277), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_390), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_430), .A2(n_289), .B(n_310), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_412), .Y(n_513) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_419), .B(n_289), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_438), .B(n_22), .Y(n_515) );
NAND3xp33_ASAP7_75t_SL g516 ( .A(n_446), .B(n_355), .C(n_340), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_422), .B(n_23), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_436), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_428), .B(n_356), .C(n_355), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_437), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_421), .A2(n_336), .B(n_313), .C(n_318), .Y(n_521) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_424), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_384), .B(n_314), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_398), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_382), .B(n_23), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_383), .B(n_25), .Y(n_526) );
AO32x2_ASAP7_75t_L g527 ( .A1(n_448), .A2(n_310), .A3(n_313), .B1(n_318), .B2(n_328), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_421), .A2(n_336), .B(n_313), .C(n_318), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_384), .B(n_310), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_382), .B(n_25), .Y(n_530) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_424), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_437), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_382), .A2(n_313), .B1(n_318), .B2(n_328), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_382), .A2(n_313), .B1(n_318), .B2(n_328), .Y(n_534) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_450), .A2(n_27), .B1(n_28), .B2(n_30), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_451), .A2(n_336), .B1(n_328), .B2(n_373), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_499), .A2(n_360), .B(n_356), .Y(n_537) );
AO31x2_ASAP7_75t_L g538 ( .A1(n_521), .A2(n_376), .A3(n_373), .B(n_360), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_520), .B(n_28), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_455), .A2(n_356), .B(n_336), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_495), .A2(n_31), .B(n_32), .C(n_33), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_490), .A2(n_336), .B(n_328), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_476), .B(n_463), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_457), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_520), .B(n_34), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_488), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_459), .A2(n_65), .B(n_64), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_506), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_525), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_488), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_465), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_528), .A2(n_68), .B(n_67), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_530), .Y(n_554) );
CKINVDCx14_ASAP7_75t_R g555 ( .A(n_494), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_456), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_516), .A2(n_70), .B(n_69), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_479), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_486), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_453), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_466), .A2(n_113), .B(n_194), .C(n_193), .Y(n_561) );
BUFx10_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_452), .A2(n_72), .B(n_71), .Y(n_564) );
O2A1O1Ixp5_ASAP7_75t_L g565 ( .A1(n_529), .A2(n_523), .B(n_515), .C(n_477), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_508), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_460), .B(n_52), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_489), .A2(n_117), .B(n_191), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_480), .A2(n_55), .B(n_57), .C(n_58), .Y(n_569) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_512), .A2(n_118), .B(n_190), .Y(n_570) );
AO32x2_ASAP7_75t_L g571 ( .A1(n_509), .A2(n_57), .A3(n_58), .B1(n_59), .B2(n_60), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_462), .B(n_62), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_508), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_487), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_496), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_449), .A2(n_123), .B(n_74), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_SL g577 ( .A1(n_505), .A2(n_126), .B(n_76), .C(n_77), .Y(n_577) );
BUFx8_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_482), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_522), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_SL g581 ( .A1(n_517), .A2(n_89), .B(n_91), .C(n_94), .Y(n_581) );
BUFx10_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
BUFx3_ASAP7_75t_L g583 ( .A(n_474), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_500), .B(n_96), .Y(n_584) );
AOI21xp5_ASAP7_75t_SL g585 ( .A1(n_482), .A2(n_99), .B(n_100), .Y(n_585) );
NOR2x1_ASAP7_75t_SL g586 ( .A(n_464), .B(n_101), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_504), .B(n_102), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_461), .B(n_491), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_502), .B(n_104), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_454), .B(n_108), .Y(n_590) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_475), .A2(n_111), .B(n_114), .Y(n_591) );
AO31x2_ASAP7_75t_L g592 ( .A1(n_533), .A2(n_116), .A3(n_122), .B(n_127), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_478), .A2(n_128), .B(n_129), .C(n_130), .Y(n_593) );
INVx5_ASAP7_75t_L g594 ( .A(n_474), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_518), .Y(n_595) );
AOI21x1_ASAP7_75t_L g596 ( .A1(n_507), .A2(n_137), .B(n_138), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_469), .A2(n_140), .B1(n_141), .B2(n_143), .Y(n_597) );
AND2x6_ASAP7_75t_L g598 ( .A(n_464), .B(n_144), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_458), .Y(n_599) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_467), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_464), .Y(n_601) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_510), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_481), .A2(n_145), .B(n_147), .Y(n_603) );
BUFx3_ASAP7_75t_L g604 ( .A(n_518), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_503), .A2(n_149), .B(n_150), .Y(n_605) );
CKINVDCx11_ASAP7_75t_R g606 ( .A(n_471), .Y(n_606) );
INVx6_ASAP7_75t_L g607 ( .A(n_484), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_532), .B(n_155), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_513), .A2(n_158), .B1(n_159), .B2(n_163), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_471), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_485), .A2(n_165), .B(n_166), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_471), .Y(n_612) );
CKINVDCx12_ASAP7_75t_R g613 ( .A(n_531), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_514), .A2(n_175), .B1(n_179), .B2(n_181), .Y(n_614) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_484), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_519), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_468), .B(n_196), .Y(n_617) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_534), .A2(n_184), .A3(n_185), .B(n_186), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_472), .B(n_497), .Y(n_619) );
AO31x2_ASAP7_75t_L g620 ( .A1(n_492), .A2(n_501), .A3(n_498), .B(n_527), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_470), .A2(n_472), .B(n_511), .C(n_484), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_594), .B(n_497), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_543), .B(n_475), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_574), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_602), .B(n_511), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_548), .B(n_575), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_599), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_567), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_551), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_544), .B(n_546), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_539), .Y(n_632) );
AO21x2_ASAP7_75t_L g633 ( .A1(n_540), .A2(n_553), .B(n_576), .Y(n_633) );
INVx6_ASAP7_75t_L g634 ( .A(n_578), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_541), .A2(n_550), .B1(n_559), .B2(n_535), .C(n_588), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_558), .A2(n_565), .B(n_569), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_594), .B(n_583), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_600), .B(n_582), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_545), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_590), .A2(n_584), .B(n_587), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_556), .Y(n_641) );
NOR2x1_ASAP7_75t_R g642 ( .A(n_560), .B(n_606), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_589), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_566), .A2(n_598), .B1(n_597), .B2(n_562), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_608), .A2(n_621), .B1(n_617), .B2(n_609), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_562), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_571), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_561), .A2(n_581), .B(n_547), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_617), .A2(n_610), .B1(n_595), .B2(n_604), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_571), .Y(n_650) );
OAI21x1_ASAP7_75t_SL g651 ( .A1(n_611), .A2(n_586), .B(n_605), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_613), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_557), .A2(n_577), .B(n_564), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_568), .A2(n_603), .B(n_593), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_612), .B(n_601), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_555), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_573), .B(n_619), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_580), .A2(n_607), .B1(n_601), .B2(n_536), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_615), .B(n_579), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_563), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_620), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_563), .B(n_579), .Y(n_662) );
NOR2x1_ASAP7_75t_R g663 ( .A(n_563), .B(n_579), .Y(n_663) );
INVxp33_ASAP7_75t_L g664 ( .A(n_585), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_596), .A2(n_538), .B(n_620), .Y(n_665) );
CKINVDCx12_ASAP7_75t_R g666 ( .A(n_614), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_538), .B(n_591), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_618), .B(n_592), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_570), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_592), .B(n_618), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_618), .B(n_415), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_575), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_574), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_552), .A2(n_364), .B1(n_343), .B2(n_465), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_574), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_575), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_543), .B(n_382), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_543), .B(n_382), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_575), .Y(n_679) );
CKINVDCx12_ASAP7_75t_R g680 ( .A(n_555), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_549), .A2(n_526), .B(n_554), .C(n_473), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_575), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_542), .A2(n_616), .B(n_537), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_575), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_542), .A2(n_616), .B(n_537), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_575), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_543), .B(n_382), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_575), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_616), .A2(n_455), .B(n_521), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_574), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_574), .Y(n_691) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
OAI21x1_ASAP7_75t_SL g693 ( .A1(n_611), .A2(n_586), .B(n_605), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_552), .B(n_450), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_552), .B(n_398), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_542), .A2(n_616), .B(n_537), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_575), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_552), .B(n_398), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_594), .B(n_483), .Y(n_699) );
INVx3_ASAP7_75t_L g700 ( .A(n_594), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_546), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_552), .A2(n_364), .B1(n_343), .B2(n_465), .Y(n_702) );
OR2x6_ASAP7_75t_L g703 ( .A(n_649), .B(n_692), .Y(n_703) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_663), .Y(n_704) );
OR2x6_ASAP7_75t_L g705 ( .A(n_692), .B(n_645), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_624), .B(n_627), .Y(n_706) );
AO21x2_ASAP7_75t_L g707 ( .A1(n_668), .A2(n_670), .B(n_667), .Y(n_707) );
INVx3_ASAP7_75t_L g708 ( .A(n_692), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_673), .B(n_675), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_662), .B(n_643), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_702), .A2(n_671), .B1(n_635), .B2(n_641), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_690), .B(n_691), .Y(n_712) );
BUFx2_ASAP7_75t_L g713 ( .A(n_663), .Y(n_713) );
OA21x2_ASAP7_75t_L g714 ( .A1(n_647), .A2(n_650), .B(n_685), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_626), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_629), .A2(n_698), .B1(n_695), .B2(n_694), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_672), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_676), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_628), .A2(n_681), .B1(n_682), .B2(n_697), .C(n_684), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_661), .Y(n_720) );
OR2x6_ASAP7_75t_L g721 ( .A(n_700), .B(n_632), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_679), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_631), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_646), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_686), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_688), .B(n_677), .Y(n_726) );
AO21x2_ASAP7_75t_L g727 ( .A1(n_683), .A2(n_696), .B(n_648), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_678), .B(n_687), .Y(n_728) );
INVxp67_ASAP7_75t_L g729 ( .A(n_701), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_665), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_689), .B(n_699), .Y(n_731) );
AO21x2_ASAP7_75t_L g732 ( .A1(n_623), .A2(n_693), .B(n_651), .Y(n_732) );
AO21x2_ASAP7_75t_L g733 ( .A1(n_636), .A2(n_689), .B(n_633), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_644), .B(n_639), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_625), .B(n_652), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_637), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_657), .Y(n_737) );
INVx3_ASAP7_75t_L g738 ( .A(n_622), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_659), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_655), .B(n_660), .Y(n_740) );
INVxp67_ASAP7_75t_L g741 ( .A(n_638), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_634), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_658), .B(n_664), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_654), .B(n_640), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_630), .B(n_653), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_642), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_666), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_656), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_663), .Y(n_749) );
CKINVDCx6p67_ASAP7_75t_R g750 ( .A(n_680), .Y(n_750) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_668), .A2(n_670), .B(n_669), .Y(n_751) );
BUFx3_ASAP7_75t_L g752 ( .A(n_692), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_674), .A2(n_552), .B1(n_450), .B2(n_702), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_647), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_626), .Y(n_755) );
OR2x6_ASAP7_75t_L g756 ( .A(n_649), .B(n_539), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_731), .B(n_754), .Y(n_757) );
BUFx3_ASAP7_75t_L g758 ( .A(n_736), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_731), .B(n_722), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_715), .B(n_755), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_725), .B(n_706), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_709), .B(n_712), .Y(n_762) );
INVx5_ASAP7_75t_SL g763 ( .A(n_750), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_753), .A2(n_747), .B1(n_734), .B2(n_711), .Y(n_764) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_728), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_726), .B(n_717), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_720), .Y(n_767) );
INVx4_ASAP7_75t_L g768 ( .A(n_703), .Y(n_768) );
AND2x4_ASAP7_75t_SL g769 ( .A(n_703), .B(n_756), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_733), .B(n_718), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_737), .B(n_723), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_730), .Y(n_772) );
INVx1_ASAP7_75t_SL g773 ( .A(n_724), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_719), .B(n_716), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_705), .B(n_743), .Y(n_775) );
OR2x6_ASAP7_75t_SL g776 ( .A(n_745), .B(n_747), .Y(n_776) );
BUFx3_ASAP7_75t_L g777 ( .A(n_736), .Y(n_777) );
AND2x4_ASAP7_75t_SL g778 ( .A(n_703), .B(n_756), .Y(n_778) );
AND2x2_ASAP7_75t_SL g779 ( .A(n_713), .B(n_749), .Y(n_779) );
OR2x6_ASAP7_75t_L g780 ( .A(n_705), .B(n_756), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_714), .B(n_744), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_781), .B(n_751), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_781), .B(n_751), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_757), .B(n_770), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_770), .B(n_707), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_773), .B(n_748), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_759), .B(n_707), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_759), .B(n_707), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_764), .A2(n_746), .B1(n_729), .B2(n_741), .C(n_721), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_779), .B(n_746), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_767), .B(n_732), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_767), .B(n_739), .Y(n_792) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_772), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_761), .B(n_740), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_771), .B(n_742), .Y(n_795) );
AND2x4_ASAP7_75t_L g796 ( .A(n_768), .B(n_727), .Y(n_796) );
NOR2x1_ASAP7_75t_L g797 ( .A(n_790), .B(n_780), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_796), .B(n_775), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_784), .B(n_765), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_794), .B(n_762), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_789), .B(n_776), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_796), .B(n_775), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_793), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_795), .B(n_776), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_786), .B(n_774), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_787), .B(n_766), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_787), .B(n_760), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_788), .B(n_775), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_808), .B(n_782), .Y(n_809) );
AO21x1_ASAP7_75t_L g810 ( .A1(n_801), .A2(n_778), .B(n_769), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_805), .B(n_804), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_798), .Y(n_812) );
AOI322xp5_ASAP7_75t_L g813 ( .A1(n_811), .A2(n_799), .A3(n_800), .B1(n_797), .B2(n_806), .C1(n_807), .C2(n_783), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_810), .A2(n_802), .B1(n_785), .B2(n_780), .Y(n_814) );
OAI21xp5_ASAP7_75t_SL g815 ( .A1(n_814), .A2(n_778), .B(n_812), .Y(n_815) );
OAI211xp5_ASAP7_75t_L g816 ( .A1(n_813), .A2(n_803), .B(n_768), .C(n_735), .Y(n_816) );
NAND3xp33_ASAP7_75t_SL g817 ( .A(n_816), .B(n_763), .C(n_768), .Y(n_817) );
AOI211xp5_ASAP7_75t_SL g818 ( .A1(n_817), .A2(n_815), .B(n_763), .C(n_704), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_818), .B(n_752), .C(n_708), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_819), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_820), .Y(n_821) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_821), .B(n_809), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_822), .A2(n_721), .B(n_792), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_823), .A2(n_708), .B(n_738), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_824), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_825), .A2(n_710), .B1(n_777), .B2(n_758), .C(n_791), .Y(n_826) );
endmodule