module fake_jpeg_17715_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_45),
.B1(n_60),
.B2(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_17),
.B1(n_22),
.B2(n_20),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_51),
.Y(n_83)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_57),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_19),
.B(n_30),
.C(n_25),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_65),
.B(n_64),
.C(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_0),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.C(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_32),
.A2(n_17),
.B1(n_22),
.B2(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_15),
.B1(n_17),
.B2(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_73),
.B1(n_61),
.B2(n_54),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_71),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_15),
.B1(n_60),
.B2(n_26),
.Y(n_99)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_15),
.B1(n_29),
.B2(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_61),
.B1(n_25),
.B2(n_30),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_53),
.B(n_57),
.C(n_49),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_95),
.B(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_92),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_61),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_45),
.B(n_43),
.C(n_63),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_79),
.B1(n_73),
.B2(n_72),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_42),
.B1(n_38),
.B2(n_51),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_108),
.B1(n_60),
.B2(n_48),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_92),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_63),
.C(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_52),
.B1(n_48),
.B2(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_99),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_124),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_52),
.B1(n_58),
.B2(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_117),
.B1(n_125),
.B2(n_127),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_72),
.B1(n_82),
.B2(n_78),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_123),
.B1(n_93),
.B2(n_97),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_121),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_84),
.B1(n_42),
.B2(n_71),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_83),
.B(n_77),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_71),
.B1(n_76),
.B2(n_59),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_73),
.B1(n_42),
.B2(n_38),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_105),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_51),
.B1(n_85),
.B2(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_94),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_18),
.C(n_28),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_125),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_28),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_29),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_112),
.B1(n_91),
.B2(n_97),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_106),
.B1(n_87),
.B2(n_104),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_120),
.B1(n_109),
.B2(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_91),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_126),
.C(n_117),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_161),
.C(n_174),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_126),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_141),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_118),
.B(n_123),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_193)
);

NOR2x1p5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_144),
.B1(n_137),
.B2(n_155),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_97),
.B1(n_85),
.B2(n_108),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_24),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_40),
.C(n_35),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_40),
.C(n_110),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_177),
.C(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_40),
.C(n_110),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_150),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_189),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_188),
.C(n_191),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_194),
.B(n_196),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_165),
.B1(n_19),
.B2(n_21),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_151),
.C(n_143),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_154),
.C(n_147),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_168),
.A3(n_171),
.B1(n_176),
.B2(n_163),
.C(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_18),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_24),
.C(n_31),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_197),
.C(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_31),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_30),
.C(n_26),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_174),
.C(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_8),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_209),
.C(n_213),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_212),
.B1(n_214),
.B2(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_167),
.C(n_172),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_180),
.B(n_165),
.CI(n_28),
.CON(n_210),
.SN(n_210)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_19),
.C(n_21),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_8),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_192),
.B(n_188),
.C(n_195),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_203),
.B(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_198),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_215),
.B1(n_13),
.B2(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_9),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_224),
.C(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_21),
.C(n_18),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_0),
.C(n_1),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_211),
.B1(n_202),
.B2(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_1),
.C(n_2),
.Y(n_227)
);

AOI31xp33_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_9),
.A3(n_12),
.B(n_11),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_5),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_203),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_6),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_240),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_219),
.B1(n_206),
.B2(n_225),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_235),
.B(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_250),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_220),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_234),
.B(n_235),
.Y(n_248)
);

NOR4xp25_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_3),
.C(n_5),
.D(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_220),
.C(n_4),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_238),
.B1(n_239),
.B2(n_3),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_5),
.B(n_250),
.C(n_245),
.D(n_249),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_253),
.B(n_258),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_262),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_254),
.B(n_259),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

XOR2x2_ASAP7_75t_R g267 ( 
.A(n_264),
.B(n_260),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);


endmodule