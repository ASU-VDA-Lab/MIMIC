module fake_netlist_6_1514_n_3082 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_3082);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_3082;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_2534;
wire n_2353;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_2480;
wire n_641;
wire n_2739;
wire n_1300;
wire n_3023;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_659;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_2971;
wire n_1713;
wire n_1111;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_3069;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_437;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_627;
wire n_1767;
wire n_595;
wire n_1779;
wire n_1465;
wire n_524;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_925;
wire n_1101;
wire n_2535;
wire n_1880;
wire n_1026;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_2693;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3037;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2667;
wire n_2539;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1774;
wire n_884;
wire n_1398;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_474;
wire n_1207;
wire n_683;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_2263;
wire n_994;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_609;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_2716;
wire n_1320;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2699;
wire n_2272;
wire n_2200;
wire n_3029;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_3045;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_799;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1045;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_430;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_841;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_2969;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_2769;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_3035;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_2600;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_3038;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_2899;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_66),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_23),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_51),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_125),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_291),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_187),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_251),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_38),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_235),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_271),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_159),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_337),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_174),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_284),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_365),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_199),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_48),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_408),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_141),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_300),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_26),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_229),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_36),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_249),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_42),
.Y(n_435)
);

BUFx8_ASAP7_75t_SL g436 ( 
.A(n_306),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_208),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_224),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_206),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_221),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_357),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_401),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_347),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_20),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_46),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_108),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_157),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_329),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_164),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_98),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_399),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_74),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_5),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_90),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_48),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_161),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_362),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_166),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_218),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_183),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_380),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_55),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_205),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_178),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_43),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_215),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_54),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_57),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_333),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_409),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_100),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_241),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_179),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_349),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_231),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_159),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_54),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_278),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_171),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_187),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_237),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_146),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_301),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_207),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_211),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_18),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_64),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_28),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_384),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_308),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_256),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_7),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_272),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_213),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_236),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_9),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_379),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_268),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_263),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_279),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_175),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_71),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_172),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_270),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_109),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_43),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_74),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_351),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_316),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_167),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_222),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_376),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_318),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_78),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_285),
.Y(n_519)
);

BUFx8_ASAP7_75t_SL g520 ( 
.A(n_51),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_180),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_180),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_0),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_196),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_158),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_7),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_173),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_361),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_156),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_150),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_348),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_161),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_332),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_276),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_28),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_239),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_60),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_264),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_149),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_406),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_32),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_324),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_9),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_343),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_72),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_155),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_25),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_38),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_214),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_375),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_267),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_287),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_137),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_36),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_21),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_363),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_154),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_230),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_403),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_77),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_114),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_134),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_153),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_257),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_216),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_277),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_297),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_387),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_41),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_114),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_95),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_65),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_244),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_364),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_153),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_217),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_262),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_238),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_296),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_163),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_122),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_32),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_103),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_395),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_280),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_109),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_243),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_3),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_265),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_330),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_197),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_116),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_252),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_175),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_204),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_154),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_56),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_195),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_293),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_118),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_353),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_15),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_202),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_39),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g605 ( 
.A(n_100),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_254),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_189),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_157),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_325),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_149),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_194),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_92),
.Y(n_612)
);

BUFx5_ASAP7_75t_L g613 ( 
.A(n_17),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_292),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_253),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_111),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_121),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_34),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_25),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_336),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_120),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_396),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_352),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_400),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_127),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_372),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_255),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_212),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_170),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_405),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_190),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_385),
.Y(n_632)
);

INVxp33_ASAP7_75t_SL g633 ( 
.A(n_60),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_172),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_178),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_17),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_163),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_339),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_135),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_183),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_62),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_26),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_58),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_130),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_33),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_340),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_266),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_21),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_371),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_107),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_93),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_65),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_126),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_119),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_147),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_354),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_116),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_140),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_103),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_66),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_13),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_123),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_392),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_73),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_46),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_309),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_77),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_99),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_171),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_304),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_240),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_303),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_319),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_294),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_31),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_11),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_19),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_53),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_84),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_193),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_22),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_320),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_232),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_112),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_166),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_382),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_367),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_123),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_150),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_108),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_331),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_90),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_133),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_5),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_68),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_97),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_219),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_40),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_317),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_15),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_174),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_0),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_86),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_370),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_307),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_143),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_223),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_120),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_33),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_315),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_20),
.Y(n_711)
);

CKINVDCx6p67_ASAP7_75t_R g712 ( 
.A(n_137),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_220),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_104),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_179),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_346),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_545),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_613),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_520),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_417),
.Y(n_720)
);

CKINVDCx14_ASAP7_75t_R g721 ( 
.A(n_649),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_598),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_504),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_662),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_613),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_667),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_613),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_613),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_613),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_613),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_421),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_613),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_664),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_664),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_664),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_531),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_485),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_712),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_712),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_664),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_664),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_451),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_451),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_451),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_579),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_451),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_451),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_485),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_592),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_592),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_592),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_420),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_442),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_482),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_453),
.B(n_1),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_411),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_420),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_447),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_484),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_435),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_432),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_435),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_447),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_492),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_412),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_456),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_453),
.B(n_1),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_545),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_432),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_432),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_490),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_600),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_461),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_468),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_600),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_495),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_698),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_698),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_415),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_429),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_431),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_479),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_481),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_425),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_426),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_488),
.Y(n_792)
);

INVxp33_ASAP7_75t_L g793 ( 
.A(n_506),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_452),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_508),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_456),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_514),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_523),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_525),
.Y(n_799)
);

BUFx2_ASAP7_75t_SL g800 ( 
.A(n_502),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_532),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_535),
.Y(n_802)
);

XNOR2xp5_ASAP7_75t_L g803 ( 
.A(n_462),
.B(n_2),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_537),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_510),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_546),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_518),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_554),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_521),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_557),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_560),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_447),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_449),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_569),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_571),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_476),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_522),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_572),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_410),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_583),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_575),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_594),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_602),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_610),
.Y(n_824)
);

INVxp33_ASAP7_75t_SL g825 ( 
.A(n_410),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_612),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_631),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_634),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_640),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_477),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_478),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_526),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_478),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_575),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_499),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_575),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_499),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_529),
.Y(n_839)
);

INVxp33_ASAP7_75t_L g840 ( 
.A(n_655),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_529),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_528),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_548),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_548),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_553),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_553),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_452),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_413),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_639),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_487),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_639),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_678),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_678),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_657),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_452),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_658),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_748),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_770),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_741),
.B(n_502),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_794),
.B(n_491),
.Y(n_861)
);

CKINVDCx11_ASAP7_75t_R g862 ( 
.A(n_732),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_759),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_770),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_770),
.Y(n_865)
);

CKINVDCx11_ASAP7_75t_R g866 ( 
.A(n_779),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_748),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_780),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_746),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_748),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_746),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_747),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_752),
.B(n_615),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_747),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_750),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_774),
.B(n_643),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_750),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_751),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_751),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_753),
.Y(n_880)
);

CKINVDCx11_ASAP7_75t_R g881 ( 
.A(n_842),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_753),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_720),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_767),
.B(n_615),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_775),
.B(n_691),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_754),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_754),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_755),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_755),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_778),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_756),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_756),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_757),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_740),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_757),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_721),
.B(n_691),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_800),
.B(n_489),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_731),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_825),
.A2(n_633),
.B1(n_605),
.B2(n_624),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_800),
.B(n_434),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_735),
.A2(n_726),
.B(n_725),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_728),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_720),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_758),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_776),
.B(n_423),
.Y(n_906)
);

BUFx8_ASAP7_75t_SL g907 ( 
.A(n_719),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_718),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_790),
.B(n_423),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_791),
.B(n_439),
.Y(n_910)
);

OA21x2_ASAP7_75t_L g911 ( 
.A1(n_729),
.A2(n_497),
.B(n_439),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_813),
.B(n_497),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_785),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_816),
.B(n_501),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_786),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_723),
.A2(n_727),
.B1(n_722),
.B2(n_724),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_758),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_772),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_718),
.Y(n_920)
);

OAI22x1_ASAP7_75t_SL g921 ( 
.A1(n_722),
.A2(n_509),
.B1(n_543),
.B2(n_505),
.Y(n_921)
);

OAI22x1_ASAP7_75t_SL g922 ( 
.A1(n_724),
.A2(n_563),
.B1(n_596),
.B2(n_555),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_787),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_760),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_772),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_796),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_796),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_845),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_760),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_794),
.Y(n_930)
);

OAI22x1_ASAP7_75t_SL g931 ( 
.A1(n_719),
.A2(n_641),
.B1(n_651),
.B2(n_608),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_733),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_781),
.B(n_643),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_845),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_682),
.B(n_501),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_734),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_717),
.Y(n_937)
);

BUFx8_ASAP7_75t_SL g938 ( 
.A(n_742),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_734),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_736),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_736),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_831),
.B(n_682),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_825),
.A2(n_627),
.B1(n_623),
.B2(n_530),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_749),
.A2(n_539),
.B1(n_541),
.B2(n_527),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_742),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_769),
.A2(n_616),
.B1(n_422),
.B2(n_427),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_788),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_737),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_737),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_738),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_850),
.B(n_710),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_738),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_739),
.B(n_492),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_847),
.B(n_710),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_847),
.B(n_494),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_739),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_744),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_744),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_745),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_745),
.A2(n_517),
.B(n_513),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_763),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_764),
.B(n_821),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_854),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_765),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_854),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_855),
.B(n_533),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_783),
.B(n_542),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_789),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_792),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_765),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_795),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_777),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_763),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_766),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_784),
.B(n_773),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_797),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_766),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_768),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_798),
.B(n_544),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_R g980 ( 
.A(n_924),
.B(n_777),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_872),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_896),
.B(n_782),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_902),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_900),
.B(n_761),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_902),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_872),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_863),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_864),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_906),
.B(n_975),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_959),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_864),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_959),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_906),
.B(n_782),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_864),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_920),
.Y(n_995)
);

CKINVDCx16_ASAP7_75t_R g996 ( 
.A(n_868),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_920),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_932),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_937),
.B(n_835),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_906),
.B(n_805),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_979),
.B(n_573),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_937),
.B(n_805),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_937),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_932),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_864),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_878),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_878),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_879),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_937),
.Y(n_1009)
);

AND2x6_ASAP7_75t_L g1010 ( 
.A(n_975),
.B(n_492),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_865),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_879),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_949),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_886),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_949),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_865),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_892),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_950),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_892),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_865),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_950),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_SL g1023 ( 
.A1(n_899),
.A2(n_803),
.B1(n_422),
.B2(n_427),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_893),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_893),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_895),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_975),
.B(n_807),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_865),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_909),
.B(n_912),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_895),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_909),
.B(n_717),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_898),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_956),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_898),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_909),
.B(n_768),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_937),
.B(n_897),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_979),
.B(n_551),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_905),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_956),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_957),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_905),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_912),
.B(n_807),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_912),
.B(n_809),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_905),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_957),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_930),
.B(n_809),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_936),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_943),
.A2(n_803),
.B1(n_433),
.B2(n_444),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_905),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_898),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_915),
.B(n_817),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_898),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_915),
.B(n_832),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_958),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_958),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_908),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_908),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_898),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_926),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_926),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_904),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_901),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_908),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_939),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_926),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_904),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_901),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_862),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_930),
.B(n_817),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_972),
.B(n_833),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_939),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_939),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_940),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_940),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_901),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_940),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_903),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_915),
.B(n_832),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_903),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_914),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_867),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_914),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_869),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_926),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_926),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_928),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_928),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_888),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_890),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_935),
.A2(n_558),
.B(n_552),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_936),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_936),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_928),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_972),
.B(n_436),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_928),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_936),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_901),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_936),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_901),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_979),
.B(n_566),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_941),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_941),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_859),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_941),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_941),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_953),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_884),
.B(n_833),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_924),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_928),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_942),
.B(n_951),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_859),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_942),
.B(n_834),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_941),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_948),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_942),
.B(n_855),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_929),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_934),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_934),
.Y(n_1120)
);

OR2x2_ASAP7_75t_SL g1121 ( 
.A(n_964),
.B(n_819),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_948),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_945),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_885),
.B(n_743),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_934),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_967),
.B(n_578),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_948),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_951),
.B(n_556),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_967),
.B(n_867),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_951),
.B(n_834),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_944),
.A2(n_561),
.B1(n_562),
.B2(n_547),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_860),
.B(n_647),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_934),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_890),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_948),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_948),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_873),
.B(n_480),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_952),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_929),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_919),
.B(n_483),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_952),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_967),
.B(n_836),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_952),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_952),
.Y(n_1144)
);

XNOR2xp5_ASAP7_75t_L g1145 ( 
.A(n_921),
.B(n_922),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_952),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_970),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_859),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_982),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_983),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_989),
.B(n_972),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_987),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_983),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_1115),
.Y(n_1154)
);

OAI22x1_ASAP7_75t_L g1155 ( 
.A1(n_1145),
.A2(n_970),
.B1(n_812),
.B2(n_837),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1029),
.B(n_492),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_985),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_1115),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1112),
.B(n_910),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1031),
.B(n_848),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_984),
.B(n_954),
.Y(n_1161)
);

BUFx4f_ASAP7_75t_L g1162 ( 
.A(n_1118),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_990),
.B(n_955),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1001),
.B(n_492),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1083),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_990),
.B(n_966),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1035),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1096),
.B(n_945),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1134),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1115),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_985),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_992),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1109),
.A2(n_894),
.B1(n_861),
.B2(n_917),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_992),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1123),
.B(n_938),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1035),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1043),
.B(n_946),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1001),
.B(n_919),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_981),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1001),
.B(n_536),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1129),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1044),
.B(n_962),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_993),
.B(n_894),
.Y(n_1183)
);

NOR2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1027),
.B(n_743),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1053),
.B(n_913),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1001),
.B(n_919),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_SL g1188 ( 
.A(n_1134),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1129),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1129),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1000),
.B(n_876),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1055),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_981),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1083),
.B(n_916),
.Y(n_1194)
);

AND2x6_ASAP7_75t_L g1195 ( 
.A(n_1058),
.B(n_536),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1080),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1108),
.B(n_536),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1132),
.B(n_960),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1080),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1124),
.B(n_923),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1129),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1114),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1031),
.B(n_876),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1118),
.B(n_933),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1114),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1091),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1130),
.B(n_1142),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1054),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1085),
.B(n_960),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1108),
.B(n_536),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1130),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1063),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1063),
.B(n_933),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_986),
.Y(n_1214)
);

BUFx4f_ASAP7_75t_L g1215 ( 
.A(n_1139),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1108),
.B(n_536),
.Y(n_1216)
);

INVx4_ASAP7_75t_SL g1217 ( 
.A(n_1010),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_986),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1139),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1085),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1142),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1117),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1090),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1115),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1054),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1128),
.B(n_947),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1090),
.B(n_960),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1147),
.B(n_762),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1006),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1068),
.B(n_445),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_991),
.Y(n_1231)
);

AND2x6_ASAP7_75t_L g1232 ( 
.A(n_1058),
.B(n_620),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_SL g1233 ( 
.A(n_1038),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1137),
.B(n_968),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1038),
.A2(n_493),
.B1(n_496),
.B2(n_486),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_996),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1068),
.B(n_771),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1059),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1059),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_1038),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1110),
.B(n_793),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1115),
.Y(n_1242)
);

AND2x2_ASAP7_75t_SL g1243 ( 
.A(n_1038),
.B(n_620),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1052),
.B(n_999),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1108),
.B(n_620),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1065),
.B(n_871),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1006),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1047),
.B(n_840),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1065),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1007),
.Y(n_1250)
);

AND2x6_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_620),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1102),
.A2(n_500),
.B1(n_503),
.B2(n_498),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1054),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_991),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1066),
.B(n_871),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1102),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1007),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1126),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1105),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1071),
.B(n_1003),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1073),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1073),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_996),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1074),
.B(n_882),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1054),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1131),
.B(n_629),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1054),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1074),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1010),
.A2(n_935),
.B1(n_911),
.B2(n_714),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1075),
.B(n_882),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_980),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1072),
.B(n_971),
.C(n_969),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1008),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_1105),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1075),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1060),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1076),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1008),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1012),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1102),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1108),
.B(n_620),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1108),
.B(n_585),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1037),
.A2(n_593),
.B1(n_603),
.B2(n_589),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1012),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1009),
.B(n_976),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1121),
.B(n_963),
.Y(n_1286)
);

INVx5_ASAP7_75t_L g1287 ( 
.A(n_1060),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1076),
.B(n_889),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1078),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1014),
.Y(n_1290)
);

INVx4_ASAP7_75t_SL g1291 ( 
.A(n_1010),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1002),
.B(n_1102),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1060),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1049),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1014),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1126),
.B(n_414),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1023),
.B(n_714),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1126),
.B(n_414),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1126),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1064),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1078),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1105),
.B(n_889),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_991),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1079),
.B(n_638),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1123),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1121),
.B(n_963),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_SL g1307 ( 
.A(n_1023),
.B(n_663),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_1010),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1070),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1145),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1079),
.B(n_965),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_1010),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1015),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1081),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1015),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1123),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1140),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1081),
.B(n_965),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1018),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1064),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1082),
.B(n_670),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1082),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1064),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1084),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1113),
.Y(n_1325)
);

AND3x2_ASAP7_75t_L g1326 ( 
.A(n_1123),
.B(n_677),
.C(n_669),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1018),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1010),
.A2(n_564),
.B1(n_519),
.B2(n_582),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1084),
.B(n_799),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1010),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_991),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_995),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1020),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1113),
.B(n_891),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1020),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_995),
.B(n_801),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1093),
.B(n_416),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_997),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_997),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1092),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1161),
.B(n_998),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1159),
.B(n_998),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1271),
.B(n_1093),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1317),
.B(n_1113),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1172),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1172),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1234),
.B(n_1200),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1230),
.B(n_802),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1234),
.B(n_1004),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1201),
.B(n_1094),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1200),
.B(n_1004),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1152),
.Y(n_1352)
);

NAND2x1_ASAP7_75t_L g1353 ( 
.A(n_1267),
.B(n_1032),
.Y(n_1353)
);

NOR3xp33_ASAP7_75t_L g1354 ( 
.A(n_1294),
.B(n_866),
.C(n_862),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1177),
.A2(n_1098),
.B1(n_1100),
.B2(n_1094),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1174),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1212),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_1013),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1174),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1201),
.B(n_1148),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1201),
.B(n_1098),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1150),
.B(n_1153),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1222),
.B(n_1013),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1226),
.B(n_1016),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1243),
.A2(n_935),
.B1(n_911),
.B2(n_681),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1177),
.A2(n_1148),
.B1(n_1103),
.B2(n_1104),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1226),
.B(n_1016),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1185),
.B(n_1019),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1185),
.B(n_1019),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1201),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1211),
.B(n_1148),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1211),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1237),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1204),
.B(n_866),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1163),
.B(n_1022),
.Y(n_1375)
);

INVxp33_ASAP7_75t_L g1376 ( 
.A(n_1228),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1241),
.B(n_881),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1243),
.B(n_671),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1162),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1182),
.B(n_1100),
.Y(n_1380)
);

INVx8_ASAP7_75t_L g1381 ( 
.A(n_1188),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1162),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1238),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1182),
.B(n_1103),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1160),
.B(n_881),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1215),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1296),
.A2(n_1092),
.B(n_1033),
.C(n_1040),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1207),
.A2(n_1106),
.B1(n_1107),
.B2(n_1104),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1149),
.B(n_1106),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1221),
.B(n_1069),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1166),
.B(n_1022),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1259),
.B(n_1033),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1203),
.B(n_582),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1221),
.B(n_1069),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1258),
.A2(n_1116),
.B1(n_1122),
.B2(n_1107),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1207),
.B(n_1069),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1274),
.B(n_1040),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1325),
.B(n_1041),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1239),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1249),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1332),
.B(n_1041),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1207),
.B(n_1069),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1220),
.B(n_1046),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1165),
.B(n_1069),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1223),
.B(n_1046),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1261),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_SL g1407 ( 
.A(n_1316),
.B(n_938),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1266),
.B(n_580),
.C(n_570),
.Y(n_1408)
);

NAND2x1_ASAP7_75t_L g1409 ( 
.A(n_1267),
.B(n_1032),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1213),
.B(n_804),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1149),
.B(n_1116),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1149),
.B(n_1122),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1181),
.B(n_1127),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_SL g1414 ( 
.A(n_1173),
.B(n_433),
.C(n_413),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1179),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1179),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1193),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1262),
.Y(n_1421)
);

INVxp33_ASAP7_75t_L g1422 ( 
.A(n_1248),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1231),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1193),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1214),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1268),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1181),
.B(n_1127),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1275),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1198),
.A2(n_1136),
.B(n_1135),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1277),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1151),
.A2(n_1136),
.B1(n_1138),
.B2(n_1135),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1289),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1307),
.A2(n_1227),
.B1(n_1209),
.B2(n_1167),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1301),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1214),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1152),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1318),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_L g1438 ( 
.A(n_1269),
.B(n_1258),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1311),
.B(n_1056),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1318),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_SL g1441 ( 
.A(n_1181),
.B(n_1099),
.Y(n_1441)
);

AND2x6_ASAP7_75t_L g1442 ( 
.A(n_1150),
.B(n_1138),
.Y(n_1442)
);

INVxp33_ASAP7_75t_SL g1443 ( 
.A(n_1168),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1183),
.B(n_1141),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1151),
.A2(n_1143),
.B1(n_1144),
.B2(n_1141),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1219),
.B(n_806),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1189),
.A2(n_1144),
.B1(n_1146),
.B2(n_1143),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1176),
.B(n_1146),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1218),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1215),
.B(n_1099),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1218),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1169),
.B(n_808),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1318),
.B(n_1057),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1296),
.B(n_586),
.C(n_581),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1286),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1187),
.B(n_1057),
.Y(n_1457)
);

NAND2xp33_ASAP7_75t_L g1458 ( 
.A(n_1269),
.B(n_1036),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1338),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1192),
.B(n_1196),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_SL g1461 ( 
.A(n_1188),
.B(n_416),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1178),
.A2(n_1048),
.B(n_1034),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1314),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1229),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1199),
.B(n_1202),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1263),
.B(n_810),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1205),
.B(n_1032),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1236),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1229),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_SL g1470 ( 
.A(n_1305),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1322),
.B(n_1034),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1324),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1306),
.B(n_1244),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1186),
.B(n_1034),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1247),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1247),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1189),
.B(n_1051),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_L g1478 ( 
.A(n_1292),
.B(n_1036),
.Y(n_1478)
);

NAND2xp33_ASAP7_75t_SL g1479 ( 
.A(n_1184),
.B(n_418),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1307),
.A2(n_911),
.B1(n_679),
.B2(n_695),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1206),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1231),
.B(n_1039),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1189),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1206),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1190),
.B(n_418),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1250),
.Y(n_1486)
);

NAND2xp33_ASAP7_75t_L g1487 ( 
.A(n_1231),
.B(n_1133),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1309),
.B(n_811),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1190),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1190),
.B(n_1051),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1298),
.B(n_1051),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1256),
.B(n_1077),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1359),
.Y(n_1493)
);

NOR2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1436),
.B(n_1305),
.Y(n_1494)
);

NOR3xp33_ASAP7_75t_SL g1495 ( 
.A(n_1414),
.B(n_1316),
.C(n_446),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1352),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1347),
.B(n_1260),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1345),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1380),
.B(n_1285),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1416),
.Y(n_1500)
);

BUFx2_ASAP7_75t_SL g1501 ( 
.A(n_1370),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1378),
.A2(n_1440),
.B1(n_1437),
.B2(n_1473),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1419),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1381),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1385),
.B(n_1236),
.C(n_1310),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1380),
.B(n_1256),
.Y(n_1506)
);

CKINVDCx6p67_ASAP7_75t_R g1507 ( 
.A(n_1470),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1346),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1420),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1384),
.B(n_1280),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1422),
.B(n_1376),
.Y(n_1511)
);

NOR2x2_ASAP7_75t_L g1512 ( 
.A(n_1424),
.B(n_1297),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1378),
.A2(n_1280),
.B1(n_1299),
.B2(n_1298),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1473),
.A2(n_1194),
.B1(n_1299),
.B2(n_1233),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1384),
.B(n_1169),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1351),
.B(n_1194),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1357),
.B(n_1194),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1349),
.B(n_1337),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1356),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1368),
.B(n_1337),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1381),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1443),
.A2(n_1155),
.B1(n_444),
.B2(n_450),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1460),
.A2(n_1171),
.B(n_1153),
.C(n_1157),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1425),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1468),
.A2(n_1297),
.B1(n_1328),
.B2(n_931),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1357),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1372),
.B(n_1272),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1369),
.B(n_1339),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1459),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1373),
.A2(n_1233),
.B1(n_1252),
.B2(n_1235),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1362),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1435),
.Y(n_1532)
);

AND2x6_ASAP7_75t_L g1533 ( 
.A(n_1370),
.B(n_1171),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1463),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1456),
.B(n_1297),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1370),
.B(n_1217),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1484),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1462),
.A2(n_1157),
.B(n_1340),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1450),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1342),
.B(n_1339),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1452),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1341),
.B(n_1339),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1472),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1456),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1383),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1370),
.B(n_1217),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1433),
.B(n_1240),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1488),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1364),
.B(n_1336),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1453),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1464),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1441),
.B(n_1170),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1367),
.B(n_1250),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1399),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1400),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1406),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1423),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1444),
.B(n_1257),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1455),
.A2(n_1283),
.B1(n_1240),
.B2(n_1164),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1444),
.B(n_1257),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1348),
.B(n_907),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1421),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1469),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1418),
.A2(n_1321),
.B(n_1304),
.C(n_1164),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1475),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1433),
.B(n_1240),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1481),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1426),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1428),
.Y(n_1569)
);

AND3x2_ASAP7_75t_SL g1570 ( 
.A(n_1476),
.B(n_1278),
.C(n_1273),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1430),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1432),
.B(n_1217),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1434),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1453),
.B(n_1291),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1466),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1343),
.B(n_1273),
.Y(n_1576)
);

NOR2x2_ASAP7_75t_L g1577 ( 
.A(n_1486),
.B(n_1278),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1423),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1381),
.B(n_1330),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1454),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1548),
.B(n_1379),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1548),
.B(n_1382),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1497),
.B(n_1401),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1495),
.B(n_1386),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1497),
.B(n_1374),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1499),
.B(n_1377),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1511),
.B(n_1465),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1550),
.B(n_1496),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1575),
.B(n_1465),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1496),
.B(n_1410),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1549),
.B(n_1408),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1516),
.B(n_1389),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1516),
.B(n_1389),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1537),
.B(n_1411),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1506),
.B(n_1375),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1517),
.B(n_1411),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1550),
.B(n_1412),
.Y(n_1600)
);

AND2x2_ASAP7_75t_SL g1601 ( 
.A(n_1506),
.B(n_1438),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1510),
.B(n_1528),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1510),
.B(n_1412),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1544),
.B(n_1393),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1514),
.B(n_1344),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1544),
.B(n_1446),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1502),
.B(n_1407),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1515),
.B(n_1391),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1574),
.B(n_1483),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1580),
.B(n_1461),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1489),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1513),
.B(n_1439),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1530),
.B(n_1457),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1529),
.B(n_1343),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1527),
.B(n_1457),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_SL g1617 ( 
.A(n_1574),
.B(n_1423),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1536),
.B(n_1423),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1534),
.B(n_1358),
.Y(n_1619)
);

NAND2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1536),
.B(n_1451),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1536),
.B(n_1365),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1546),
.B(n_1365),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1527),
.B(n_1175),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1535),
.B(n_1543),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1545),
.B(n_1554),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1555),
.B(n_1363),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1556),
.B(n_1354),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1562),
.B(n_1354),
.Y(n_1628)
);

NAND2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1546),
.B(n_1480),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1546),
.B(n_1480),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1568),
.B(n_1403),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_SL g1632 ( 
.A(n_1572),
.B(n_1485),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1604),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1601),
.B(n_1523),
.Y(n_1636)
);

NAND2x1_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1533),
.Y(n_1637)
);

AND3x1_ASAP7_75t_SL g1638 ( 
.A(n_1613),
.B(n_702),
.C(n_696),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1587),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1592),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1590),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1593),
.A2(n_1525),
.B1(n_1505),
.B2(n_617),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1588),
.A2(n_617),
.B1(n_582),
.B2(n_1540),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1616),
.A2(n_1566),
.B(n_1547),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1633),
.B(n_1523),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1633),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1605),
.A2(n_1538),
.B(n_1429),
.Y(n_1648)
);

A2O1A1Ixp33_ASAP7_75t_SL g1649 ( 
.A1(n_1583),
.A2(n_1531),
.B(n_1448),
.C(n_1561),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1500),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1625),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1603),
.B(n_1542),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1594),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1589),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1619),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1586),
.A2(n_1479),
.B1(n_1566),
.B2(n_1547),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1596),
.B(n_1538),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1614),
.B(n_1576),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1607),
.A2(n_617),
.B1(n_1571),
.B2(n_1569),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1584),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1631),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1612),
.B(n_1553),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1599),
.B(n_1500),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1626),
.B(n_1498),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1609),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1615),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1611),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1627),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1611),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1531),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1600),
.Y(n_1673)
);

AO22x1_ASAP7_75t_L g1674 ( 
.A1(n_1632),
.A2(n_1533),
.B1(n_1519),
.B2(n_1508),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1621),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1624),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1623),
.Y(n_1677)
);

AOI22x1_ASAP7_75t_L g1678 ( 
.A1(n_1629),
.A2(n_1531),
.B1(n_1552),
.B2(n_1493),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1585),
.B(n_1503),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1597),
.B(n_1503),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1622),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1630),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1677),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1635),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1491),
.B(n_1552),
.Y(n_1688)
);

AO21x2_ASAP7_75t_L g1689 ( 
.A1(n_1648),
.A2(n_1645),
.B(n_1649),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1640),
.Y(n_1690)
);

INVx5_ASAP7_75t_L g1691 ( 
.A(n_1683),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1648),
.A2(n_1387),
.B(n_1610),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1650),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1677),
.Y(n_1696)
);

AOI22x1_ASAP7_75t_L g1697 ( 
.A1(n_1670),
.A2(n_1522),
.B1(n_1501),
.B2(n_1552),
.Y(n_1697)
);

BUFx4f_ASAP7_75t_L g1698 ( 
.A(n_1640),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1646),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1677),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1659),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1677),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1678),
.A2(n_1648),
.B(n_1659),
.Y(n_1703)
);

AOI22x1_ASAP7_75t_L g1704 ( 
.A1(n_1682),
.A2(n_1501),
.B1(n_1573),
.B2(n_1493),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1657),
.B(n_1591),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1677),
.Y(n_1707)
);

AOI22x1_ASAP7_75t_L g1708 ( 
.A1(n_1682),
.A2(n_1578),
.B1(n_1509),
.B2(n_1532),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1646),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1650),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1645),
.A2(n_1649),
.B(n_1658),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1659),
.A2(n_1683),
.B(n_1637),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1676),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1659),
.A2(n_1366),
.B(n_1395),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1658),
.A2(n_1559),
.B(n_1156),
.Y(n_1717)
);

BUFx12f_ASAP7_75t_L g1718 ( 
.A(n_1662),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1665),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1640),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1665),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1637),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1643),
.A2(n_1628),
.B(n_1564),
.Y(n_1723)
);

AOI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1674),
.A2(n_1156),
.B(n_1304),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1635),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1680),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1674),
.A2(n_1478),
.B(n_1458),
.Y(n_1727)
);

BUFx10_ASAP7_75t_L g1728 ( 
.A(n_1642),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1643),
.A2(n_1582),
.B(n_1581),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1637),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1683),
.A2(n_1474),
.B(n_1477),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1676),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1657),
.B(n_1509),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1650),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1635),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_SL g1736 ( 
.A(n_1641),
.B(n_1507),
.Y(n_1736)
);

AOI22x1_ASAP7_75t_L g1737 ( 
.A1(n_1682),
.A2(n_1578),
.B1(n_1524),
.B2(n_1539),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1665),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1640),
.B(n_1579),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1669),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1669),
.Y(n_1741)
);

BUFx5_ASAP7_75t_L g1742 ( 
.A(n_1663),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1669),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1682),
.B(n_1557),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1671),
.Y(n_1745)
);

AO21x2_ASAP7_75t_L g1746 ( 
.A1(n_1654),
.A2(n_1355),
.B(n_1431),
.Y(n_1746)
);

AOI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1664),
.A2(n_1321),
.B(n_1180),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1671),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1683),
.A2(n_1490),
.B(n_1471),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_SL g1750 ( 
.A1(n_1655),
.A2(n_1654),
.B(n_1664),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1655),
.A2(n_1445),
.B(n_1180),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1639),
.B(n_907),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1634),
.B(n_1524),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1653),
.Y(n_1754)
);

CKINVDCx16_ASAP7_75t_R g1755 ( 
.A(n_1671),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1640),
.B(n_1532),
.Y(n_1756)
);

INVx6_ASAP7_75t_L g1757 ( 
.A(n_1672),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1653),
.Y(n_1758)
);

NAND2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1682),
.B(n_1557),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1683),
.A2(n_1447),
.B(n_1157),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1640),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1680),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1653),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1676),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1636),
.A2(n_1487),
.B(n_1482),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1651),
.B(n_1539),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1656),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1681),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1634),
.B(n_1541),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1762),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1685),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1685),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1767),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_R g1774 ( 
.A1(n_1752),
.A2(n_689),
.B1(n_856),
.B2(n_815),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1762),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1763),
.Y(n_1776)
);

BUFx8_ASAP7_75t_SL g1777 ( 
.A(n_1718),
.Y(n_1777)
);

INVx6_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1763),
.Y(n_1779)
);

BUFx12f_ASAP7_75t_L g1780 ( 
.A(n_1767),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1687),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1718),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1723),
.A2(n_1675),
.B1(n_1639),
.B2(n_1660),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1738),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1697),
.A2(n_1675),
.B1(n_1636),
.B2(n_1680),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1687),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1762),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1738),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1697),
.A2(n_1661),
.B1(n_1644),
.B2(n_1675),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1705),
.B(n_1673),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1762),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1729),
.A2(n_1638),
.B1(n_1668),
.B2(n_1663),
.Y(n_1793)
);

CKINVDCx6p67_ASAP7_75t_R g1794 ( 
.A(n_1728),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1754),
.Y(n_1795)
);

CKINVDCx6p67_ASAP7_75t_R g1796 ( 
.A(n_1728),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1728),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1717),
.A2(n_1638),
.B1(n_1668),
.B2(n_1673),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1693),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1740),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1754),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1758),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1755),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1693),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1758),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1717),
.A2(n_1661),
.B1(n_1644),
.B2(n_1673),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1727),
.A2(n_1652),
.B(n_1660),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1719),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1728),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1717),
.A2(n_450),
.B1(n_454),
.B2(n_446),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1740),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1706),
.A2(n_1652),
.B1(n_1666),
.B2(n_1651),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1719),
.Y(n_1813)
);

INVx6_ASAP7_75t_L g1814 ( 
.A(n_1726),
.Y(n_1814)
);

OAI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1736),
.A2(n_1666),
.B1(n_1651),
.B2(n_1667),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1726),
.Y(n_1816)
);

BUFx2_ASAP7_75t_SL g1817 ( 
.A(n_1726),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1750),
.A2(n_455),
.B1(n_457),
.B2(n_454),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1711),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1721),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1698),
.A2(n_1507),
.B1(n_1579),
.B2(n_1651),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1740),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1711),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1750),
.A2(n_457),
.B1(n_458),
.B2(n_455),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1740),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1721),
.Y(n_1826)
);

BUFx12f_ASAP7_75t_L g1827 ( 
.A(n_1740),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1734),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1734),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1714),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1735),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1705),
.A2(n_460),
.B1(n_464),
.B2(n_458),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1768),
.B(n_1681),
.Y(n_1833)
);

CKINVDCx12_ASAP7_75t_R g1834 ( 
.A(n_1739),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1720),
.B(n_1681),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1712),
.A2(n_464),
.B1(n_466),
.B2(n_460),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1732),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1712),
.A2(n_467),
.B1(n_469),
.B2(n_466),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1712),
.A2(n_469),
.B1(n_470),
.B2(n_467),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1748),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1691),
.B(n_1679),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1764),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1746),
.A2(n_473),
.B1(n_475),
.B2(n_470),
.Y(n_1843)
);

INVx6_ASAP7_75t_L g1844 ( 
.A(n_1748),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1698),
.A2(n_1579),
.B1(n_1667),
.B2(n_1651),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1695),
.B(n_1699),
.Y(n_1846)
);

INVx6_ASAP7_75t_L g1847 ( 
.A(n_1748),
.Y(n_1847)
);

BUFx12f_ASAP7_75t_L g1848 ( 
.A(n_1748),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1748),
.Y(n_1849)
);

BUFx4f_ASAP7_75t_SL g1850 ( 
.A(n_1745),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1725),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1735),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1766),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1741),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1742),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1742),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1698),
.A2(n_1579),
.B1(n_1667),
.B2(n_1672),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1746),
.A2(n_475),
.B1(n_668),
.B2(n_473),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1695),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1741),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1699),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1742),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1741),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1710),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1746),
.A2(n_675),
.B1(n_676),
.B2(n_668),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1703),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1691),
.A2(n_1679),
.B1(n_676),
.B2(n_684),
.Y(n_1867)
);

NAND2x1p5_ASAP7_75t_L g1868 ( 
.A(n_1691),
.B(n_1679),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1743),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1735),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1743),
.Y(n_1871)
);

INVx6_ASAP7_75t_L g1872 ( 
.A(n_1755),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1710),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1756),
.A2(n_680),
.B1(n_684),
.B2(n_675),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1742),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1742),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1743),
.Y(n_1877)
);

CKINVDCx11_ASAP7_75t_R g1878 ( 
.A(n_1696),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1684),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1757),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1757),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1757),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1696),
.Y(n_1883)
);

BUFx12f_ASAP7_75t_L g1884 ( 
.A(n_1696),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1742),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1742),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1742),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1742),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1684),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1696),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1720),
.B(n_1761),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1696),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1769),
.B(n_1667),
.Y(n_1893)
);

INVx6_ASAP7_75t_L g1894 ( 
.A(n_1700),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1684),
.Y(n_1895)
);

INVx4_ASAP7_75t_SL g1896 ( 
.A(n_1722),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1707),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1739),
.A2(n_1667),
.B1(n_1672),
.B2(n_1504),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1756),
.A2(n_685),
.B1(n_688),
.B2(n_680),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1707),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1756),
.A2(n_688),
.B1(n_690),
.B2(n_685),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1756),
.A2(n_692),
.B1(n_693),
.B2(n_690),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1707),
.Y(n_1903)
);

BUFx10_ASAP7_75t_L g1904 ( 
.A(n_1766),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1709),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1753),
.B(n_1672),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1757),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1709),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1709),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1691),
.A2(n_693),
.B1(n_694),
.B2(n_692),
.Y(n_1910)
);

CKINVDCx11_ASAP7_75t_R g1911 ( 
.A(n_1700),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1739),
.A2(n_1672),
.B1(n_1504),
.B2(n_1521),
.Y(n_1912)
);

BUFx2_ASAP7_75t_SL g1913 ( 
.A(n_1686),
.Y(n_1913)
);

BUFx12f_ASAP7_75t_L g1914 ( 
.A(n_1700),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1761),
.B(n_1521),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1715),
.Y(n_1916)
);

INVx3_ASAP7_75t_SL g1917 ( 
.A(n_1766),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1739),
.A2(n_1388),
.B1(n_1448),
.B2(n_700),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1686),
.B(n_673),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1690),
.B(n_1694),
.Y(n_1920)
);

INVx4_ASAP7_75t_R g1921 ( 
.A(n_1715),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1891),
.B(n_1690),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1866),
.A2(n_1703),
.B(n_1713),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1800),
.Y(n_1924)
);

OA21x2_ASAP7_75t_L g1925 ( 
.A1(n_1866),
.A2(n_1876),
.B(n_1875),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1783),
.A2(n_1691),
.B(n_1708),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1771),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1800),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1780),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1807),
.A2(n_1688),
.B(n_1731),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1784),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1772),
.Y(n_1932)
);

OA21x2_ASAP7_75t_L g1933 ( 
.A1(n_1886),
.A2(n_1713),
.B(n_1731),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1836),
.A2(n_1839),
.B1(n_1838),
.B2(n_1843),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1793),
.B(n_1700),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1836),
.A2(n_1839),
.B1(n_1838),
.B2(n_1843),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1783),
.A2(n_1691),
.B(n_1708),
.Y(n_1937)
);

OA21x2_ASAP7_75t_L g1938 ( 
.A1(n_1888),
.A2(n_1749),
.B(n_1688),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1807),
.A2(n_1737),
.B(n_1704),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1860),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1793),
.B(n_1700),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1858),
.A2(n_1716),
.B(n_1749),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1781),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1786),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1812),
.A2(n_1737),
.B(n_1704),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1808),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1813),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1855),
.A2(n_1716),
.B(n_1724),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1858),
.A2(n_1865),
.B1(n_1810),
.B2(n_1790),
.Y(n_1949)
);

OAI221xp5_ASAP7_75t_L g1950 ( 
.A1(n_1832),
.A2(n_701),
.B1(n_703),
.B2(n_700),
.C(n_694),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1820),
.Y(n_1951)
);

OAI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1810),
.A2(n_703),
.B(n_706),
.C(n_701),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1865),
.A2(n_1724),
.B(n_1747),
.Y(n_1953)
);

BUFx12f_ASAP7_75t_L g1954 ( 
.A(n_1773),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1791),
.B(n_1690),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1790),
.A2(n_704),
.B(n_707),
.C(n_699),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1844),
.Y(n_1957)
);

A2O1A1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1818),
.A2(n_716),
.B(n_708),
.C(n_709),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1826),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1812),
.A2(n_1739),
.B(n_1751),
.Y(n_1960)
);

OA21x2_ASAP7_75t_L g1961 ( 
.A1(n_1856),
.A2(n_1760),
.B(n_1747),
.Y(n_1961)
);

AO31x2_ASAP7_75t_L g1962 ( 
.A1(n_1862),
.A2(n_1689),
.A3(n_1733),
.B(n_1692),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1885),
.A2(n_1760),
.B(n_1766),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1851),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1815),
.A2(n_1751),
.B(n_1617),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1859),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1861),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1830),
.B(n_1701),
.Y(n_1968)
);

AO21x2_ASAP7_75t_L g1969 ( 
.A1(n_1887),
.A2(n_1689),
.B(n_1815),
.Y(n_1969)
);

BUFx4f_ASAP7_75t_SL g1970 ( 
.A(n_1782),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1867),
.A2(n_1751),
.B(n_1689),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1818),
.A2(n_708),
.B(n_709),
.C(n_706),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1864),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1789),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1832),
.A2(n_715),
.B1(n_711),
.B2(n_604),
.C(n_607),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1835),
.B(n_1694),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1867),
.A2(n_1620),
.B(n_1765),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1799),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1851),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1871),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_SL g1981 ( 
.A1(n_1803),
.A2(n_1694),
.B1(n_1702),
.B2(n_1715),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1873),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1806),
.A2(n_1765),
.B(n_1692),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1917),
.B(n_1702),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1797),
.B(n_1702),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1787),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1806),
.A2(n_856),
.B(n_838),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1777),
.Y(n_1988)
);

AOI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1919),
.A2(n_838),
.B(n_836),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1809),
.B(n_1702),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1877),
.B(n_1701),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1800),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1795),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1804),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1785),
.A2(n_1765),
.B(n_1692),
.Y(n_1995)
);

AOI22xp33_ASAP7_75t_SL g1996 ( 
.A1(n_1872),
.A2(n_1702),
.B1(n_1730),
.B2(n_1722),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1821),
.A2(n_1759),
.B(n_1744),
.Y(n_1997)
);

OAI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1824),
.A2(n_715),
.B1(n_711),
.B2(n_611),
.C(n_618),
.Y(n_1998)
);

AOI211x1_ASAP7_75t_L g1999 ( 
.A1(n_1846),
.A2(n_818),
.B(n_820),
.C(n_814),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1819),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1823),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1801),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1785),
.A2(n_1759),
.B(n_1744),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1816),
.B(n_1701),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1829),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1802),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1837),
.B(n_1842),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1824),
.A2(n_1759),
.B1(n_1744),
.B2(n_1730),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1910),
.A2(n_1798),
.B(n_1918),
.Y(n_2009)
);

OAI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1794),
.A2(n_1722),
.B1(n_1730),
.B2(n_1701),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1912),
.A2(n_1868),
.B(n_1841),
.Y(n_2011)
);

BUFx8_ASAP7_75t_L g2012 ( 
.A(n_1915),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1910),
.A2(n_1722),
.B(n_1730),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1805),
.B(n_1722),
.Y(n_2014)
);

OAI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1874),
.A2(n_1730),
.B1(n_597),
.B2(n_619),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1798),
.A2(n_621),
.B(n_625),
.C(n_588),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1774),
.A2(n_564),
.B1(n_519),
.B2(n_822),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1828),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1776),
.Y(n_2019)
);

OAI21x1_ASAP7_75t_L g2020 ( 
.A1(n_1841),
.A2(n_1405),
.B(n_1404),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1889),
.A2(n_841),
.B(n_839),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1779),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_L g2023 ( 
.A1(n_1868),
.A2(n_1417),
.B(n_1415),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1833),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1845),
.A2(n_1397),
.B(n_1392),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1893),
.B(n_839),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1879),
.Y(n_2027)
);

INVxp67_ASAP7_75t_L g2028 ( 
.A(n_1775),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1900),
.Y(n_2029)
);

AND2x2_ASAP7_75t_SL g2030 ( 
.A(n_1816),
.B(n_1512),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1857),
.A2(n_1398),
.B(n_1371),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1831),
.B(n_841),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1844),
.Y(n_2033)
);

HB1xp67_ASAP7_75t_L g2034 ( 
.A(n_1852),
.Y(n_2034)
);

OA21x2_ASAP7_75t_L g2035 ( 
.A1(n_1903),
.A2(n_844),
.B(n_843),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1905),
.B(n_843),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1898),
.A2(n_1360),
.B(n_1449),
.Y(n_2037)
);

OAI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1883),
.A2(n_1467),
.B(n_1361),
.Y(n_2038)
);

OA21x2_ASAP7_75t_L g2039 ( 
.A1(n_1908),
.A2(n_846),
.B(n_844),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1870),
.B(n_846),
.Y(n_2040)
);

OAI21x1_ASAP7_75t_L g2041 ( 
.A1(n_1883),
.A2(n_1361),
.B(n_1350),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1872),
.A2(n_564),
.B1(n_519),
.B2(n_823),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1909),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1895),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1874),
.A2(n_826),
.B(n_824),
.Y(n_2045)
);

OAI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1840),
.A2(n_1350),
.B(n_1390),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1897),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1796),
.B(n_849),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1916),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1906),
.B(n_1863),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1863),
.B(n_1840),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1917),
.B(n_849),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1811),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1920),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1890),
.B(n_851),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1894),
.Y(n_2056)
);

AO31x2_ASAP7_75t_L g2057 ( 
.A1(n_1770),
.A2(n_828),
.A3(n_829),
.B(n_827),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1890),
.B(n_851),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1872),
.A2(n_1901),
.B1(n_1902),
.B2(n_1899),
.Y(n_2059)
);

BUFx4f_ASAP7_75t_L g2060 ( 
.A(n_1787),
.Y(n_2060)
);

OA21x2_ASAP7_75t_L g2061 ( 
.A1(n_1892),
.A2(n_853),
.B(n_852),
.Y(n_2061)
);

INVx1_ASAP7_75t_SL g2062 ( 
.A(n_1844),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1890),
.B(n_852),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1907),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_1787),
.Y(n_2065)
);

A2O1A1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_1899),
.A2(n_636),
.B(n_642),
.C(n_635),
.Y(n_2066)
);

INVx6_ASAP7_75t_L g2067 ( 
.A(n_1787),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1901),
.A2(n_1360),
.B(n_1394),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1902),
.A2(n_1154),
.B(n_1570),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1825),
.Y(n_2070)
);

CKINVDCx8_ASAP7_75t_R g2071 ( 
.A(n_1913),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1788),
.A2(n_1492),
.B(n_1541),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1881),
.A2(n_1492),
.B(n_1427),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_1817),
.A2(n_648),
.B1(n_650),
.B2(n_645),
.C(n_644),
.Y(n_2074)
);

CKINVDCx11_ASAP7_75t_R g2075 ( 
.A(n_1827),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1890),
.B(n_853),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1788),
.B(n_652),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1800),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1894),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2027),
.Y(n_2080)
);

AOI211xp5_ASAP7_75t_L g2081 ( 
.A1(n_1950),
.A2(n_654),
.B(n_659),
.C(n_653),
.Y(n_2081)
);

AOI211xp5_ASAP7_75t_L g2082 ( 
.A1(n_1950),
.A2(n_661),
.B(n_665),
.C(n_660),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1934),
.A2(n_1850),
.B1(n_1778),
.B2(n_1814),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1955),
.B(n_1853),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2005),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1936),
.A2(n_1850),
.B1(n_1778),
.B2(n_1814),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1949),
.A2(n_1853),
.B1(n_1882),
.B2(n_1880),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_2009),
.A2(n_1869),
.B1(n_1854),
.B2(n_1814),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2059),
.A2(n_1778),
.B1(n_1792),
.B2(n_1770),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_2016),
.A2(n_1792),
.B1(n_1847),
.B2(n_1894),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_1970),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2024),
.B(n_1822),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_2075),
.Y(n_2093)
);

OAI21xp33_ASAP7_75t_L g2094 ( 
.A1(n_2017),
.A2(n_424),
.B(n_419),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2015),
.A2(n_1847),
.B1(n_1848),
.B2(n_1884),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2029),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1939),
.A2(n_1849),
.B(n_1822),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_1998),
.A2(n_1975),
.B1(n_1958),
.B2(n_1972),
.C(n_2015),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_2064),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2050),
.B(n_1822),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2050),
.B(n_1822),
.Y(n_2101)
);

CKINVDCx11_ASAP7_75t_R g2102 ( 
.A(n_1954),
.Y(n_2102)
);

AO221x2_ASAP7_75t_L g2103 ( 
.A1(n_2010),
.A2(n_1921),
.B1(n_830),
.B2(n_1834),
.C(n_1896),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1998),
.A2(n_1847),
.B1(n_1911),
.B2(n_1878),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_1975),
.A2(n_1904),
.B1(n_1849),
.B2(n_1878),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2034),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1927),
.Y(n_2107)
);

OAI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2042),
.A2(n_1849),
.B1(n_428),
.B2(n_430),
.C(n_424),
.Y(n_2108)
);

OAI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_1935),
.A2(n_1911),
.B(n_428),
.C(n_430),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2054),
.B(n_1849),
.Y(n_2110)
);

AOI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_1952),
.A2(n_437),
.B(n_438),
.C(n_419),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1922),
.B(n_1904),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1964),
.B(n_973),
.Y(n_2113)
);

OAI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1977),
.A2(n_1914),
.B1(n_1896),
.B2(n_1551),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_1941),
.A2(n_973),
.B1(n_974),
.B2(n_961),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_1930),
.A2(n_1896),
.B(n_1563),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2030),
.A2(n_974),
.B1(n_977),
.B2(n_961),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_2074),
.A2(n_2008),
.B1(n_2048),
.B2(n_2052),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1932),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1956),
.A2(n_1563),
.B1(n_1565),
.B2(n_1551),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1943),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2011),
.B(n_918),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2074),
.A2(n_977),
.B1(n_978),
.B2(n_961),
.Y(n_2123)
);

INVx5_ASAP7_75t_SL g2124 ( 
.A(n_2032),
.Y(n_2124)
);

AO22x1_ASAP7_75t_L g2125 ( 
.A1(n_2012),
.A2(n_1988),
.B1(n_2053),
.B2(n_1940),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2008),
.A2(n_977),
.B1(n_978),
.B2(n_961),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2043),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2044),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_L g2129 ( 
.A1(n_1926),
.A2(n_1565),
.B(n_1329),
.Y(n_2129)
);

AOI222xp33_ASAP7_75t_L g2130 ( 
.A1(n_2045),
.A2(n_441),
.B1(n_438),
.B2(n_443),
.C1(n_440),
.C2(n_437),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1976),
.B(n_2),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2071),
.A2(n_441),
.B1(n_443),
.B2(n_440),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2007),
.B(n_918),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1981),
.A2(n_977),
.B1(n_978),
.B2(n_961),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1984),
.B(n_3),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2066),
.A2(n_459),
.B1(n_463),
.B2(n_448),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1996),
.A2(n_459),
.B1(n_463),
.B2(n_448),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1945),
.A2(n_1512),
.B1(n_471),
.B2(n_472),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1944),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_1979),
.B(n_925),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_1968),
.B(n_2007),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1946),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2028),
.B(n_4),
.Y(n_2143)
);

OA21x2_ASAP7_75t_L g2144 ( 
.A1(n_1971),
.A2(n_927),
.B(n_925),
.Y(n_2144)
);

INVx4_ASAP7_75t_SL g2145 ( 
.A(n_1929),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2070),
.B(n_2047),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_1942),
.A2(n_978),
.B1(n_977),
.B2(n_1326),
.Y(n_2147)
);

AOI221xp5_ASAP7_75t_L g2148 ( 
.A1(n_1999),
.A2(n_472),
.B1(n_474),
.B2(n_471),
.C(n_465),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_2012),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1947),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1951),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_1942),
.A2(n_978),
.B1(n_474),
.B2(n_666),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2049),
.B(n_4),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1991),
.B(n_6),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1991),
.B(n_6),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_1983),
.A2(n_672),
.B1(n_674),
.B2(n_666),
.C(n_465),
.Y(n_2156)
);

OAI221xp5_ASAP7_75t_L g2157 ( 
.A1(n_2077),
.A2(n_683),
.B1(n_686),
.B2(n_674),
.C(n_672),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1959),
.Y(n_2158)
);

AOI222xp33_ASAP7_75t_L g2159 ( 
.A1(n_2045),
.A2(n_697),
.B1(n_686),
.B2(n_705),
.C1(n_687),
.C2(n_683),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1986),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2003),
.A2(n_697),
.B1(n_705),
.B2(n_687),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1966),
.Y(n_2162)
);

BUFx2_ASAP7_75t_L g2163 ( 
.A(n_2078),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2018),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2069),
.A2(n_713),
.B1(n_1533),
.B2(n_927),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2056),
.B(n_8),
.Y(n_2166)
);

A2O1A1Ixp33_ASAP7_75t_L g2167 ( 
.A1(n_1937),
.A2(n_713),
.B(n_511),
.C(n_512),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_2067),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2069),
.A2(n_515),
.B1(n_516),
.B2(n_507),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1967),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2061),
.A2(n_1557),
.B1(n_1572),
.B2(n_534),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2079),
.B(n_1557),
.Y(n_2172)
);

AOI222xp33_ASAP7_75t_L g2173 ( 
.A1(n_1953),
.A2(n_549),
.B1(n_538),
.B2(n_550),
.C1(n_540),
.C2(n_524),
.Y(n_2173)
);

AOI21xp33_ASAP7_75t_L g2174 ( 
.A1(n_2077),
.A2(n_8),
.B(n_10),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1980),
.B(n_10),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2025),
.A2(n_1965),
.B(n_1960),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_1968),
.B(n_11),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2019),
.B(n_12),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1973),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1982),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1993),
.Y(n_2181)
);

AOI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2032),
.A2(n_567),
.B1(n_568),
.B2(n_565),
.C(n_559),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2002),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2006),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1987),
.A2(n_576),
.B1(n_577),
.B2(n_574),
.Y(n_2185)
);

NAND5xp2_ASAP7_75t_SL g2186 ( 
.A(n_2013),
.B(n_1995),
.C(n_1953),
.D(n_2068),
.E(n_2037),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2061),
.A2(n_1987),
.B1(n_1985),
.B2(n_2040),
.Y(n_2187)
);

AOI22xp33_ASAP7_75t_L g2188 ( 
.A1(n_2040),
.A2(n_2026),
.B1(n_1990),
.B2(n_2031),
.Y(n_2188)
);

OAI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_2026),
.A2(n_1557),
.B1(n_587),
.B2(n_590),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2067),
.Y(n_2190)
);

AOI22xp33_ASAP7_75t_SL g2191 ( 
.A1(n_1997),
.A2(n_591),
.B1(n_595),
.B2(n_584),
.Y(n_2191)
);

OAI221xp5_ASAP7_75t_L g2192 ( 
.A1(n_2036),
.A2(n_606),
.B1(n_609),
.B2(n_601),
.C(n_599),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2036),
.A2(n_2033),
.B1(n_1957),
.B2(n_2055),
.Y(n_2193)
);

BUFx4f_ASAP7_75t_SL g2194 ( 
.A(n_1986),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2060),
.A2(n_2062),
.B1(n_2004),
.B2(n_2051),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_1924),
.Y(n_2196)
);

OAI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2055),
.A2(n_622),
.B(n_614),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_1948),
.A2(n_1427),
.B(n_1413),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2022),
.Y(n_2199)
);

OAI22xp33_ASAP7_75t_L g2200 ( 
.A1(n_2076),
.A2(n_628),
.B1(n_630),
.B2(n_626),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1986),
.Y(n_2201)
);

OA21x2_ASAP7_75t_L g2202 ( 
.A1(n_2014),
.A2(n_646),
.B(n_632),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2065),
.Y(n_2203)
);

AOI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_2058),
.A2(n_1533),
.B1(n_1442),
.B2(n_656),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2058),
.B(n_891),
.C(n_934),
.Y(n_2205)
);

BUFx5_ASAP7_75t_L g2206 ( 
.A(n_1923),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_1969),
.A2(n_1533),
.B1(n_1572),
.B2(n_14),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2051),
.B(n_12),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2063),
.A2(n_2076),
.B1(n_2062),
.B2(n_1969),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_1924),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2060),
.A2(n_1570),
.B1(n_1577),
.B2(n_1402),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2014),
.B(n_13),
.Y(n_2212)
);

OR2x6_ASAP7_75t_L g2213 ( 
.A(n_2004),
.B(n_1413),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1928),
.B(n_14),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1931),
.Y(n_2215)
);

OAI211xp5_ASAP7_75t_L g2216 ( 
.A1(n_2063),
.A2(n_1989),
.B(n_1978),
.C(n_1974),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1994),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_1928),
.A2(n_1570),
.B1(n_1577),
.B2(n_1396),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2065),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2000),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2001),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2065),
.A2(n_1255),
.B1(n_1264),
.B2(n_1246),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_1925),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1992),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1992),
.B(n_1962),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1925),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2073),
.A2(n_1533),
.B1(n_1442),
.B2(n_1362),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_SL g2228 ( 
.A1(n_2021),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2020),
.A2(n_1442),
.B1(n_1362),
.B2(n_1288),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1963),
.B(n_16),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2021),
.A2(n_1442),
.B1(n_1362),
.B2(n_1270),
.Y(n_2231)
);

AOI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_2035),
.A2(n_1442),
.B1(n_1362),
.B2(n_1284),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2035),
.A2(n_1334),
.B(n_1302),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2039),
.A2(n_1284),
.B1(n_1290),
.B2(n_1279),
.Y(n_2234)
);

AO31x2_ASAP7_75t_L g2235 ( 
.A1(n_1933),
.A2(n_1290),
.A3(n_1295),
.B(n_1279),
.Y(n_2235)
);

AOI221xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2057),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.C(n_27),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_2023),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_2164),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2122),
.B(n_2230),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2107),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2141),
.B(n_2177),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2226),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_2122),
.B(n_2057),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2101),
.B(n_1962),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_2102),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2119),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_SL g2247 ( 
.A1(n_2098),
.A2(n_2039),
.B1(n_1963),
.B2(n_1933),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2106),
.B(n_1962),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2103),
.A2(n_2046),
.B1(n_2041),
.B2(n_2038),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2163),
.B(n_1923),
.Y(n_2250)
);

AO21x2_ASAP7_75t_L g2251 ( 
.A1(n_2223),
.A2(n_2072),
.B(n_2057),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2121),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2139),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2093),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2196),
.B(n_1938),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2142),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2150),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_2093),
.Y(n_2258)
);

INVx2_ASAP7_75t_SL g2259 ( 
.A(n_2160),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2151),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2206),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_2093),
.Y(n_2262)
);

BUFx4f_ASAP7_75t_SL g2263 ( 
.A(n_2099),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2085),
.B(n_1961),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_2103),
.A2(n_1961),
.B1(n_1938),
.B2(n_1313),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2206),
.Y(n_2266)
);

NOR2x1_ASAP7_75t_L g2267 ( 
.A(n_2149),
.B(n_1197),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2206),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2113),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2168),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2162),
.Y(n_2271)
);

AO21x2_ASAP7_75t_L g2272 ( 
.A1(n_2225),
.A2(n_1210),
.B(n_1197),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2092),
.B(n_24),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2080),
.B(n_27),
.Y(n_2274)
);

INVx4_ASAP7_75t_R g2275 ( 
.A(n_2091),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2206),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2146),
.B(n_29),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2170),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2140),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2168),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2210),
.B(n_29),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2179),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2180),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2206),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2158),
.Y(n_2285)
);

INVx8_ASAP7_75t_L g2286 ( 
.A(n_2214),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_2084),
.B(n_30),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2096),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2127),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2215),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2176),
.B(n_30),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2156),
.A2(n_1313),
.B1(n_1315),
.B2(n_1295),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2181),
.Y(n_2293)
);

INVxp67_ASAP7_75t_L g2294 ( 
.A(n_2212),
.Y(n_2294)
);

INVx5_ASAP7_75t_L g2295 ( 
.A(n_2214),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2208),
.B(n_31),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2183),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_SL g2298 ( 
.A1(n_2202),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2210),
.B(n_35),
.Y(n_2299)
);

AND2x2_ASAP7_75t_SL g2300 ( 
.A(n_2202),
.B(n_37),
.Y(n_2300)
);

AND2x2_ASAP7_75t_SL g2301 ( 
.A(n_2161),
.B(n_39),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2224),
.B(n_40),
.Y(n_2302)
);

AOI221xp5_ASAP7_75t_L g2303 ( 
.A1(n_2186),
.A2(n_44),
.B1(n_41),
.B2(n_42),
.C(n_45),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2097),
.B(n_44),
.Y(n_2304)
);

NOR2x1_ASAP7_75t_SL g2305 ( 
.A(n_2195),
.B(n_45),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_2201),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2184),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_2219),
.B(n_47),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_2160),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2199),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2112),
.B(n_47),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2190),
.B(n_49),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_2203),
.B(n_49),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2220),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2217),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2100),
.B(n_50),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2221),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2110),
.B(n_50),
.Y(n_2318)
);

NOR2x1_ASAP7_75t_L g2319 ( 
.A(n_2216),
.B(n_1210),
.Y(n_2319)
);

AO31x2_ASAP7_75t_L g2320 ( 
.A1(n_2089),
.A2(n_55),
.A3(n_52),
.B(n_53),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2128),
.B(n_52),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2153),
.Y(n_2322)
);

INVx8_ASAP7_75t_L g2323 ( 
.A(n_2213),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2203),
.B(n_56),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2209),
.B(n_57),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2133),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2178),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2237),
.B(n_2088),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2160),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2143),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2116),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2154),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2193),
.B(n_58),
.Y(n_2333)
);

AOI22xp33_ASAP7_75t_L g2334 ( 
.A1(n_2130),
.A2(n_1319),
.B1(n_1327),
.B2(n_1315),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2166),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_2194),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2235),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2235),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2155),
.B(n_59),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2129),
.B(n_59),
.Y(n_2340)
);

BUFx3_ASAP7_75t_L g2341 ( 
.A(n_2135),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2131),
.B(n_61),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_R g2343 ( 
.A(n_2118),
.B(n_61),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2235),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2172),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2145),
.Y(n_2346)
);

OAI211xp5_ASAP7_75t_L g2347 ( 
.A1(n_2081),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2124),
.B(n_63),
.Y(n_2348)
);

AOI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2174),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2172),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2198),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2124),
.B(n_67),
.Y(n_2352)
);

AOI222xp33_ASAP7_75t_L g2353 ( 
.A1(n_2094),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.C1(n_72),
.C2(n_73),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2145),
.B(n_75),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_2125),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2213),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2087),
.B(n_75),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2104),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2213),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2083),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2175),
.B(n_76),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2188),
.B(n_2187),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2086),
.B(n_2144),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2144),
.B(n_79),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2242),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2303),
.A2(n_2159),
.B1(n_2173),
.B2(n_2152),
.Y(n_2366)
);

BUFx3_ASAP7_75t_L g2367 ( 
.A(n_2258),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2242),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2261),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2310),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_2254),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2261),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2327),
.B(n_2279),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_L g2374 ( 
.A(n_2343),
.B(n_2104),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2240),
.Y(n_2375)
);

OAI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2300),
.A2(n_2167),
.B(n_2169),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2239),
.B(n_2095),
.Y(n_2377)
);

AOI21xp33_ASAP7_75t_SL g2378 ( 
.A1(n_2355),
.A2(n_2138),
.B(n_2114),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2246),
.Y(n_2379)
);

INVxp67_ASAP7_75t_L g2380 ( 
.A(n_2269),
.Y(n_2380)
);

INVxp67_ASAP7_75t_SL g2381 ( 
.A(n_2305),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2266),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2238),
.Y(n_2383)
);

A2O1A1Ixp33_ASAP7_75t_L g2384 ( 
.A1(n_2347),
.A2(n_2082),
.B(n_2081),
.C(n_2094),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_2239),
.B(n_2207),
.Y(n_2385)
);

OAI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2300),
.A2(n_2169),
.B(n_2191),
.Y(n_2386)
);

AO31x2_ASAP7_75t_L g2387 ( 
.A1(n_2266),
.A2(n_2234),
.A3(n_2171),
.B(n_2090),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2327),
.B(n_2236),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2239),
.B(n_2105),
.Y(n_2389)
);

O2A1O1Ixp33_ASAP7_75t_L g2390 ( 
.A1(n_2291),
.A2(n_2082),
.B(n_2108),
.C(n_2157),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2362),
.A2(n_2228),
.B(n_2109),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2252),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2268),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2253),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2256),
.Y(n_2395)
);

OAI21xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2353),
.A2(n_2136),
.B(n_2148),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2257),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2268),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2346),
.Y(n_2399)
);

AO21x2_ASAP7_75t_L g2400 ( 
.A1(n_2276),
.A2(n_2185),
.B(n_2205),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2260),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2276),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2358),
.A2(n_2228),
.B(n_2189),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2262),
.Y(n_2404)
);

AOI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2360),
.A2(n_2236),
.B(n_2137),
.Y(n_2405)
);

AOI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2343),
.A2(n_2192),
.B1(n_2165),
.B2(n_2123),
.Y(n_2406)
);

INVxp67_ASAP7_75t_SL g2407 ( 
.A(n_2304),
.Y(n_2407)
);

INVxp67_ASAP7_75t_L g2408 ( 
.A(n_2241),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2290),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2284),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2350),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2298),
.A2(n_2245),
.B(n_2349),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2345),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_2301),
.A2(n_2197),
.B1(n_2147),
.B2(n_2117),
.Y(n_2414)
);

OAI21xp33_ASAP7_75t_L g2415 ( 
.A1(n_2247),
.A2(n_2115),
.B(n_2111),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2355),
.B(n_2222),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2270),
.B(n_2280),
.Y(n_2417)
);

BUFx3_ASAP7_75t_L g2418 ( 
.A(n_2258),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2345),
.Y(n_2419)
);

OAI221xp5_ASAP7_75t_L g2420 ( 
.A1(n_2294),
.A2(n_2111),
.B1(n_2132),
.B2(n_2182),
.C(n_2185),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2284),
.Y(n_2421)
);

AOI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2328),
.A2(n_2211),
.B1(n_2200),
.B2(n_2218),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2285),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_R g2424 ( 
.A(n_2254),
.B(n_80),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2262),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2271),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2280),
.B(n_2126),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2285),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2278),
.Y(n_2429)
);

A2O1A1Ixp33_ASAP7_75t_L g2430 ( 
.A1(n_2301),
.A2(n_2134),
.B(n_2227),
.C(n_2204),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2357),
.A2(n_2205),
.B1(n_2120),
.B2(n_2229),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2322),
.B(n_2231),
.Y(n_2432)
);

OAI21xp33_ASAP7_75t_SL g2433 ( 
.A1(n_2328),
.A2(n_2232),
.B(n_2233),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2304),
.A2(n_1327),
.B1(n_1333),
.B2(n_1319),
.Y(n_2434)
);

OR2x6_ASAP7_75t_L g2435 ( 
.A(n_2262),
.B(n_80),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2282),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2326),
.B(n_81),
.Y(n_2437)
);

OA21x2_ASAP7_75t_L g2438 ( 
.A1(n_2264),
.A2(n_1245),
.B(n_1216),
.Y(n_2438)
);

A2O1A1Ixp33_ASAP7_75t_L g2439 ( 
.A1(n_2354),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2288),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2288),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2289),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2319),
.A2(n_82),
.B(n_83),
.Y(n_2443)
);

INVx2_ASAP7_75t_SL g2444 ( 
.A(n_2254),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2357),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2304),
.A2(n_85),
.B(n_87),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2254),
.Y(n_2447)
);

NAND4xp25_ASAP7_75t_L g2448 ( 
.A(n_2354),
.B(n_89),
.C(n_87),
.D(n_88),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2283),
.Y(n_2449)
);

BUFx3_ASAP7_75t_L g2450 ( 
.A(n_2306),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2293),
.Y(n_2451)
);

OAI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2325),
.A2(n_88),
.B(n_89),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2316),
.B(n_91),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2322),
.B(n_91),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_SL g2455 ( 
.A1(n_2325),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_2455)
);

OA21x2_ASAP7_75t_L g2456 ( 
.A1(n_2351),
.A2(n_1245),
.B(n_1216),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2331),
.Y(n_2457)
);

HB1xp67_ASAP7_75t_L g2458 ( 
.A(n_2289),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2297),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2307),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2255),
.Y(n_2461)
);

AO31x2_ASAP7_75t_L g2462 ( 
.A1(n_2329),
.A2(n_96),
.A3(n_94),
.B(n_95),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2255),
.Y(n_2463)
);

INVx2_ASAP7_75t_SL g2464 ( 
.A(n_2275),
.Y(n_2464)
);

AOI21xp33_ASAP7_75t_L g2465 ( 
.A1(n_2363),
.A2(n_96),
.B(n_97),
.Y(n_2465)
);

AO21x2_ASAP7_75t_L g2466 ( 
.A1(n_2281),
.A2(n_1281),
.B(n_98),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2250),
.Y(n_2467)
);

OAI21x1_ASAP7_75t_L g2468 ( 
.A1(n_2331),
.A2(n_99),
.B(n_101),
.Y(n_2468)
);

OAI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_2295),
.A2(n_104),
.B1(n_101),
.B2(n_102),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2250),
.Y(n_2470)
);

CKINVDCx14_ASAP7_75t_R g2471 ( 
.A(n_2336),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2314),
.Y(n_2472)
);

HB1xp67_ASAP7_75t_L g2473 ( 
.A(n_2356),
.Y(n_2473)
);

OAI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2267),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_2474)
);

AND2x4_ASAP7_75t_L g2475 ( 
.A(n_2243),
.B(n_105),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2331),
.Y(n_2476)
);

OA21x2_ASAP7_75t_L g2477 ( 
.A1(n_2248),
.A2(n_2338),
.B(n_2337),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2370),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2375),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2399),
.B(n_2359),
.Y(n_2480)
);

INVx1_ASAP7_75t_SL g2481 ( 
.A(n_2424),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2471),
.A2(n_2295),
.B1(n_2249),
.B2(n_2323),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2477),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2471),
.A2(n_2295),
.B1(n_2323),
.B2(n_2341),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2373),
.B(n_2315),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2383),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2425),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2417),
.B(n_2259),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2477),
.Y(n_2489)
);

OR2x2_ASAP7_75t_L g2490 ( 
.A(n_2388),
.B(n_2317),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_2374),
.A2(n_2323),
.B1(n_2363),
.B2(n_2340),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2473),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2409),
.B(n_2320),
.Y(n_2493)
);

OAI33xp33_ASAP7_75t_L g2494 ( 
.A1(n_2416),
.A2(n_2330),
.A3(n_2321),
.B1(n_2296),
.B2(n_2273),
.B3(n_2287),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2379),
.Y(n_2495)
);

INVx4_ASAP7_75t_L g2496 ( 
.A(n_2435),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2407),
.B(n_2259),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2392),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2377),
.B(n_2248),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2464),
.B(n_2263),
.Y(n_2500)
);

INVx4_ASAP7_75t_L g2501 ( 
.A(n_2435),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2413),
.B(n_2309),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2477),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2374),
.A2(n_2333),
.B(n_2286),
.Y(n_2504)
);

INVx5_ASAP7_75t_SL g2505 ( 
.A(n_2435),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_R g2506 ( 
.A(n_2450),
.B(n_2263),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2450),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2411),
.B(n_2320),
.Y(n_2508)
);

BUFx2_ASAP7_75t_L g2509 ( 
.A(n_2404),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2381),
.A2(n_2243),
.B1(n_2323),
.B2(n_2340),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2475),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2419),
.B(n_2309),
.Y(n_2512)
);

OAI31xp33_ASAP7_75t_L g2513 ( 
.A1(n_2405),
.A2(n_2333),
.A3(n_2352),
.B(n_2348),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2475),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2475),
.B(n_2335),
.Y(n_2515)
);

INVx2_ASAP7_75t_SL g2516 ( 
.A(n_2367),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_2404),
.Y(n_2517)
);

AOI211xp5_ASAP7_75t_L g2518 ( 
.A1(n_2386),
.A2(n_2376),
.B(n_2378),
.C(n_2403),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2391),
.B(n_2335),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2389),
.B(n_2309),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2385),
.B(n_2447),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2447),
.B(n_2309),
.Y(n_2522)
);

INVx5_ASAP7_75t_SL g2523 ( 
.A(n_2466),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2447),
.B(n_2295),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2476),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2404),
.B(n_2341),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2433),
.B(n_2243),
.Y(n_2527)
);

A2O1A1Ixp33_ASAP7_75t_L g2528 ( 
.A1(n_2384),
.A2(n_2348),
.B(n_2352),
.C(n_2361),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2476),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2394),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2408),
.B(n_2281),
.Y(n_2531)
);

OAI211xp5_ASAP7_75t_L g2532 ( 
.A1(n_2424),
.A2(n_2364),
.B(n_2299),
.C(n_2277),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2367),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2416),
.A2(n_2340),
.B1(n_2286),
.B2(n_2332),
.Y(n_2534)
);

INVx4_ASAP7_75t_L g2535 ( 
.A(n_2418),
.Y(n_2535)
);

INVxp67_ASAP7_75t_L g2536 ( 
.A(n_2418),
.Y(n_2536)
);

AOI22xp33_ASAP7_75t_L g2537 ( 
.A1(n_2415),
.A2(n_2286),
.B1(n_2364),
.B2(n_2313),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2395),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2440),
.B(n_2320),
.Y(n_2539)
);

AO21x2_ASAP7_75t_L g2540 ( 
.A1(n_2465),
.A2(n_2299),
.B(n_2324),
.Y(n_2540)
);

OAI211xp5_ASAP7_75t_SL g2541 ( 
.A1(n_2412),
.A2(n_2318),
.B(n_2265),
.C(n_2244),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2380),
.B(n_2316),
.Y(n_2542)
);

NOR2x1_ASAP7_75t_SL g2543 ( 
.A(n_2400),
.B(n_2277),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2397),
.Y(n_2544)
);

AO21x2_ASAP7_75t_L g2545 ( 
.A1(n_2439),
.A2(n_2324),
.B(n_2312),
.Y(n_2545)
);

BUFx2_ASAP7_75t_SL g2546 ( 
.A(n_2371),
.Y(n_2546)
);

INVx2_ASAP7_75t_SL g2547 ( 
.A(n_2371),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2444),
.B(n_2311),
.Y(n_2548)
);

OAI31xp33_ASAP7_75t_SL g2549 ( 
.A1(n_2452),
.A2(n_2313),
.A3(n_2361),
.B(n_2308),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2401),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2457),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2457),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2461),
.B(n_2311),
.Y(n_2553)
);

INVx4_ASAP7_75t_L g2554 ( 
.A(n_2454),
.Y(n_2554)
);

AO21x2_ASAP7_75t_L g2555 ( 
.A1(n_2439),
.A2(n_2312),
.B(n_2274),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2461),
.B(n_2302),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2453),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2457),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2426),
.Y(n_2559)
);

INVx4_ASAP7_75t_L g2560 ( 
.A(n_2466),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2429),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2463),
.B(n_2302),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2463),
.B(n_2274),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2467),
.B(n_2320),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2436),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2506),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2520),
.B(n_2458),
.Y(n_2567)
);

NOR3xp33_ASAP7_75t_SL g2568 ( 
.A(n_2484),
.B(n_2448),
.C(n_2474),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2492),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2520),
.B(n_2467),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2486),
.Y(n_2571)
);

INVx5_ASAP7_75t_L g2572 ( 
.A(n_2560),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2507),
.B(n_2521),
.Y(n_2573)
);

AO21x1_ASAP7_75t_L g2574 ( 
.A1(n_2518),
.A2(n_2469),
.B(n_2443),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2519),
.B(n_2432),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2507),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2507),
.B(n_2470),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2515),
.B(n_2437),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2521),
.B(n_2470),
.Y(n_2579)
);

AND2x4_ASAP7_75t_SL g2580 ( 
.A(n_2496),
.B(n_2501),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2528),
.B(n_2446),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2480),
.B(n_2423),
.Y(n_2582)
);

NOR2x1_ASAP7_75t_L g2583 ( 
.A(n_2560),
.B(n_2313),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2480),
.B(n_2488),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2487),
.Y(n_2585)
);

INVx2_ASAP7_75t_SL g2586 ( 
.A(n_2509),
.Y(n_2586)
);

NOR2x1_ASAP7_75t_L g2587 ( 
.A(n_2560),
.B(n_2308),
.Y(n_2587)
);

NAND2x1p5_ASAP7_75t_L g2588 ( 
.A(n_2496),
.B(n_2468),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2535),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2487),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2542),
.B(n_2472),
.Y(n_2591)
);

NAND2x1_ASAP7_75t_L g2592 ( 
.A(n_2496),
.B(n_2365),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2509),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2517),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2528),
.B(n_2427),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2478),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2501),
.B(n_2423),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2488),
.B(n_2428),
.Y(n_2598)
);

HB1xp67_ASAP7_75t_L g2599 ( 
.A(n_2497),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2517),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2479),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2517),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_R g2603 ( 
.A(n_2481),
.B(n_2445),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2495),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2497),
.B(n_2428),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2498),
.Y(n_2606)
);

INVxp67_ASAP7_75t_L g2607 ( 
.A(n_2546),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2526),
.B(n_2441),
.Y(n_2608)
);

INVxp67_ASAP7_75t_L g2609 ( 
.A(n_2546),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2526),
.B(n_2441),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2501),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2522),
.B(n_2442),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2545),
.B(n_2449),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2530),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2535),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2545),
.B(n_2451),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2522),
.B(n_2442),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2535),
.B(n_2516),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2516),
.B(n_2365),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2538),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2533),
.B(n_2368),
.Y(n_2621)
);

NAND2x1p5_ASAP7_75t_L g2622 ( 
.A(n_2524),
.B(n_2468),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2483),
.Y(n_2623)
);

NOR2xp67_ASAP7_75t_L g2624 ( 
.A(n_2533),
.B(n_2368),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2545),
.B(n_2554),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2499),
.B(n_2387),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2547),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2544),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2550),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2500),
.Y(n_2630)
);

INVx2_ASAP7_75t_SL g2631 ( 
.A(n_2524),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2559),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2561),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2483),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2565),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2554),
.B(n_2459),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2489),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2547),
.B(n_2460),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2499),
.B(n_2387),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2554),
.B(n_2513),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2563),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2511),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2563),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2511),
.B(n_2369),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2502),
.B(n_2387),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2514),
.B(n_2455),
.Y(n_2646)
);

AND2x4_ASAP7_75t_SL g2647 ( 
.A(n_2548),
.B(n_2514),
.Y(n_2647)
);

INVxp67_ASAP7_75t_L g2648 ( 
.A(n_2573),
.Y(n_2648)
);

XNOR2x2_ASAP7_75t_L g2649 ( 
.A(n_2581),
.B(n_2504),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2584),
.B(n_2573),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2572),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2572),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2572),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2584),
.B(n_2505),
.Y(n_2654)
);

NOR4xp25_ASAP7_75t_L g2655 ( 
.A(n_2595),
.B(n_2536),
.C(n_2557),
.D(n_2384),
.Y(n_2655)
);

INVx1_ASAP7_75t_SL g2656 ( 
.A(n_2566),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2572),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2599),
.B(n_2505),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2586),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2586),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2618),
.B(n_2630),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_2647),
.Y(n_2662)
);

NOR2x1_ASAP7_75t_R g2663 ( 
.A(n_2630),
.B(n_2308),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2623),
.Y(n_2664)
);

BUFx3_ASAP7_75t_L g2665 ( 
.A(n_2618),
.Y(n_2665)
);

CKINVDCx16_ASAP7_75t_R g2666 ( 
.A(n_2603),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2647),
.B(n_2502),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_SL g2668 ( 
.A(n_2587),
.B(n_2494),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2567),
.B(n_2512),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2623),
.Y(n_2670)
);

XOR2x2_ASAP7_75t_L g2671 ( 
.A(n_2640),
.B(n_2543),
.Y(n_2671)
);

NOR3xp33_ASAP7_75t_L g2672 ( 
.A(n_2607),
.B(n_2482),
.C(n_2396),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2634),
.Y(n_2673)
);

NAND4xp75_ASAP7_75t_L g2674 ( 
.A(n_2574),
.B(n_2625),
.C(n_2583),
.D(n_2568),
.Y(n_2674)
);

NAND4xp75_ASAP7_75t_L g2675 ( 
.A(n_2574),
.B(n_2527),
.C(n_2564),
.D(n_2505),
.Y(n_2675)
);

XNOR2xp5_ASAP7_75t_L g2676 ( 
.A(n_2580),
.B(n_2366),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_SL g2677 ( 
.A(n_2609),
.B(n_2512),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2572),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2589),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2567),
.B(n_2505),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2634),
.Y(n_2681)
);

XNOR2xp5_ASAP7_75t_L g2682 ( 
.A(n_2580),
.B(n_2366),
.Y(n_2682)
);

NAND3xp33_ASAP7_75t_L g2683 ( 
.A(n_2613),
.B(n_2445),
.C(n_2493),
.Y(n_2683)
);

NAND4xp75_ASAP7_75t_SL g2684 ( 
.A(n_2570),
.B(n_2564),
.C(n_2438),
.D(n_2531),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2637),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2585),
.B(n_2531),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2570),
.B(n_2553),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2590),
.B(n_2548),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2611),
.B(n_2537),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2592),
.Y(n_2690)
);

NAND4xp75_ASAP7_75t_L g2691 ( 
.A(n_2616),
.B(n_2510),
.C(n_2523),
.D(n_2422),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2611),
.B(n_2555),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2589),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2624),
.Y(n_2694)
);

NAND4xp75_ASAP7_75t_L g2695 ( 
.A(n_2615),
.B(n_2523),
.C(n_2489),
.D(n_2503),
.Y(n_2695)
);

OAI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2646),
.A2(n_2523),
.B1(n_2491),
.B2(n_2534),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2579),
.B(n_2553),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2637),
.Y(n_2698)
);

XOR2x2_ASAP7_75t_L g2699 ( 
.A(n_2588),
.B(n_2555),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2579),
.B(n_2556),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2576),
.B(n_2555),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2642),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2589),
.Y(n_2703)
);

NAND4xp75_ASAP7_75t_L g2704 ( 
.A(n_2615),
.B(n_2523),
.C(n_2503),
.D(n_2342),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2582),
.B(n_2562),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2602),
.Y(n_2706)
);

HB1xp67_ASAP7_75t_L g2707 ( 
.A(n_2627),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2576),
.B(n_2642),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2641),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2661),
.B(n_2643),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2707),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_SL g2712 ( 
.A(n_2666),
.B(n_2631),
.Y(n_2712)
);

INVxp67_ASAP7_75t_SL g2713 ( 
.A(n_2694),
.Y(n_2713)
);

AND2x4_ASAP7_75t_SL g2714 ( 
.A(n_2661),
.B(n_2569),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2690),
.Y(n_2715)
);

OR2x2_ASAP7_75t_L g2716 ( 
.A(n_2656),
.B(n_2575),
.Y(n_2716)
);

INVx4_ASAP7_75t_L g2717 ( 
.A(n_2678),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2690),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2700),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2665),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2700),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2688),
.B(n_2571),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2665),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2655),
.B(n_2593),
.Y(n_2724)
);

INVx2_ASAP7_75t_SL g2725 ( 
.A(n_2667),
.Y(n_2725)
);

INVx1_ASAP7_75t_SL g2726 ( 
.A(n_2699),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2686),
.B(n_2578),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2705),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_L g2729 ( 
.A(n_2654),
.B(n_2532),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2650),
.Y(n_2730)
);

OAI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2675),
.A2(n_2588),
.B1(n_2622),
.B2(n_2493),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2650),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2705),
.Y(n_2733)
);

NAND3xp33_ASAP7_75t_L g2734 ( 
.A(n_2668),
.B(n_2549),
.C(n_2636),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2667),
.B(n_2631),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2697),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2677),
.B(n_2603),
.Y(n_2737)
);

INVxp67_ASAP7_75t_L g2738 ( 
.A(n_2663),
.Y(n_2738)
);

NAND2xp33_ASAP7_75t_SL g2739 ( 
.A(n_2669),
.B(n_2540),
.Y(n_2739)
);

OR2x2_ASAP7_75t_L g2740 ( 
.A(n_2648),
.B(n_2591),
.Y(n_2740)
);

AOI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2675),
.A2(n_2541),
.B1(n_2540),
.B2(n_2598),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2669),
.B(n_2598),
.Y(n_2742)
);

INVx1_ASAP7_75t_SL g2743 ( 
.A(n_2699),
.Y(n_2743)
);

OAI21xp33_ASAP7_75t_L g2744 ( 
.A1(n_2671),
.A2(n_2582),
.B(n_2608),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2697),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2674),
.B(n_2596),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2674),
.B(n_2601),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2687),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2691),
.A2(n_2622),
.B1(n_2508),
.B2(n_2406),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2702),
.B(n_2490),
.Y(n_2750)
);

HB1xp67_ASAP7_75t_L g2751 ( 
.A(n_2687),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2678),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2680),
.B(n_2556),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2689),
.B(n_2490),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2676),
.B(n_2682),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2664),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2751),
.Y(n_2757)
);

OAI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2749),
.A2(n_2691),
.B(n_2671),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_2752),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2730),
.B(n_2708),
.Y(n_2760)
);

OAI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2734),
.A2(n_2749),
.B1(n_2741),
.B2(n_2724),
.Y(n_2761)
);

O2A1O1Ixp5_ASAP7_75t_L g2762 ( 
.A1(n_2731),
.A2(n_2683),
.B(n_2696),
.C(n_2658),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2731),
.A2(n_2701),
.B(n_2693),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2752),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2752),
.Y(n_2765)
);

OAI221xp5_ASAP7_75t_L g2766 ( 
.A1(n_2734),
.A2(n_2672),
.B1(n_2676),
.B2(n_2682),
.C(n_2662),
.Y(n_2766)
);

OAI21xp33_ASAP7_75t_L g2767 ( 
.A1(n_2712),
.A2(n_2744),
.B(n_2724),
.Y(n_2767)
);

AOI21xp33_ASAP7_75t_L g2768 ( 
.A1(n_2712),
.A2(n_2680),
.B(n_2692),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2717),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2713),
.B(n_2659),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2737),
.B(n_2660),
.C(n_2709),
.Y(n_2771)
);

XNOR2xp5_ASAP7_75t_L g2772 ( 
.A(n_2753),
.B(n_2649),
.Y(n_2772)
);

INVxp67_ASAP7_75t_L g2773 ( 
.A(n_2735),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2732),
.B(n_2709),
.Y(n_2774)
);

A2O1A1Ixp33_ASAP7_75t_L g2775 ( 
.A1(n_2726),
.A2(n_2649),
.B(n_2508),
.C(n_2390),
.Y(n_2775)
);

NAND3xp33_ASAP7_75t_L g2776 ( 
.A(n_2746),
.B(n_2747),
.C(n_2755),
.Y(n_2776)
);

OAI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2746),
.A2(n_2704),
.B(n_2695),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2717),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2719),
.Y(n_2779)
);

INVx2_ASAP7_75t_SL g2780 ( 
.A(n_2735),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_SL g2781 ( 
.A(n_2716),
.B(n_2597),
.Y(n_2781)
);

AOI21xp33_ASAP7_75t_L g2782 ( 
.A1(n_2729),
.A2(n_2738),
.B(n_2726),
.Y(n_2782)
);

AOI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2743),
.A2(n_2681),
.B1(n_2685),
.B2(n_2673),
.C(n_2670),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2725),
.B(n_2679),
.Y(n_2784)
);

AOI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2747),
.A2(n_2693),
.B(n_2679),
.Y(n_2785)
);

OAI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2743),
.A2(n_2704),
.B1(n_2695),
.B2(n_2539),
.Y(n_2786)
);

OAI22xp33_ASAP7_75t_L g2787 ( 
.A1(n_2754),
.A2(n_2539),
.B1(n_2602),
.B2(n_2420),
.Y(n_2787)
);

AOI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2742),
.A2(n_2540),
.B1(n_2577),
.B2(n_2608),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2721),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2728),
.Y(n_2790)
);

OAI221xp5_ASAP7_75t_SL g2791 ( 
.A1(n_2722),
.A2(n_2706),
.B1(n_2639),
.B2(n_2626),
.C(n_2703),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2733),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2736),
.A2(n_2577),
.B1(n_2610),
.B2(n_2605),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2739),
.B(n_2711),
.C(n_2720),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2766),
.B(n_2714),
.Y(n_2795)
);

AOI31xp33_ASAP7_75t_SL g2796 ( 
.A1(n_2782),
.A2(n_2723),
.A3(n_2727),
.B(n_2740),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2780),
.Y(n_2797)
);

AOI211x1_ASAP7_75t_SL g2798 ( 
.A1(n_2761),
.A2(n_2718),
.B(n_2715),
.C(n_2706),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2759),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2773),
.B(n_2710),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2764),
.Y(n_2801)
);

OAI21xp33_ASAP7_75t_L g2802 ( 
.A1(n_2758),
.A2(n_2767),
.B(n_2775),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2761),
.B(n_2745),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2778),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2770),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2769),
.B(n_2748),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2765),
.B(n_2703),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2757),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2776),
.B(n_2756),
.Y(n_2809)
);

NOR4xp25_ASAP7_75t_SL g2810 ( 
.A(n_2791),
.B(n_2698),
.C(n_2604),
.D(n_2614),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2768),
.B(n_2750),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2774),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2760),
.Y(n_2813)
);

INVxp67_ASAP7_75t_L g2814 ( 
.A(n_2781),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2784),
.B(n_2606),
.Y(n_2815)
);

OAI21xp5_ASAP7_75t_SL g2816 ( 
.A1(n_2758),
.A2(n_2777),
.B(n_2772),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2793),
.Y(n_2817)
);

OAI21xp33_ASAP7_75t_L g2818 ( 
.A1(n_2777),
.A2(n_2610),
.B(n_2619),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2779),
.B(n_2605),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2789),
.B(n_2651),
.Y(n_2820)
);

AOI22xp33_ASAP7_75t_SL g2821 ( 
.A1(n_2786),
.A2(n_2639),
.B1(n_2626),
.B2(n_2597),
.Y(n_2821)
);

OA211x2_ASAP7_75t_L g2822 ( 
.A1(n_2783),
.A2(n_2771),
.B(n_2794),
.C(n_2762),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2785),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2790),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2792),
.Y(n_2825)
);

OAI322xp33_ASAP7_75t_L g2826 ( 
.A1(n_2786),
.A2(n_2651),
.A3(n_2657),
.B1(n_2653),
.B2(n_2652),
.C1(n_2632),
.C2(n_2620),
.Y(n_2826)
);

AOI222xp33_ASAP7_75t_L g2827 ( 
.A1(n_2802),
.A2(n_2787),
.B1(n_2763),
.B2(n_2628),
.C1(n_2633),
.C2(n_2635),
.Y(n_2827)
);

AOI222xp33_ASAP7_75t_L g2828 ( 
.A1(n_2816),
.A2(n_2811),
.B1(n_2809),
.B2(n_2823),
.C1(n_2803),
.C2(n_2814),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2810),
.A2(n_2788),
.B(n_2653),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2797),
.B(n_2612),
.Y(n_2830)
);

NAND3xp33_ASAP7_75t_L g2831 ( 
.A(n_2821),
.B(n_2809),
.C(n_2795),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2797),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2818),
.B(n_2597),
.Y(n_2833)
);

OAI21xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2803),
.A2(n_2684),
.B(n_2645),
.Y(n_2834)
);

INVx1_ASAP7_75t_SL g2835 ( 
.A(n_2819),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2804),
.Y(n_2836)
);

OR2x2_ASAP7_75t_L g2837 ( 
.A(n_2800),
.B(n_2629),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2798),
.B(n_2619),
.Y(n_2838)
);

NAND4xp25_ASAP7_75t_L g2839 ( 
.A(n_2822),
.B(n_2657),
.C(n_2652),
.D(n_2594),
.Y(n_2839)
);

NAND3xp33_ASAP7_75t_L g2840 ( 
.A(n_2812),
.B(n_2600),
.C(n_2594),
.Y(n_2840)
);

INVxp67_ASAP7_75t_L g2841 ( 
.A(n_2807),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2807),
.Y(n_2842)
);

OAI221xp5_ASAP7_75t_L g2843 ( 
.A1(n_2796),
.A2(n_2406),
.B1(n_2600),
.B2(n_2621),
.C(n_2645),
.Y(n_2843)
);

OAI32xp33_ASAP7_75t_L g2844 ( 
.A1(n_2799),
.A2(n_2621),
.A3(n_2558),
.B1(n_2552),
.B2(n_2551),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2806),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2806),
.Y(n_2846)
);

OAI22x1_ASAP7_75t_L g2847 ( 
.A1(n_2813),
.A2(n_2638),
.B1(n_2644),
.B2(n_2617),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2820),
.Y(n_2848)
);

AOI21xp33_ASAP7_75t_SL g2849 ( 
.A1(n_2801),
.A2(n_2638),
.B(n_2617),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2815),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2808),
.Y(n_2851)
);

OAI322xp33_ASAP7_75t_L g2852 ( 
.A1(n_2838),
.A2(n_2817),
.A3(n_2805),
.B1(n_2824),
.B2(n_2820),
.C1(n_2825),
.C2(n_2826),
.Y(n_2852)
);

NOR2xp67_ASAP7_75t_L g2853 ( 
.A(n_2847),
.B(n_2638),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2830),
.B(n_2832),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2829),
.A2(n_2612),
.B(n_2644),
.Y(n_2855)
);

AOI221xp5_ASAP7_75t_L g2856 ( 
.A1(n_2834),
.A2(n_2644),
.B1(n_2558),
.B2(n_2552),
.C(n_2551),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2835),
.B(n_2562),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2843),
.B(n_2839),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2833),
.B(n_2485),
.Y(n_2859)
);

NAND3xp33_ASAP7_75t_L g2860 ( 
.A(n_2828),
.B(n_2529),
.C(n_2525),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2836),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2849),
.B(n_2485),
.Y(n_2862)
);

NOR3x1_ASAP7_75t_L g2863 ( 
.A(n_2831),
.B(n_2462),
.C(n_2525),
.Y(n_2863)
);

A2O1A1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2834),
.A2(n_2529),
.B(n_2339),
.C(n_2342),
.Y(n_2864)
);

BUFx2_ASAP7_75t_L g2865 ( 
.A(n_2841),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2827),
.A2(n_2339),
.B(n_2400),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2842),
.B(n_2369),
.Y(n_2867)
);

NOR3x1_ASAP7_75t_L g2868 ( 
.A(n_2840),
.B(n_2462),
.C(n_2286),
.Y(n_2868)
);

AOI31xp33_ASAP7_75t_L g2869 ( 
.A1(n_2850),
.A2(n_2414),
.A3(n_2434),
.B(n_2431),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2848),
.B(n_2845),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2855),
.A2(n_2846),
.B(n_2840),
.Y(n_2871)
);

O2A1O1Ixp33_ASAP7_75t_L g2872 ( 
.A1(n_2852),
.A2(n_2851),
.B(n_2837),
.C(n_2844),
.Y(n_2872)
);

OR2x2_ASAP7_75t_L g2873 ( 
.A(n_2854),
.B(n_2372),
.Y(n_2873)
);

NAND3xp33_ASAP7_75t_L g2874 ( 
.A(n_2858),
.B(n_2414),
.C(n_2382),
.Y(n_2874)
);

NAND4xp75_ASAP7_75t_L g2875 ( 
.A(n_2863),
.B(n_2438),
.C(n_2382),
.D(n_2393),
.Y(n_2875)
);

OAI221xp5_ASAP7_75t_SL g2876 ( 
.A1(n_2866),
.A2(n_2430),
.B1(n_2431),
.B2(n_2421),
.C(n_2393),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2857),
.B(n_2372),
.Y(n_2877)
);

NOR3xp33_ASAP7_75t_L g2878 ( 
.A(n_2865),
.B(n_2430),
.C(n_2402),
.Y(n_2878)
);

AOI32xp33_ASAP7_75t_L g2879 ( 
.A1(n_2862),
.A2(n_2859),
.A3(n_2861),
.B1(n_2856),
.B2(n_2870),
.Y(n_2879)
);

OAI211xp5_ASAP7_75t_L g2880 ( 
.A1(n_2853),
.A2(n_2402),
.B(n_2410),
.C(n_2398),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2860),
.A2(n_2438),
.B1(n_2410),
.B2(n_2421),
.Y(n_2881)
);

OAI21xp33_ASAP7_75t_SL g2882 ( 
.A1(n_2869),
.A2(n_2398),
.B(n_2462),
.Y(n_2882)
);

OAI321xp33_ASAP7_75t_L g2883 ( 
.A1(n_2867),
.A2(n_2462),
.A3(n_2334),
.B1(n_2292),
.B2(n_2387),
.C(n_2337),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2873),
.Y(n_2884)
);

AND4x1_ASAP7_75t_L g2885 ( 
.A(n_2871),
.B(n_2868),
.C(n_2864),
.D(n_111),
.Y(n_2885)
);

O2A1O1Ixp33_ASAP7_75t_L g2886 ( 
.A1(n_2872),
.A2(n_112),
.B(n_106),
.C(n_110),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2882),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2877),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2878),
.Y(n_2889)
);

OAI22x1_ASAP7_75t_L g2890 ( 
.A1(n_2874),
.A2(n_2456),
.B1(n_2344),
.B2(n_2338),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2876),
.Y(n_2891)
);

OAI22x1_ASAP7_75t_L g2892 ( 
.A1(n_2879),
.A2(n_2456),
.B1(n_2344),
.B2(n_115),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2880),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2875),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2883),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2881),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_SL g2897 ( 
.A(n_2885),
.B(n_2334),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2891),
.Y(n_2898)
);

OAI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2886),
.A2(n_2456),
.B(n_110),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2885),
.B(n_113),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2893),
.B(n_2887),
.Y(n_2901)
);

NOR3xp33_ASAP7_75t_L g2902 ( 
.A(n_2888),
.B(n_113),
.C(n_115),
.Y(n_2902)
);

OAI211xp5_ASAP7_75t_L g2903 ( 
.A1(n_2894),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2895),
.A2(n_2272),
.B1(n_2251),
.B2(n_122),
.Y(n_2904)
);

OAI221xp5_ASAP7_75t_SL g2905 ( 
.A1(n_2896),
.A2(n_117),
.B1(n_121),
.B2(n_124),
.C(n_125),
.Y(n_2905)
);

AOI221xp5_ASAP7_75t_L g2906 ( 
.A1(n_2889),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.C(n_128),
.Y(n_2906)
);

NAND4xp75_ASAP7_75t_L g2907 ( 
.A(n_2884),
.B(n_2892),
.C(n_2890),
.D(n_130),
.Y(n_2907)
);

NOR3xp33_ASAP7_75t_L g2908 ( 
.A(n_2886),
.B(n_128),
.C(n_129),
.Y(n_2908)
);

NAND3xp33_ASAP7_75t_SL g2909 ( 
.A(n_2885),
.B(n_129),
.C(n_131),
.Y(n_2909)
);

AOI211xp5_ASAP7_75t_L g2910 ( 
.A1(n_2886),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_2889),
.B(n_132),
.Y(n_2911)
);

NAND5xp2_ASAP7_75t_L g2912 ( 
.A(n_2886),
.B(n_134),
.C(n_135),
.D(n_136),
.E(n_138),
.Y(n_2912)
);

AOI221xp5_ASAP7_75t_L g2913 ( 
.A1(n_2886),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.C(n_140),
.Y(n_2913)
);

AOI32xp33_ASAP7_75t_L g2914 ( 
.A1(n_2900),
.A2(n_139),
.A3(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_2914)
);

NOR4xp75_ASAP7_75t_L g2915 ( 
.A(n_2901),
.B(n_145),
.C(n_142),
.D(n_144),
.Y(n_2915)
);

AOI211xp5_ASAP7_75t_L g2916 ( 
.A1(n_2909),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2916)
);

OAI222xp33_ASAP7_75t_L g2917 ( 
.A1(n_2898),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.C1(n_152),
.C2(n_155),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2907),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2902),
.B(n_2251),
.Y(n_2919)
);

NAND4xp25_ASAP7_75t_L g2920 ( 
.A(n_2908),
.B(n_2910),
.C(n_2912),
.D(n_2897),
.Y(n_2920)
);

AOI222xp33_ASAP7_75t_L g2921 ( 
.A1(n_2899),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.C1(n_156),
.C2(n_158),
.Y(n_2921)
);

AOI31xp33_ASAP7_75t_L g2922 ( 
.A1(n_2913),
.A2(n_164),
.A3(n_160),
.B(n_162),
.Y(n_2922)
);

AOI221xp5_ASAP7_75t_L g2923 ( 
.A1(n_2905),
.A2(n_160),
.B1(n_162),
.B2(n_165),
.C(n_167),
.Y(n_2923)
);

OAI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2911),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2906),
.B(n_2903),
.Y(n_2925)
);

O2A1O1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2904),
.A2(n_168),
.B(n_169),
.C(n_173),
.Y(n_2926)
);

O2A1O1Ixp33_ASAP7_75t_SL g2927 ( 
.A1(n_2909),
.A2(n_176),
.B(n_177),
.C(n_181),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2908),
.B(n_176),
.Y(n_2928)
);

AOI221xp5_ASAP7_75t_SL g2929 ( 
.A1(n_2920),
.A2(n_177),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2922),
.B(n_182),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2927),
.B(n_184),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2915),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2924),
.Y(n_2933)
);

OAI211xp5_ASAP7_75t_SL g2934 ( 
.A1(n_2918),
.A2(n_185),
.B(n_186),
.C(n_188),
.Y(n_2934)
);

O2A1O1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_2925),
.A2(n_185),
.B(n_186),
.C(n_188),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2928),
.B(n_2272),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2928),
.Y(n_2937)
);

OAI211xp5_ASAP7_75t_L g2938 ( 
.A1(n_2921),
.A2(n_189),
.B(n_190),
.C(n_191),
.Y(n_2938)
);

OR2x2_ASAP7_75t_L g2939 ( 
.A(n_2919),
.B(n_191),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2914),
.B(n_192),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2929),
.B(n_2916),
.Y(n_2941)
);

NAND4xp75_ASAP7_75t_L g2942 ( 
.A(n_2940),
.B(n_2923),
.C(n_2926),
.D(n_2917),
.Y(n_2942)
);

AOI22x1_ASAP7_75t_SL g2943 ( 
.A1(n_2932),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_2943)
);

OAI211xp5_ASAP7_75t_L g2944 ( 
.A1(n_2938),
.A2(n_195),
.B(n_1281),
.C(n_1282),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2931),
.Y(n_2945)
);

NAND4xp75_ASAP7_75t_L g2946 ( 
.A(n_2930),
.B(n_2937),
.C(n_2936),
.D(n_2933),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2939),
.Y(n_2947)
);

O2A1O1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2935),
.A2(n_1282),
.B(n_200),
.C(n_201),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2934),
.Y(n_2949)
);

NAND4xp75_ASAP7_75t_L g2950 ( 
.A(n_2929),
.B(n_198),
.C(n_203),
.D(n_209),
.Y(n_2950)
);

OAI211xp5_ASAP7_75t_L g2951 ( 
.A1(n_2938),
.A2(n_210),
.B(n_225),
.C(n_226),
.Y(n_2951)
);

OAI211xp5_ASAP7_75t_SL g2952 ( 
.A1(n_2949),
.A2(n_870),
.B(n_857),
.C(n_233),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2942),
.A2(n_2941),
.B1(n_2945),
.B2(n_2946),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2950),
.B(n_227),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2947),
.B(n_228),
.Y(n_2955)
);

NOR3xp33_ASAP7_75t_L g2956 ( 
.A(n_2951),
.B(n_870),
.C(n_857),
.Y(n_2956)
);

NAND3xp33_ASAP7_75t_SL g2957 ( 
.A(n_2944),
.B(n_2948),
.C(n_2943),
.Y(n_2957)
);

OAI221xp5_ASAP7_75t_SL g2958 ( 
.A1(n_2949),
.A2(n_234),
.B1(n_242),
.B2(n_245),
.C(n_246),
.Y(n_2958)
);

NAND3xp33_ASAP7_75t_SL g2959 ( 
.A(n_2951),
.B(n_247),
.C(n_248),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2949),
.B(n_250),
.Y(n_2960)
);

OAI211xp5_ASAP7_75t_SL g2961 ( 
.A1(n_2949),
.A2(n_258),
.B(n_259),
.C(n_260),
.Y(n_2961)
);

NOR3xp33_ASAP7_75t_SL g2962 ( 
.A(n_2946),
.B(n_261),
.C(n_269),
.Y(n_2962)
);

AOI221xp5_ASAP7_75t_L g2963 ( 
.A1(n_2949),
.A2(n_880),
.B1(n_887),
.B2(n_874),
.C(n_877),
.Y(n_2963)
);

NOR3xp33_ASAP7_75t_L g2964 ( 
.A(n_2946),
.B(n_858),
.C(n_273),
.Y(n_2964)
);

XNOR2xp5_ASAP7_75t_L g2965 ( 
.A(n_2953),
.B(n_274),
.Y(n_2965)
);

OR3x1_ASAP7_75t_L g2966 ( 
.A(n_2957),
.B(n_2959),
.C(n_2961),
.Y(n_2966)
);

XNOR2xp5_ASAP7_75t_L g2967 ( 
.A(n_2962),
.B(n_275),
.Y(n_2967)
);

XNOR2x1_ASAP7_75t_L g2968 ( 
.A(n_2954),
.B(n_281),
.Y(n_2968)
);

AND2x4_ASAP7_75t_L g2969 ( 
.A(n_2960),
.B(n_282),
.Y(n_2969)
);

AND4x1_ASAP7_75t_L g2970 ( 
.A(n_2964),
.B(n_283),
.C(n_286),
.D(n_288),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2955),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2958),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2967),
.Y(n_2973)
);

CKINVDCx20_ASAP7_75t_R g2974 ( 
.A(n_2965),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2968),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2969),
.Y(n_2976)
);

AOI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2966),
.A2(n_2952),
.B1(n_2956),
.B2(n_2963),
.Y(n_2977)
);

AOI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2972),
.A2(n_1251),
.B1(n_1232),
.B2(n_1195),
.Y(n_2978)
);

AOI211xp5_ASAP7_75t_SL g2979 ( 
.A1(n_2971),
.A2(n_289),
.B(n_290),
.C(n_295),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2970),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2967),
.Y(n_2981)
);

AO22x2_ASAP7_75t_L g2982 ( 
.A1(n_2968),
.A2(n_1291),
.B1(n_299),
.B2(n_302),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2966),
.A2(n_1232),
.B1(n_1251),
.B2(n_1195),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2966),
.A2(n_1232),
.B1(n_1251),
.B2(n_1195),
.Y(n_2984)
);

OAI22x1_ASAP7_75t_L g2985 ( 
.A1(n_2967),
.A2(n_298),
.B1(n_305),
.B2(n_310),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2967),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2967),
.Y(n_2987)
);

OAI22x1_ASAP7_75t_L g2988 ( 
.A1(n_2967),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2988)
);

AOI31xp33_ASAP7_75t_L g2989 ( 
.A1(n_2965),
.A2(n_314),
.A3(n_321),
.B(n_322),
.Y(n_2989)
);

HB1xp67_ASAP7_75t_L g2990 ( 
.A(n_2967),
.Y(n_2990)
);

OAI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2974),
.A2(n_1335),
.B1(n_1333),
.B2(n_875),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2980),
.A2(n_875),
.B1(n_887),
.B2(n_877),
.Y(n_2992)
);

AOI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2985),
.A2(n_1232),
.B1(n_1251),
.B2(n_1195),
.Y(n_2993)
);

HB1xp67_ASAP7_75t_L g2994 ( 
.A(n_2988),
.Y(n_2994)
);

INVx2_ASAP7_75t_SL g2995 ( 
.A(n_2982),
.Y(n_2995)
);

AOI31xp33_ASAP7_75t_L g2996 ( 
.A1(n_2975),
.A2(n_323),
.A3(n_326),
.B(n_327),
.Y(n_2996)
);

AOI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2973),
.A2(n_1195),
.B1(n_1291),
.B2(n_953),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2976),
.Y(n_2998)
);

OAI31xp33_ASAP7_75t_L g2999 ( 
.A1(n_2982),
.A2(n_2987),
.A3(n_2981),
.B(n_2990),
.Y(n_2999)
);

HB1xp67_ASAP7_75t_L g3000 ( 
.A(n_2986),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2977),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2989),
.Y(n_3002)
);

INVx1_ASAP7_75t_SL g3003 ( 
.A(n_2978),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2979),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2983),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2984),
.A2(n_953),
.B1(n_887),
.B2(n_874),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2980),
.B(n_328),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2980),
.Y(n_3008)
);

AND2x2_ASAP7_75t_SL g3009 ( 
.A(n_2980),
.B(n_874),
.Y(n_3009)
);

AOI31xp33_ASAP7_75t_L g3010 ( 
.A1(n_2980),
.A2(n_334),
.A3(n_335),
.B(n_338),
.Y(n_3010)
);

AOI22xp5_ASAP7_75t_L g3011 ( 
.A1(n_2974),
.A2(n_953),
.B1(n_887),
.B2(n_874),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2980),
.B(n_341),
.Y(n_3012)
);

AOI31xp33_ASAP7_75t_L g3013 ( 
.A1(n_2980),
.A2(n_344),
.A3(n_345),
.B(n_350),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2982),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2974),
.A2(n_953),
.B1(n_874),
.B2(n_880),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2982),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2980),
.B(n_355),
.Y(n_3017)
);

AOI222xp33_ASAP7_75t_L g3018 ( 
.A1(n_2998),
.A2(n_880),
.B1(n_877),
.B2(n_875),
.C1(n_366),
.C2(n_368),
.Y(n_3018)
);

OR5x1_ASAP7_75t_L g3019 ( 
.A(n_2999),
.B(n_358),
.C(n_359),
.D(n_360),
.E(n_369),
.Y(n_3019)
);

NAND3xp33_ASAP7_75t_L g3020 ( 
.A(n_3000),
.B(n_880),
.C(n_877),
.Y(n_3020)
);

OAI22xp5_ASAP7_75t_SL g3021 ( 
.A1(n_2995),
.A2(n_373),
.B1(n_377),
.B2(n_378),
.Y(n_3021)
);

OAI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_3008),
.A2(n_875),
.B1(n_1208),
.B2(n_1323),
.Y(n_3022)
);

NOR2x1p5_ASAP7_75t_L g3023 ( 
.A(n_3007),
.B(n_381),
.Y(n_3023)
);

OR5x1_ASAP7_75t_L g3024 ( 
.A(n_3014),
.B(n_383),
.C(n_386),
.D(n_388),
.E(n_389),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_3017),
.A2(n_1254),
.B1(n_1331),
.B2(n_1231),
.Y(n_3025)
);

AO22x1_ASAP7_75t_L g3026 ( 
.A1(n_3002),
.A2(n_390),
.B1(n_393),
.B2(n_394),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_SL g3027 ( 
.A1(n_3004),
.A2(n_2994),
.B1(n_3001),
.B2(n_3012),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_3016),
.A2(n_3005),
.B1(n_3003),
.B2(n_3009),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2993),
.A2(n_1303),
.B1(n_1331),
.B2(n_1254),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_2991),
.A2(n_1303),
.B1(n_1331),
.B2(n_1254),
.Y(n_3030)
);

AOI221xp5_ASAP7_75t_L g3031 ( 
.A1(n_2992),
.A2(n_1303),
.B1(n_858),
.B2(n_1026),
.C(n_1024),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_3006),
.A2(n_1030),
.B1(n_1026),
.B2(n_1025),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_3011),
.A2(n_1030),
.B1(n_1025),
.B2(n_1024),
.Y(n_3033)
);

O2A1O1Ixp33_ASAP7_75t_L g3034 ( 
.A1(n_2996),
.A2(n_397),
.B(n_398),
.C(n_402),
.Y(n_3034)
);

NOR4xp25_ASAP7_75t_L g3035 ( 
.A(n_3010),
.B(n_3013),
.C(n_3015),
.D(n_2997),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_SL g3036 ( 
.A1(n_2995),
.A2(n_407),
.B1(n_1158),
.B2(n_1224),
.Y(n_3036)
);

AOI221xp5_ASAP7_75t_L g3037 ( 
.A1(n_3008),
.A2(n_1293),
.B1(n_1300),
.B2(n_1276),
.C(n_1265),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_SL g3038 ( 
.A1(n_2995),
.A2(n_1158),
.B1(n_1224),
.B2(n_1170),
.Y(n_3038)
);

OR5x1_ASAP7_75t_L g3039 ( 
.A(n_2999),
.B(n_1308),
.C(n_1312),
.D(n_1320),
.E(n_1323),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_3017),
.B(n_1111),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_SL g3041 ( 
.A1(n_2995),
.A2(n_1158),
.B1(n_1224),
.B2(n_1170),
.Y(n_3041)
);

AOI31xp33_ASAP7_75t_L g3042 ( 
.A1(n_3027),
.A2(n_1050),
.A3(n_1125),
.B(n_1120),
.Y(n_3042)
);

OAI22xp33_ASAP7_75t_SL g3043 ( 
.A1(n_3040),
.A2(n_1409),
.B1(n_1353),
.B2(n_1276),
.Y(n_3043)
);

AOI31xp33_ASAP7_75t_L g3044 ( 
.A1(n_3028),
.A2(n_1095),
.A3(n_1133),
.B(n_1125),
.Y(n_3044)
);

AOI31xp33_ASAP7_75t_L g3045 ( 
.A1(n_3020),
.A2(n_1089),
.A3(n_1119),
.B(n_1111),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_3036),
.A2(n_1089),
.B1(n_1050),
.B2(n_1120),
.Y(n_3046)
);

AOI31xp33_ASAP7_75t_L g3047 ( 
.A1(n_3019),
.A2(n_1088),
.A3(n_1119),
.B(n_1097),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_3018),
.A2(n_1088),
.B1(n_1039),
.B2(n_1097),
.Y(n_3048)
);

AOI31xp33_ASAP7_75t_L g3049 ( 
.A1(n_3031),
.A2(n_1087),
.A3(n_1042),
.B(n_1095),
.Y(n_3049)
);

AOI31xp33_ASAP7_75t_L g3050 ( 
.A1(n_3022),
.A2(n_1087),
.A3(n_1042),
.B(n_1045),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_3038),
.A2(n_1061),
.B1(n_1086),
.B2(n_1067),
.Y(n_3051)
);

AOI31xp33_ASAP7_75t_L g3052 ( 
.A1(n_3024),
.A2(n_1062),
.A3(n_1061),
.B(n_1086),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_3041),
.A2(n_1062),
.B1(n_1067),
.B2(n_1045),
.Y(n_3053)
);

OAI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_3023),
.A2(n_1208),
.B1(n_1323),
.B2(n_1320),
.Y(n_3054)
);

AOI31xp33_ASAP7_75t_L g3055 ( 
.A1(n_3029),
.A2(n_1048),
.A3(n_1308),
.B(n_1312),
.Y(n_3055)
);

AOI31xp33_ASAP7_75t_L g3056 ( 
.A1(n_3032),
.A2(n_1077),
.A3(n_1101),
.B(n_1005),
.Y(n_3056)
);

OAI221xp5_ASAP7_75t_L g3057 ( 
.A1(n_3046),
.A2(n_3034),
.B1(n_3025),
.B2(n_3030),
.C(n_3035),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_SL g3058 ( 
.A1(n_3054),
.A2(n_3039),
.B1(n_3021),
.B2(n_3033),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_3047),
.B(n_3037),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3042),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3044),
.Y(n_3061)
);

CKINVDCx20_ASAP7_75t_R g3062 ( 
.A(n_3052),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_3048),
.Y(n_3063)
);

NAND5xp2_ASAP7_75t_L g3064 ( 
.A(n_3051),
.B(n_3026),
.C(n_1158),
.D(n_1287),
.E(n_1242),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_3045),
.Y(n_3065)
);

BUFx3_ASAP7_75t_L g3066 ( 
.A(n_3049),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_3050),
.A2(n_1077),
.B(n_1101),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_3058),
.Y(n_3068)
);

AOI21xp33_ASAP7_75t_SL g3069 ( 
.A1(n_3057),
.A2(n_3056),
.B(n_3055),
.Y(n_3069)
);

OA21x2_ASAP7_75t_L g3070 ( 
.A1(n_3059),
.A2(n_3053),
.B(n_3043),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3062),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_3065),
.A2(n_1028),
.B(n_1011),
.Y(n_3072)
);

NAND3xp33_ASAP7_75t_L g3073 ( 
.A(n_3063),
.B(n_994),
.C(n_1021),
.Y(n_3073)
);

OAI31xp33_ASAP7_75t_L g3074 ( 
.A1(n_3064),
.A2(n_1225),
.A3(n_1253),
.B(n_988),
.Y(n_3074)
);

OR2x6_ASAP7_75t_L g3075 ( 
.A(n_3060),
.B(n_1017),
.Y(n_3075)
);

NAND3xp33_ASAP7_75t_L g3076 ( 
.A(n_3068),
.B(n_3061),
.C(n_3066),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_3071),
.B(n_3067),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_3074),
.B(n_1011),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_3078),
.Y(n_3079)
);

XNOR2xp5_ASAP7_75t_L g3080 ( 
.A(n_3079),
.B(n_3076),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_L g3081 ( 
.A1(n_3080),
.A2(n_3077),
.B1(n_3075),
.B2(n_3070),
.Y(n_3081)
);

AOI211xp5_ASAP7_75t_L g3082 ( 
.A1(n_3081),
.A2(n_3069),
.B(n_3072),
.C(n_3073),
.Y(n_3082)
);


endmodule