module real_jpeg_4162_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_286;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_228;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_1),
.B(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_3),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_4),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_5),
.Y(n_225)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_7),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_7),
.B(n_188),
.Y(n_187)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_9),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_9),
.B(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_11),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_12),
.B(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_14),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_14),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_14),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_14),
.B(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_179),
.B1(n_180),
.B2(n_292),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_18),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_177),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_150),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_20),
.B(n_150),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.C(n_57),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_23),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_37),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_26),
.B(n_31),
.C(n_38),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_27),
.B(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_29),
.Y(n_146)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_30),
.Y(n_239)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_35),
.Y(n_148)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_43),
.A2(n_57),
.B1(n_58),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_51),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_44),
.A2(n_51),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_44),
.Y(n_158)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_47),
.B(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_50),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_51),
.Y(n_159)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_55),
.Y(n_171)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_56),
.Y(n_209)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_59),
.Y(n_173)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_62),
.Y(n_249)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_82),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_76),
.B(n_122),
.Y(n_198)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_78),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_82),
.Y(n_294)
);

FAx1_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.CI(n_95),
.CON(n_82),
.SN(n_82)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_84),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_136),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_117),
.C(n_119),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_117),
.B1(n_118),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_106),
.C(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_103),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_103),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_116),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_114),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_131),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_120),
.A2(n_121),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_284)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_174),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_151),
.A2(n_152),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_155),
.B(n_174),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_172),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_156),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_160),
.B(n_172),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_168),
.B(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_286),
.B(n_291),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_273),
.B(n_285),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_231),
.B(n_272),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_216),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_184),
.B(n_216),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_199),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_200),
.C(n_213),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_186),
.B(n_194),
.C(n_198),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_189),
.B1(n_190),
.B2(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_213),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.C(n_210),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_229),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_220),
.B1(n_229),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_266),
.B(n_271),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_253),
.B(n_265),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_244),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_243),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_240),
.C(n_243),
.Y(n_267)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_261),
.B(n_264),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_281),
.C(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);


endmodule