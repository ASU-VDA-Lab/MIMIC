module fake_jpeg_8302_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx2_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_43),
.Y(n_52)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_31),
.B1(n_22),
.B2(n_43),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_56),
.B1(n_59),
.B2(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_38),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_63),
.B1(n_17),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_68),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_34),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_81),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_89),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_37),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_39),
.C(n_61),
.Y(n_123)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_128)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_41),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_39),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_48),
.B1(n_38),
.B2(n_40),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_122),
.B1(n_127),
.B2(n_101),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_70),
.B(n_80),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_36),
.B(n_39),
.C(n_46),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_48),
.B1(n_40),
.B2(n_37),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_66),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_48),
.B1(n_40),
.B2(n_41),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_88),
.B1(n_82),
.B2(n_89),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_76),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_39),
.C(n_41),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_98),
.C(n_25),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_135),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_140),
.B(n_143),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_150),
.C(n_104),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_74),
.Y(n_136)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_114),
.B1(n_112),
.B2(n_115),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_41),
.B(n_93),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_111),
.B(n_73),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_142),
.B1(n_144),
.B2(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_32),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_86),
.B1(n_84),
.B2(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_32),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_30),
.Y(n_145)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_0),
.Y(n_147)
);

NAND2x1p5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_1),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_158),
.B(n_160),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_27),
.B1(n_26),
.B2(n_3),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_108),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_111),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_27),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_85),
.B(n_83),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_167),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_129),
.B(n_107),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_165),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_109),
.A3(n_120),
.B1(n_108),
.B2(n_128),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_173),
.B(n_177),
.Y(n_212)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_107),
.C(n_114),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_150),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_192),
.B1(n_153),
.B2(n_139),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_112),
.B(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_186),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_26),
.C(n_27),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_178),
.B(n_182),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_184),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_160),
.B1(n_137),
.B2(n_131),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_156),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_26),
.B(n_9),
.C(n_15),
.D(n_4),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_9),
.C(n_15),
.Y(n_187)
);

BUFx12f_ASAP7_75t_SL g215 ( 
.A(n_187),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_111),
.B1(n_2),
.B2(n_3),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_146),
.B1(n_144),
.B2(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_202),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_199),
.B(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_205),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_214),
.B1(n_216),
.B2(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_226),
.C(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_163),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_197),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_163),
.CI(n_161),
.CON(n_223),
.SN(n_223)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_134),
.C(n_191),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_168),
.B1(n_166),
.B2(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_238),
.B1(n_207),
.B2(n_211),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_168),
.B1(n_170),
.B2(n_162),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_189),
.B1(n_162),
.B2(n_143),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_212),
.B(n_185),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_191),
.C(n_158),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_210),
.C(n_205),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_252),
.B1(n_224),
.B2(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_247),
.Y(n_270)
);

AOI211xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_224),
.B(n_235),
.C(n_177),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_203),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_258),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_250),
.C(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_214),
.C(n_217),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_195),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_149),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_200),
.B1(n_215),
.B2(n_140),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_220),
.C(n_237),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_265),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_233),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_266),
.B1(n_242),
.B2(n_256),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_242),
.B(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_226),
.B1(n_223),
.B2(n_236),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_253),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_223),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_251),
.B(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_202),
.C(n_147),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_4),
.B(n_5),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_278),
.B(n_281),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_254),
.CI(n_243),
.CON(n_274),
.SN(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_283),
.B1(n_5),
.B2(n_7),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_244),
.B1(n_215),
.B2(n_138),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_138),
.B1(n_186),
.B2(n_8),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_138),
.B(n_8),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_5),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_286),
.B(n_288),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_269),
.B(n_262),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.C(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_7),
.C(n_8),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_277),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_280),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_274),
.B1(n_278),
.B2(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_10),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_12),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_299),
.B(n_12),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_287),
.A2(n_282),
.B(n_11),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_10),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_10),
.A3(n_12),
.B1(n_14),
.B2(n_293),
.C1(n_297),
.C2(n_298),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_302),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_14),
.Y(n_309)
);


endmodule