module fake_jpeg_665_n_222 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_1),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_66),
.B1(n_60),
.B2(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_91),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_62),
.C(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_66),
.B1(n_60),
.B2(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_63),
.B1(n_68),
.B2(n_55),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_68),
.B1(n_73),
.B2(n_61),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_97),
.B1(n_67),
.B2(n_55),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_54),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_119),
.Y(n_135)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_72),
.B1(n_77),
.B2(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_78),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_73),
.B1(n_85),
.B2(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_69),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_126),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_93),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_40),
.C(n_39),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_95),
.B1(n_93),
.B2(n_59),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_111),
.B1(n_102),
.B2(n_56),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_129),
.C(n_2),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_118),
.C(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_93),
.B1(n_57),
.B2(n_72),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_140),
.B1(n_141),
.B2(n_43),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_138),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_77),
.B(n_71),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_3),
.B(n_4),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_57),
.B1(n_72),
.B2(n_59),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_157),
.B(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_111),
.B1(n_56),
.B2(n_4),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_52),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_6),
.C(n_9),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_124),
.B1(n_122),
.B2(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_2),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_154),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_127),
.B1(n_139),
.B2(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_160),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_42),
.C(n_41),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_3),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_5),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_165),
.B(n_10),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_171),
.Y(n_191)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_179),
.Y(n_194)
);

OAI322xp33_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_176),
.A3(n_172),
.B1(n_181),
.B2(n_178),
.C1(n_21),
.C2(n_22),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_12),
.B(n_16),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_38),
.B(n_37),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_29),
.B(n_28),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_35),
.C(n_34),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_162),
.C(n_166),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_145),
.B1(n_165),
.B2(n_148),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_17),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_160),
.B1(n_31),
.B2(n_30),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_180),
.B1(n_168),
.B2(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_175),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_173),
.B1(n_19),
.B2(n_20),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_182),
.B(n_170),
.Y(n_197)
);

AND3x1_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_189),
.C(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_177),
.C(n_169),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

OA21x2_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_27),
.B(n_18),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_173),
.C(n_18),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_195),
.B1(n_188),
.B2(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_211),
.B1(n_198),
.B2(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_199),
.C(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_203),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_208),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_216),
.C(n_210),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_19),
.B(n_20),
.Y(n_220)
);

OAI211xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_24),
.Y(n_222)
);


endmodule