module real_jpeg_32851_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_12),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_1),
.Y(n_36)
);

CKINVDCx11_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx2_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2x1p5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_22),
.Y(n_31)
);

AOI221xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.C(n_49),
.Y(n_42)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AND2x4_ASAP7_75t_SL g46 ( 
.A(n_4),
.B(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_7),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_30),
.Y(n_29)
);

OAI211xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_15),
.B(n_25),
.C(n_42),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_27),
.B1(n_34),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

AND2x4_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_13),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_14),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_28),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_28),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_29),
.B(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI221xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.C(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);


endmodule