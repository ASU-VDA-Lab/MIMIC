module real_jpeg_13595_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_249, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_249;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_54),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_4),
.A2(n_36),
.B1(n_38),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_4),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_29),
.C(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_62),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_98),
.B(n_154),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_50),
.B(n_63),
.C(n_181),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_36),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_45),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_8),
.A2(n_36),
.B1(n_38),
.B2(n_68),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_68),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_36),
.B1(n_38),
.B2(n_57),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_57),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_12),
.B(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_25),
.B1(n_29),
.B2(n_59),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_36),
.B1(n_38),
.B2(n_59),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_15),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_15),
.A2(n_30),
.B1(n_36),
.B2(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_25),
.B1(n_29),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_103),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.C(n_60),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_22),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_23),
.B(n_33),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_24),
.A2(n_27),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_24),
.A2(n_27),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_24),
.B(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_25),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_25),
.B(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_27),
.B(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_31),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_36),
.B(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_38),
.A2(n_64),
.B(n_139),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_39),
.A2(n_46),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_39),
.A2(n_44),
.B1(n_46),
.B2(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_39),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_39),
.B(n_141),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_39),
.A2(n_46),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_43),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_43),
.B(n_139),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_43),
.A2(n_151),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_46),
.B(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_58),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_48),
.A2(n_55),
.B(n_139),
.C(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_56),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_49),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_50),
.A2(n_52),
.A3(n_55),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_66),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_65),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_61),
.A2(n_66),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_61),
.A2(n_89),
.B1(n_116),
.B2(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_67),
.Y(n_117)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_84),
.B2(n_85),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_83),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_95),
.B2(n_102),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_89),
.A2(n_117),
.B(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_93),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_99),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_98),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_98),
.A2(n_99),
.B1(n_124),
.B2(n_183),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_99),
.A2(n_160),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_139),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_99),
.A2(n_168),
.B(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_108),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_104),
.B(n_106),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_108),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_118),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_236)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_232),
.A3(n_241),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_214),
.B(n_231),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_193),
.B(n_213),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_176),
.B(n_192),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_156),
.B(n_175),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_137),
.A2(n_140),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_164),
.B(n_174),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_158),
.B(n_162),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B(n_173),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_177),
.B(n_178),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_187),
.C(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_182),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_206),
.B2(n_207),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_209),
.C(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_201),
.C(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_216),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_228),
.C(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_226),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_223),
.C(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_235),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);


endmodule