module fake_jpeg_7249_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_57),
.B1(n_64),
.B2(n_66),
.Y(n_90)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_75),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_64),
.B1(n_18),
.B2(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_72),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_19),
.B(n_30),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_76),
.B(n_96),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_73),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_30),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_47),
.C(n_37),
.Y(n_117)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_81),
.Y(n_127)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_18),
.B(n_31),
.C(n_34),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_95),
.B1(n_37),
.B2(n_35),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_16),
.B1(n_44),
.B2(n_43),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_22),
.B1(n_29),
.B2(n_34),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_102),
.B1(n_59),
.B2(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_130),
.B1(n_91),
.B2(n_69),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_31),
.B(n_34),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_88),
.B(n_26),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_47),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_1),
.Y(n_142)
);

AO21x1_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_82),
.B(n_72),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_35),
.B1(n_51),
.B2(n_59),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_51),
.B1(n_54),
.B2(n_25),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_67),
.A3(n_79),
.B1(n_81),
.B2(n_95),
.Y(n_122)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_44),
.B1(n_40),
.B2(n_43),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_51),
.B1(n_25),
.B2(n_40),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_94),
.B1(n_83),
.B2(n_77),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_25),
.B1(n_28),
.B2(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_102),
.B1(n_28),
.B2(n_26),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_143),
.B1(n_145),
.B2(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_138),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVxp33_ASAP7_75t_SL g172 ( 
.A(n_136),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_93),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_146),
.C(n_156),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_157),
.B(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_26),
.Y(n_192)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_91),
.B1(n_94),
.B2(n_82),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_44),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_160),
.Y(n_166)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_80),
.B1(n_85),
.B2(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_131),
.B1(n_130),
.B2(n_108),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_101),
.B1(n_28),
.B2(n_20),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_105),
.B1(n_109),
.B2(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_155),
.B(n_158),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_110),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_28),
.C(n_92),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_104),
.B(n_10),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_105),
.B1(n_124),
.B2(n_109),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_197),
.B(n_15),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_178),
.B1(n_182),
.B2(n_187),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_122),
.B1(n_108),
.B2(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_110),
.B1(n_106),
.B2(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_185),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_190),
.B1(n_193),
.B2(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_137),
.C(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_112),
.B1(n_128),
.B2(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_112),
.B1(n_128),
.B2(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_4),
.B(n_5),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_134),
.A2(n_129),
.B1(n_116),
.B2(n_28),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_135),
.A2(n_116),
.B1(n_28),
.B2(n_26),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_142),
.B(n_148),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_139),
.A2(n_28),
.B1(n_20),
.B2(n_26),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_1),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_142),
.A2(n_26),
.B1(n_15),
.B2(n_13),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_215),
.B1(n_197),
.B2(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_135),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_164),
.C(n_194),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_149),
.B(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_206),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_162),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_211),
.C(n_222),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_1),
.B(n_2),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_209),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_152),
.C(n_3),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_193),
.B1(n_170),
.B2(n_165),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_221),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_168),
.A2(n_2),
.B(n_3),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_192),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_2),
.C(n_4),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_175),
.C(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_4),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_244),
.B1(n_210),
.B2(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_200),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_179),
.B1(n_181),
.B2(n_169),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_242),
.B1(n_249),
.B2(n_251),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_170),
.C(n_188),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_246),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_180),
.B1(n_174),
.B2(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_223),
.B1(n_218),
.B2(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_165),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_167),
.B1(n_175),
.B2(n_6),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_204),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NOR2x1_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_224),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_12),
.B(n_10),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_227),
.B1(n_216),
.B2(n_201),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_262),
.B1(n_229),
.B2(n_235),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_227),
.B1(n_206),
.B2(n_220),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_211),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_269),
.C(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_251),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_226),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_226),
.C(n_6),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_228),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_242),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_285),
.Y(n_299)
);

AO221x1_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_234),
.B1(n_233),
.B2(n_236),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_261),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_267),
.C(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_288),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_233),
.C(n_8),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_269),
.C(n_254),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_11),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_297),
.C(n_303),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_257),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_253),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_293),
.B(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_280),
.B1(n_289),
.B2(n_282),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_273),
.B1(n_274),
.B2(n_7),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_276),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_281),
.C(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_313),
.C(n_11),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_280),
.C(n_284),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_273),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_315),
.B(n_314),
.C(n_7),
.Y(n_324)
);

HB1xp67_ASAP7_75t_SL g326 ( 
.A(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_321),
.Y(n_328)
);

AOI321xp33_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_329),
.A3(n_330),
.B1(n_304),
.B2(n_311),
.C(n_313),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_322),
.B(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_327),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_325),
.C(n_11),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_12),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_8),
.Y(n_335)
);


endmodule