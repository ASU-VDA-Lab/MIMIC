module fake_jpeg_20572_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

NAND2xp67_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_51),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_40),
.C(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_43),
.Y(n_86)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_55),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_82),
.C(n_4),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_86),
.C(n_37),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_45),
.B1(n_54),
.B2(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_84),
.B1(n_9),
.B2(n_11),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_41),
.C(n_47),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_56),
.B1(n_48),
.B2(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_42),
.B1(n_38),
.B2(n_3),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_2),
.Y(n_92)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_103),
.C(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_92),
.B1(n_95),
.B2(n_94),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_107),
.C(n_110),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_106),
.B1(n_94),
.B2(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_18),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_25),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_29),
.B(n_31),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_33),
.Y(n_118)
);


endmodule