module real_jpeg_20169_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_0),
.A2(n_30),
.B1(n_74),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_0),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_74),
.B1(n_79),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_97),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_97),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_97),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_74),
.B1(n_79),
.B2(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_27),
.B1(n_31),
.B2(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_151),
.Y(n_207)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_6),
.A2(n_74),
.B1(n_79),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_129),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_129),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_7),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_7),
.B(n_76),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_7),
.A2(n_14),
.B(n_35),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_60),
.B1(n_158),
.B2(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_7),
.B(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_7),
.B(n_47),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_7),
.A2(n_47),
.B(n_231),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_34),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_39),
.B1(n_74),
.B2(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_31),
.B(n_33),
.C(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_106),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_105),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_55),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_25),
.A2(n_41),
.B(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_26),
.Y(n_142)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_27),
.A2(n_36),
.B(n_149),
.C(n_198),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_27),
.B(n_45),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_31),
.A2(n_46),
.A3(n_48),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_33),
.A2(n_41),
.B1(n_66),
.B2(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_37),
.B(n_93),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_33),
.A2(n_41),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_33),
.B(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_33),
.A2(n_41),
.B1(n_202),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_33),
.A2(n_41),
.B1(n_222),
.B2(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_34),
.B(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_66),
.B(n_67),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_41),
.A2(n_67),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_43)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_44),
.A2(n_50),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_44),
.A2(n_50),
.B1(n_180),
.B2(n_235),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_47),
.B(n_73),
.Y(n_155)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_48),
.A2(n_75),
.B1(n_148),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_51),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_50),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_50),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_50),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_70),
.B1(n_82),
.B2(n_83),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_65),
.B1(n_83),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_63),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_60),
.A2(n_119),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_60),
.A2(n_62),
.B1(n_192),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_60),
.A2(n_90),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_61),
.A2(n_91),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_61),
.A2(n_64),
.B(n_121),
.Y(n_229)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_89),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_77),
.B(n_80),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_71),
.A2(n_96),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_71),
.A2(n_128),
.B1(n_130),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_72),
.A2(n_76),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_74),
.B(n_149),
.CON(n_148),
.SN(n_148)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_78),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_76),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.C(n_99),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_86),
.B(n_92),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_87),
.A2(n_157),
.B(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_102),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_102),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_112),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_126),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_113),
.A2(n_114),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_122),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_276),
.B(n_281),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_183),
.B(n_261),
.C(n_275),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_168),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_135),
.B(n_168),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_152),
.B2(n_167),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_138),
.B(n_139),
.C(n_167),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_158),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_153),
.B(n_160),
.C(n_164),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_156),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_169),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_178),
.B(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_260),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_255),
.B(n_259),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_243),
.B(n_254),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_225),
.B(n_242),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_214),
.B(n_224),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_203),
.B(n_213),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_195),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_199),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_208),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_240),
.B2(n_241),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_252),
.C(n_253),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_269),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule