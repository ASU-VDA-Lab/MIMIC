module fake_jpeg_18979_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_1),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_21),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_5),
.B1(n_11),
.B2(n_8),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_19),
.C(n_16),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_9),
.B1(n_13),
.B2(n_15),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

FAx1_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_19),
.CI(n_17),
.CON(n_29),
.SN(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_29),
.C(n_32),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_24),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_29),
.B1(n_33),
.B2(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_36),
.C(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_27),
.Y(n_45)
);


endmodule