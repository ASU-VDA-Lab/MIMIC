module fake_jpeg_14507_n_41 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_37;
wire n_29;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_8),
.Y(n_22)
);

HAxp5_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_4),
.CON(n_23),
.SN(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_1),
.C(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_13),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_35),
.B(n_34),
.C(n_30),
.D(n_28),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_31),
.Y(n_38)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_31),
.A3(n_29),
.B1(n_22),
.B2(n_26),
.C1(n_23),
.C2(n_20),
.Y(n_40)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_22),
.C(n_27),
.Y(n_41)
);


endmodule