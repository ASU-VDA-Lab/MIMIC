module fake_jpeg_9283_n_30 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_5),
.A2(n_7),
.B1(n_3),
.B2(n_6),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

OAI221xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_9),
.B2(n_11),
.C(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_15),
.C(n_14),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_2),
.B(n_8),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_14),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_22),
.Y(n_30)
);


endmodule