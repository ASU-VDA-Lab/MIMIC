module real_jpeg_12048_n_16 (n_5, n_4, n_8, n_0, n_12, n_251, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_251;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_69),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_70),
.B1(n_73),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_80),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_80),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_70),
.B1(n_73),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_7),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_114),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_114),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_10),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_11),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_73),
.B(n_76),
.C(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_70),
.B1(n_73),
.B2(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_13),
.B(n_81),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_103),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_13),
.A2(n_24),
.B1(n_36),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_13),
.B(n_109),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_14),
.A2(n_64),
.B1(n_70),
.B2(n_73),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_64),
.Y(n_152)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_142),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_20),
.B(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_94),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_21),
.B(n_82),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_22),
.B(n_55),
.C(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_23),
.B(n_39),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_24),
.A2(n_36),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_24),
.A2(n_36),
.B1(n_213),
.B2(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_24),
.A2(n_85),
.B(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_25),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_25),
.A2(n_35),
.B(n_86),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_25),
.A2(n_30),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_26),
.B(n_41),
.C(n_103),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_26),
.B(n_219),
.Y(n_218)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_36),
.A2(n_87),
.B(n_100),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_36),
.B(n_103),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_49),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_40),
.B(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_40),
.B(n_103),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_45),
.A2(n_58),
.B(n_182),
.C(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_45),
.B(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_46),
.B(n_59),
.C(n_61),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_52),
.A2(n_92),
.B(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_52),
.A2(n_124),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_52),
.A2(n_91),
.B1(n_189),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_52),
.A2(n_91),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_52),
.A2(n_91),
.B1(n_198),
.B2(n_208),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_56),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_56),
.A2(n_106),
.B1(n_109),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_56),
.A2(n_109),
.B1(n_170),
.B2(n_183),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_57),
.A2(n_107),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_62),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_77),
.B(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g183 ( 
.A(n_62),
.B(n_103),
.CON(n_183),
.SN(n_183)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_74),
.B1(n_79),
.B2(n_81),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_74),
.A2(n_81),
.B1(n_113),
.B2(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_93),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_93),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_152),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_110),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_96),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_104),
.B(n_110),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_140),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_138),
.B2(n_139),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_158),
.B1(n_174),
.B2(n_249),
.C(n_251),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_144),
.B(n_146),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_157),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_153),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_172),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_159),
.B(n_172),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_160),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_164),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_168),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_248),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_243),
.B(n_247),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_199),
.B(n_242),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_194),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_178),
.B(n_194),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_191),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_186),
.C(n_191),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_185),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B(n_190),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_197),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_237),
.B(n_241),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_227),
.B(n_236),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_216),
.B(n_226),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_209),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B(n_225),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_232),
.C(n_235),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_246),
.Y(n_247)
);


endmodule