module fake_jpeg_21031_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_44),
.B1(n_38),
.B2(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_14),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_18),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_67),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_20),
.B1(n_44),
.B2(n_38),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_79),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_17),
.B(n_29),
.C(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_51),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_34),
.B1(n_33),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_89),
.B1(n_93),
.B2(n_43),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_33),
.B1(n_34),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_78),
.B1(n_51),
.B2(n_19),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_84),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_88),
.Y(n_94)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_51),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_43),
.B1(n_42),
.B2(n_24),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_22),
.B(n_51),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_97),
.B(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_115),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_4),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_6),
.C(n_8),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_72),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_131),
.Y(n_144)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_99),
.B1(n_102),
.B2(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_102),
.B1(n_111),
.B2(n_103),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_141),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_130),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_127),
.C(n_117),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_114),
.B(n_105),
.Y(n_141)
);

AO21x2_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_101),
.B(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_95),
.B1(n_115),
.B2(n_98),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_95),
.B1(n_126),
.B2(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_153),
.B1(n_142),
.B2(n_152),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_155),
.B1(n_156),
.B2(n_122),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_154),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_129),
.B(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_145),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_139),
.C(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_151),
.C(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_160),
.C(n_163),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_152),
.B1(n_132),
.B2(n_142),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_165),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_149),
.B1(n_141),
.B2(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_171),
.B1(n_163),
.B2(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_141),
.B1(n_95),
.B2(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_140),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_178),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_92),
.B1(n_98),
.B2(n_88),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.C(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_70),
.B1(n_90),
.B2(n_65),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

NOR4xp25_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_181),
.D(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_82),
.C(n_87),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_84),
.B1(n_10),
.B2(n_11),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_9),
.Y(n_187)
);


endmodule