module fake_jpeg_18589_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_5),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_9),
.B1(n_10),
.B2(n_20),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_3),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

OA22x2_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_8),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_20),
.B(n_14),
.C(n_16),
.D(n_12),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_25),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_25),
.B1(n_15),
.B2(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_18),
.B1(n_19),
.B2(n_13),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.C(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_32),
.Y(n_34)
);


endmodule