module real_aes_7892_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_0), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_1), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g456 ( .A(n_1), .Y(n_456) );
INVx1_ASAP7_75t_L g486 ( .A(n_2), .Y(n_486) );
INVx1_ASAP7_75t_L g198 ( .A(n_3), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_4), .A2(n_39), .B1(n_159), .B2(n_516), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g166 ( .A1(n_5), .A2(n_140), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_6), .B(n_133), .Y(n_499) );
AND2x6_ASAP7_75t_L g145 ( .A(n_7), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_8), .A2(n_248), .B(n_249), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_9), .B(n_40), .Y(n_112) );
INVx1_ASAP7_75t_L g173 ( .A(n_10), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_11), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g138 ( .A(n_12), .Y(n_138) );
INVx1_ASAP7_75t_L g480 ( .A(n_13), .Y(n_480) );
INVx1_ASAP7_75t_L g254 ( .A(n_14), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_15), .B(n_181), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_16), .A2(n_102), .B1(n_113), .B2(n_775), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_17), .B(n_134), .Y(n_557) );
AO32x2_ASAP7_75t_L g529 ( .A1(n_18), .A2(n_133), .A3(n_178), .B1(n_508), .B2(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_19), .A2(n_63), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_19), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_20), .B(n_159), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_21), .B(n_154), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_22), .B(n_134), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_23), .A2(n_51), .B1(n_159), .B2(n_516), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_24), .B(n_140), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_25), .A2(n_77), .B1(n_159), .B2(n_181), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_26), .B(n_159), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_27), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_28), .A2(n_252), .B(n_253), .C(n_255), .Y(n_251) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_29), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_30), .B(n_175), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_31), .B(n_171), .Y(n_200) );
INVx1_ASAP7_75t_L g187 ( .A(n_32), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_33), .B(n_175), .Y(n_546) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_35), .B(n_159), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_36), .B(n_175), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_37), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_38), .A2(n_145), .B(n_149), .C(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g185 ( .A(n_41), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_42), .B(n_171), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_43), .B(n_159), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_44), .A2(n_87), .B1(n_217), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_45), .B(n_159), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_46), .B(n_159), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_47), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_48), .A2(n_70), .B1(n_760), .B2(n_761), .Y(n_759) );
CKINVDCx16_ASAP7_75t_R g761 ( .A(n_48), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_49), .B(n_485), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_50), .B(n_140), .Y(n_242) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_52), .A2(n_61), .B1(n_159), .B2(n_181), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_53), .A2(n_149), .B1(n_181), .B2(n_183), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_54), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_55), .B(n_159), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_56), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_57), .B(n_159), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_58), .A2(n_158), .B(n_170), .C(n_172), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_59), .Y(n_230) );
INVx1_ASAP7_75t_L g168 ( .A(n_60), .Y(n_168) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
INVx1_ASAP7_75t_L g122 ( .A(n_63), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_64), .B(n_159), .Y(n_487) );
INVx1_ASAP7_75t_L g137 ( .A(n_65), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
AO32x2_ASAP7_75t_L g513 ( .A1(n_67), .A2(n_133), .A3(n_234), .B1(n_508), .B2(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g506 ( .A(n_68), .Y(n_506) );
INVx1_ASAP7_75t_L g541 ( .A(n_69), .Y(n_541) );
INVx1_ASAP7_75t_L g760 ( .A(n_70), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_SL g153 ( .A1(n_71), .A2(n_154), .B(n_155), .C(n_158), .Y(n_153) );
INVxp67_ASAP7_75t_L g156 ( .A(n_72), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_73), .B(n_181), .Y(n_542) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_75), .Y(n_191) );
INVx1_ASAP7_75t_L g223 ( .A(n_76), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_78), .A2(n_145), .B(n_149), .C(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_79), .B(n_516), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_80), .B(n_181), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_81), .B(n_199), .Y(n_213) );
INVx2_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_83), .B(n_154), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_84), .B(n_181), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_85), .A2(n_145), .B(n_149), .C(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g107 ( .A(n_86), .Y(n_107) );
OR2x2_ASAP7_75t_L g453 ( .A(n_86), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g464 ( .A(n_86), .B(n_455), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_88), .A2(n_100), .B1(n_181), .B2(n_182), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_89), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_90), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_91), .A2(n_145), .B(n_149), .C(n_237), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_92), .Y(n_244) );
INVx1_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_94), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_95), .B(n_199), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_96), .B(n_181), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_97), .B(n_133), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_99), .A2(n_140), .B(n_147), .Y(n_139) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_104), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x2_ASAP7_75t_L g467 ( .A(n_107), .B(n_455), .Y(n_467) );
NOR2x2_ASAP7_75t_L g771 ( .A(n_107), .B(n_454), .Y(n_771) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g455 ( .A(n_112), .B(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_460), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g774 ( .A(n_116), .Y(n_774) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_450), .B(n_457), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_449), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g449 ( .A(n_124), .Y(n_449) );
INVx1_ASAP7_75t_SL g465 ( .A(n_124), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_124), .A2(n_763), .B1(n_765), .B2(n_766), .Y(n_762) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND4x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_367), .C(n_414), .D(n_434), .Y(n_125) );
NOR3xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_297), .C(n_322), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_205), .B(n_257), .C(n_287), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_176), .Y(n_129) );
INVx3_ASAP7_75t_SL g339 ( .A(n_130), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_130), .B(n_270), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_130), .B(n_192), .Y(n_420) );
AND2x2_ASAP7_75t_L g443 ( .A(n_130), .B(n_309), .Y(n_443) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_164), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g261 ( .A(n_132), .B(n_165), .Y(n_261) );
INVx3_ASAP7_75t_L g274 ( .A(n_132), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_132), .B(n_164), .Y(n_279) );
OR2x2_ASAP7_75t_L g330 ( .A(n_132), .B(n_271), .Y(n_330) );
BUFx2_ASAP7_75t_L g350 ( .A(n_132), .Y(n_350) );
AND2x2_ASAP7_75t_L g360 ( .A(n_132), .B(n_271), .Y(n_360) );
AND2x2_ASAP7_75t_L g366 ( .A(n_132), .B(n_177), .Y(n_366) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_161), .Y(n_132) );
INVx4_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_492), .B(n_499), .Y(n_491) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_135), .B(n_136), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g248 ( .A(n_140), .Y(n_248) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_141), .B(n_145), .Y(n_189) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g485 ( .A(n_142), .Y(n_485) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
INVx4_ASAP7_75t_SL g160 ( .A(n_145), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_145), .A2(n_479), .B(n_483), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_145), .A2(n_493), .B(n_496), .Y(n_492) );
BUFx3_ASAP7_75t_L g508 ( .A(n_145), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_145), .A2(n_521), .B(n_525), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_145), .A2(n_540), .B(n_543), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_153), .C(n_160), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_148), .A2(n_160), .B(n_168), .C(n_169), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_148), .A2(n_160), .B(n_250), .C(n_251), .Y(n_249) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
INVx1_ASAP7_75t_L g516 ( .A(n_150), .Y(n_516) );
INVx1_ASAP7_75t_L g524 ( .A(n_154), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_157), .B(n_173), .Y(n_172) );
INVx5_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g514 ( .A1(n_157), .A2(n_171), .B1(n_515), .B2(n_517), .Y(n_514) );
O2A1O1Ixp5_ASAP7_75t_SL g540 ( .A1(n_158), .A2(n_199), .B(n_541), .C(n_542), .Y(n_540) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_159), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_160), .A2(n_180), .B1(n_188), .B2(n_189), .Y(n_179) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_162), .A2(n_166), .B(n_174), .Y(n_165) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_163), .B(n_220), .Y(n_219) );
AO21x1_ASAP7_75t_L g552 ( .A1(n_163), .A2(n_553), .B(n_556), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_163), .B(n_508), .C(n_553), .Y(n_571) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_165), .B(n_271), .Y(n_285) );
INVx2_ASAP7_75t_L g295 ( .A(n_165), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_165), .B(n_274), .Y(n_308) );
OR2x2_ASAP7_75t_L g319 ( .A(n_165), .B(n_271), .Y(n_319) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_165), .B(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g377 ( .A(n_165), .Y(n_377) );
AND2x2_ASAP7_75t_L g423 ( .A(n_165), .B(n_177), .Y(n_423) );
O2A1O1Ixp5_ASAP7_75t_L g505 ( .A1(n_170), .A2(n_484), .B(n_506), .C(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_170), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_171), .A2(n_488), .B1(n_531), .B2(n_532), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_171), .A2(n_488), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g204 ( .A(n_175), .Y(n_204) );
INVx2_ASAP7_75t_L g234 ( .A(n_175), .Y(n_234) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_175), .A2(n_247), .B(n_256), .Y(n_246) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_175), .A2(n_520), .B(n_528), .Y(n_519) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_175), .A2(n_539), .B(n_546), .Y(n_538) );
INVx3_ASAP7_75t_SL g296 ( .A(n_176), .Y(n_296) );
OR2x2_ASAP7_75t_L g349 ( .A(n_176), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
INVx3_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g338 ( .A(n_177), .B(n_193), .Y(n_338) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_177), .Y(n_406) );
AOI33xp33_ASAP7_75t_L g410 ( .A1(n_177), .A2(n_339), .A3(n_346), .B1(n_355), .B2(n_411), .B3(n_412), .Y(n_410) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_190), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_178), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_178), .A2(n_194), .B(n_202), .Y(n_193) );
INVx2_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
INVx2_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_183) );
INVx2_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
INVx4_ASAP7_75t_L g252 ( .A(n_184), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g259 ( .A(n_192), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_192), .B(n_274), .Y(n_273) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_192), .B(n_334), .C(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g359 ( .A(n_192), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_192), .B(n_366), .Y(n_369) );
AND2x2_ASAP7_75t_L g422 ( .A(n_192), .B(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
OR2x2_ASAP7_75t_L g372 ( .A(n_193), .B(n_271), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g488 ( .A(n_199), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_199), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_199), .A2(n_503), .B(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_201), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_204), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_204), .B(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_231), .Y(n_205) );
AOI32xp33_ASAP7_75t_L g323 ( .A1(n_206), .A2(n_324), .A3(n_326), .B1(n_328), .B2(n_331), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_206), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g426 ( .A(n_206), .Y(n_426) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g358 ( .A(n_207), .B(n_342), .Y(n_358) );
AND2x2_ASAP7_75t_L g378 ( .A(n_207), .B(n_304), .Y(n_378) );
AND2x2_ASAP7_75t_L g446 ( .A(n_207), .B(n_364), .Y(n_446) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_221), .Y(n_207) );
INVx3_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_208), .B(n_265), .Y(n_281) );
OR2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_264), .Y(n_286) );
INVx1_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_208), .B(n_275), .Y(n_301) );
AND2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_208), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g356 ( .A(n_208), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_208), .B(n_441), .Y(n_440) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_218), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
INVx1_ASAP7_75t_L g228 ( .A(n_218), .Y(n_228) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_218), .A2(n_478), .B(n_489), .Y(n_477) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_218), .A2(n_501), .B(n_509), .Y(n_500) );
INVx2_ASAP7_75t_L g265 ( .A(n_221), .Y(n_265) );
AND2x2_ASAP7_75t_L g311 ( .A(n_221), .B(n_232), .Y(n_311) );
AND2x2_ASAP7_75t_L g321 ( .A(n_221), .B(n_246), .Y(n_321) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .B(n_229), .Y(n_221) );
INVx2_ASAP7_75t_L g441 ( .A(n_231), .Y(n_441) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_245), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_232), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g342 ( .A(n_232), .B(n_305), .Y(n_342) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g290 ( .A(n_233), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_233), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_233), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_233), .B(n_265), .Y(n_387) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_243), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_241), .Y(n_237) );
AND2x2_ASAP7_75t_L g266 ( .A(n_245), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g327 ( .A(n_245), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_245), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g364 ( .A(n_245), .Y(n_364) );
INVx1_ASAP7_75t_L g397 ( .A(n_245), .Y(n_397) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g275 ( .A(n_246), .B(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_252), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g482 ( .A(n_252), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_252), .A2(n_544), .B(n_545), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B1(n_268), .B2(n_275), .C(n_276), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_259), .B(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_259), .B(n_342), .Y(n_419) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_261), .B(n_309), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_261), .B(n_270), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_261), .B(n_284), .Y(n_413) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
AND2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g388 ( .A(n_266), .Y(n_388) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_267), .B(n_290), .Y(n_336) );
AND2x2_ASAP7_75t_L g400 ( .A(n_267), .B(n_326), .Y(n_400) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g309 ( .A(n_271), .B(n_278), .Y(n_309) );
AND2x2_ASAP7_75t_L g405 ( .A(n_272), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_274), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_275), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_275), .B(n_282), .Y(n_370) );
AND2x2_ASAP7_75t_L g390 ( .A(n_275), .B(n_290), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_275), .B(n_355), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .A3(n_282), .B1(n_283), .B2(n_286), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_SL g284 ( .A(n_278), .Y(n_284) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_278), .B(n_308), .Y(n_325) );
OR2x2_ASAP7_75t_L g329 ( .A(n_278), .B(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_278), .B(n_377), .Y(n_430) );
INVx1_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_280), .A2(n_371), .B1(n_417), .B2(n_420), .C(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_281), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g331 ( .A(n_281), .B(n_304), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_281), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g409 ( .A(n_281), .B(n_342), .Y(n_409) );
INVxp67_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g415 ( .A(n_284), .B(n_402), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_284), .B(n_365), .Y(n_438) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_286), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g431 ( .A(n_286), .B(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_291), .B(n_294), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_289), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g384 ( .A(n_293), .B(n_304), .Y(n_384) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g402 ( .A(n_295), .B(n_360), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_295), .B(n_359), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_296), .B(n_308), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .C(n_312), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_298), .A2(n_333), .B1(n_337), .B2(n_340), .C(n_343), .Y(n_332) );
AOI31xp33_ASAP7_75t_L g427 ( .A1(n_298), .A2(n_428), .A3(n_429), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_308), .B2(n_310), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g428 ( .A(n_308), .Y(n_428) );
INVx1_ASAP7_75t_L g391 ( .A(n_309), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g434 ( .A1(n_311), .A2(n_435), .B(n_437), .C(n_439), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_316), .B2(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_317), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_319), .A2(n_353), .B1(n_372), .B2(n_408), .C(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g403 ( .A(n_320), .Y(n_403) );
INVx1_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_332), .C(n_347), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_374), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_326), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g433 ( .A(n_327), .Y(n_433) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g371 ( .A(n_334), .B(n_354), .Y(n_371) );
INVx1_ASAP7_75t_L g346 ( .A(n_335), .Y(n_346) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_338), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_338), .B(n_376), .Y(n_375) );
NOR4xp25_ASAP7_75t_L g343 ( .A(n_339), .B(n_344), .C(n_345), .D(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_352), .B1(n_358), .B2(n_359), .C1(n_361), .C2(n_365), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g445 ( .A(n_349), .Y(n_445) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_361), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_366), .A2(n_422), .B(n_424), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_379), .C(n_392), .D(n_407), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_372), .C(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g448 ( .A(n_369), .Y(n_448) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_376), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_385), .B2(n_386), .C1(n_389), .C2(n_391), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_415), .B(n_416), .C(n_427), .Y(n_414) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_398), .B1(n_399), .B2(n_401), .C1(n_403), .C2(n_404), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_409), .A2(n_412), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_442), .B(n_444), .C(n_447), .Y(n_439) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g458 ( .A(n_453), .Y(n_458) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_457), .A2(n_461), .B(n_773), .Y(n_460) );
NOR2xp33_ASAP7_75t_SL g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OAI222xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_759), .B1(n_762), .B2(n_767), .C1(n_768), .C2(n_772), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_466), .B2(n_468), .Y(n_462) );
INVx2_ASAP7_75t_L g764 ( .A(n_463), .Y(n_764) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g765 ( .A(n_467), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_468), .Y(n_766) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_469), .B(n_725), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_629), .C(n_713), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_572), .C(n_594), .D(n_610), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_510), .B1(n_533), .B2(n_551), .C(n_558), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_490), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_474), .B(n_551), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_474), .B(n_612), .C(n_625), .D(n_627), .Y(n_624) );
INVxp67_ASAP7_75t_L g741 ( .A(n_474), .Y(n_741) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g623 ( .A(n_475), .B(n_561), .Y(n_623) );
AND2x2_ASAP7_75t_L g647 ( .A(n_475), .B(n_490), .Y(n_647) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g614 ( .A(n_476), .B(n_550), .Y(n_614) );
AND2x2_ASAP7_75t_L g654 ( .A(n_476), .B(n_635), .Y(n_654) );
AND2x2_ASAP7_75t_L g671 ( .A(n_476), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_476), .B(n_491), .Y(n_695) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g549 ( .A(n_477), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g566 ( .A(n_477), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g578 ( .A(n_477), .B(n_491), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_477), .B(n_500), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B(n_487), .C(n_488), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_488), .A2(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_L g581 ( .A(n_490), .B(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_490), .A2(n_631), .B1(n_634), .B2(n_636), .C(n_640), .Y(n_630) );
AND2x2_ASAP7_75t_L g689 ( .A(n_490), .B(n_654), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_490), .B(n_671), .Y(n_723) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
INVx3_ASAP7_75t_L g550 ( .A(n_491), .Y(n_550) );
AND2x2_ASAP7_75t_L g598 ( .A(n_491), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g652 ( .A(n_491), .B(n_567), .Y(n_652) );
AND2x2_ASAP7_75t_L g710 ( .A(n_491), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g551 ( .A(n_500), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
INVx1_ASAP7_75t_L g622 ( .A(n_500), .Y(n_622) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_500), .Y(n_628) );
AND2x2_ASAP7_75t_L g673 ( .A(n_500), .B(n_550), .Y(n_673) );
OR2x2_ASAP7_75t_L g712 ( .A(n_500), .B(n_552), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_505), .B(n_508), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_510), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .Y(n_510) );
AND2x2_ASAP7_75t_L g708 ( .A(n_511), .B(n_705), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_511), .B(n_690), .Y(n_740) );
BUFx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g639 ( .A(n_512), .B(n_563), .Y(n_639) );
AND2x2_ASAP7_75t_L g688 ( .A(n_512), .B(n_536), .Y(n_688) );
INVx1_ASAP7_75t_L g734 ( .A(n_512), .Y(n_734) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_513), .Y(n_548) );
AND2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_563), .Y(n_589) );
INVx1_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
AND2x2_ASAP7_75t_L g612 ( .A(n_513), .B(n_529), .Y(n_612) );
AND2x2_ASAP7_75t_L g680 ( .A(n_518), .B(n_588), .Y(n_680) );
INVx2_ASAP7_75t_L g745 ( .A(n_518), .Y(n_745) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
AND2x2_ASAP7_75t_L g562 ( .A(n_519), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g575 ( .A(n_519), .B(n_537), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_519), .B(n_536), .Y(n_603) );
INVx1_ASAP7_75t_L g609 ( .A(n_519), .Y(n_609) );
INVx1_ASAP7_75t_L g626 ( .A(n_519), .Y(n_626) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_519), .Y(n_638) );
INVx2_ASAP7_75t_L g706 ( .A(n_519), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g563 ( .A(n_529), .Y(n_563) );
BUFx2_ASAP7_75t_L g660 ( .A(n_529), .Y(n_660) );
AND2x2_ASAP7_75t_L g705 ( .A(n_529), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_547), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_535), .B(n_642), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_535), .A2(n_704), .B(n_718), .Y(n_728) );
AND2x2_ASAP7_75t_L g753 ( .A(n_535), .B(n_639), .Y(n_753) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g675 ( .A(n_537), .Y(n_675) );
AND2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_538), .Y(n_588) );
INVx2_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_538), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g561 ( .A(n_548), .Y(n_561) );
OR2x2_ASAP7_75t_L g574 ( .A(n_548), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g642 ( .A(n_548), .B(n_638), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_548), .B(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g743 ( .A(n_548), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_548), .B(n_680), .Y(n_755) );
AND2x2_ASAP7_75t_L g634 ( .A(n_549), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g657 ( .A(n_549), .B(n_551), .Y(n_657) );
INVx2_ASAP7_75t_L g569 ( .A(n_550), .Y(n_569) );
AND2x2_ASAP7_75t_L g597 ( .A(n_550), .B(n_570), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_550), .B(n_622), .Y(n_678) );
AND2x2_ASAP7_75t_L g592 ( .A(n_551), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g739 ( .A(n_551), .Y(n_739) );
AND2x2_ASAP7_75t_L g751 ( .A(n_551), .B(n_614), .Y(n_751) );
AND2x2_ASAP7_75t_L g577 ( .A(n_552), .B(n_567), .Y(n_577) );
INVx1_ASAP7_75t_L g672 ( .A(n_552), .Y(n_672) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g570 ( .A(n_557), .B(n_571), .Y(n_570) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_561), .B(n_608), .Y(n_617) );
OR2x2_ASAP7_75t_L g749 ( .A(n_561), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g666 ( .A(n_562), .B(n_607), .Y(n_666) );
AND2x2_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g733 ( .A(n_562), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g757 ( .A(n_562), .B(n_604), .Y(n_757) );
NOR2xp67_ASAP7_75t_L g715 ( .A(n_563), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g744 ( .A(n_563), .B(n_607), .Y(n_744) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
AND2x2_ASAP7_75t_L g596 ( .A(n_566), .B(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g758 ( .A(n_566), .Y(n_758) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g593 ( .A(n_569), .Y(n_593) );
AND2x2_ASAP7_75t_L g644 ( .A(n_569), .B(n_577), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_569), .B(n_712), .Y(n_738) );
INVx2_ASAP7_75t_L g583 ( .A(n_570), .Y(n_583) );
INVx3_ASAP7_75t_L g635 ( .A(n_570), .Y(n_635) );
OR2x2_ASAP7_75t_L g663 ( .A(n_570), .B(n_664), .Y(n_663) );
AOI311xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .A3(n_578), .B(n_579), .C(n_590), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_573), .A2(n_611), .B(n_613), .C(n_615), .Y(n_610) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g595 ( .A(n_575), .Y(n_595) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g613 ( .A(n_577), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_577), .B(n_593), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_577), .B(n_578), .Y(n_746) );
AND2x2_ASAP7_75t_L g668 ( .A(n_578), .B(n_582), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_585), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g726 ( .A(n_582), .B(n_614), .Y(n_726) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_583), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_L g611 ( .A(n_587), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g656 ( .A(n_589), .Y(n_656) );
AND2x4_ASAP7_75t_L g718 ( .A(n_589), .B(n_687), .Y(n_718) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_592), .A2(n_658), .B1(n_670), .B2(n_674), .C1(n_676), .C2(n_680), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_598), .C(n_601), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_595), .B(n_639), .Y(n_662) );
INVx1_ASAP7_75t_L g684 ( .A(n_597), .Y(n_684) );
INVx1_ASAP7_75t_L g618 ( .A(n_599), .Y(n_618) );
OR2x2_ASAP7_75t_L g683 ( .A(n_600), .B(n_684), .Y(n_683) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_604), .B(n_608), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_602), .B(n_620), .C(n_621), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_602), .A2(n_639), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_606), .Y(n_659) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_607), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g716 ( .A(n_607), .Y(n_716) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_607), .Y(n_732) );
INVx2_ASAP7_75t_L g690 ( .A(n_608), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_612), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g664 ( .A(n_614), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B1(n_619), .B2(n_623), .C(n_624), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_618), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g752 ( .A(n_618), .Y(n_752) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g633 ( .A(n_625), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_625), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g691 ( .A(n_625), .B(n_639), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_625), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g724 ( .A(n_625), .B(n_659), .Y(n_724) );
BUFx3_ASAP7_75t_L g687 ( .A(n_626), .Y(n_687) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND5xp2_ASAP7_75t_L g629 ( .A(n_630), .B(n_648), .C(n_669), .D(n_681), .E(n_696), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI32xp33_ASAP7_75t_L g721 ( .A1(n_633), .A2(n_660), .A3(n_676), .B1(n_722), .B2(n_724), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_635), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g645 ( .A(n_639), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_645), .B2(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_655), .B1(n_657), .B2(n_658), .C(n_661), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g720 ( .A(n_652), .B(n_671), .Y(n_720) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_657), .A2(n_718), .B1(n_736), .B2(n_741), .C(n_742), .Y(n_735) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g701 ( .A(n_660), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_667), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g679 ( .A(n_671), .Y(n_679) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B1(n_689), .B2(n_690), .C1(n_691), .C2(n_692), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_690), .A2(n_737), .B1(n_739), .B2(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_702), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_707), .B(n_709), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g750 ( .A(n_705), .Y(n_750) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B(n_719), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_729), .C(n_754), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g730 ( .A(n_726), .Y(n_730) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI211xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_735), .C(n_747), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .B(n_746), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI21xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g767 ( .A(n_759), .Y(n_767) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
endmodule