module real_jpeg_14254_n_6 (n_5, n_4, n_0, n_1, n_41, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_41;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_15),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_18),
.B(n_22),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_10),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B(n_23),
.C(n_32),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_14),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_14),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

AOI211xp5_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_12),
.B(n_28),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

OAI322xp33_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_21),
.A3(n_28),
.B1(n_33),
.B2(n_34),
.C1(n_35),
.C2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);


endmodule