module fake_aes_4083_n_565 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_565);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_565;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_20), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_64), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_37), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_42), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_28), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_33), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_0), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_57), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_9), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_54), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_70), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_52), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_22), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_44), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_74), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_7), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_36), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_72), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_7), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_18), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_66), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_27), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_80), .Y(n_117) );
BUFx8_ASAP7_75t_L g118 ( .A(n_105), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_102), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_107), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_84), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
NAND2xp33_ASAP7_75t_SL g125 ( .A(n_105), .B(n_2), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_111), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_92), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_90), .B(n_5), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_84), .B(n_6), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_140), .B(n_94), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_126), .B(n_93), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_138), .B(n_97), .Y(n_144) );
BUFx10_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_120), .Y(n_147) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_122), .A2(n_99), .B(n_114), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
NOR2xp33_ASAP7_75t_SL g151 ( .A(n_118), .B(n_88), .Y(n_151) );
OR2x2_ASAP7_75t_L g152 ( .A(n_140), .B(n_108), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_138), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_118), .B(n_115), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_128), .A2(n_88), .B1(n_96), .B2(n_95), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_123), .B(n_100), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_115), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_124), .B(n_98), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_124), .B(n_104), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_162), .B(n_127), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_161), .A2(n_125), .B1(n_137), .B2(n_134), .Y(n_171) );
NAND2xp33_ASAP7_75t_SL g172 ( .A(n_156), .B(n_96), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_143), .A2(n_137), .B(n_134), .Y(n_173) );
NOR2xp67_ASAP7_75t_L g174 ( .A(n_146), .B(n_119), .Y(n_174) );
BUFx6f_ASAP7_75t_SL g175 ( .A(n_161), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_145), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_167), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_164), .B(n_127), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_147), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_155), .B(n_98), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_145), .Y(n_184) );
NAND3xp33_ASAP7_75t_L g185 ( .A(n_161), .B(n_133), .C(n_121), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_167), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_141), .B(n_133), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_158), .B(n_135), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_166), .B(n_119), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_166), .B(n_121), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_166), .A2(n_139), .B1(n_103), .B2(n_116), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_144), .B(n_132), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_155), .B(n_110), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_149), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_155), .B(n_132), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
NOR2xp33_ASAP7_75t_R g204 ( .A(n_179), .B(n_102), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_175), .A2(n_159), .B1(n_112), .B2(n_144), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_172), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_188), .A2(n_152), .B(n_142), .C(n_149), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_170), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_SL g209 ( .A1(n_173), .A2(n_131), .B(n_165), .C(n_154), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_190), .A2(n_152), .B(n_165), .C(n_160), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_170), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_169), .A2(n_155), .B(n_148), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_178), .A2(n_148), .B(n_163), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_180), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_185), .A2(n_154), .B(n_157), .C(n_160), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_180), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_186), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_183), .B(n_144), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
BUFx8_ASAP7_75t_SL g220 ( .A(n_189), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_185), .A2(n_163), .B(n_157), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_SL g223 ( .A1(n_192), .A2(n_153), .B(n_150), .C(n_163), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_183), .B(n_148), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_198), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_168), .B(n_145), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_193), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_183), .B(n_148), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_191), .B(n_153), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_174), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_192), .B(n_153), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_193), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_208), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_205), .A2(n_175), .B1(n_189), .B2(n_171), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_193), .B(n_187), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_218), .B(n_201), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_208), .B(n_189), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_212), .A2(n_202), .B(n_197), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_208), .B(n_189), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_222), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_211), .Y(n_248) );
NOR2x1_ASAP7_75t_SL g249 ( .A(n_227), .B(n_201), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_218), .B(n_194), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_227), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_207), .B(n_171), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_222), .A2(n_175), .B1(n_189), .B2(n_199), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_226), .A2(n_174), .B1(n_112), .B2(n_181), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_211), .A2(n_187), .B(n_195), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_218), .B(n_200), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_231), .B(n_200), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_217), .A2(n_177), .B(n_195), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_219), .B(n_182), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_203), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_231), .B(n_200), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_219), .A2(n_196), .B(n_177), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_210), .B(n_182), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_225), .B(n_182), .Y(n_265) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_209), .A2(n_89), .B(n_167), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_238), .B(n_225), .Y(n_267) );
AOI21xp33_ASAP7_75t_L g268 ( .A1(n_252), .A2(n_223), .B(n_230), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_238), .B(n_230), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_240), .A2(n_233), .B(n_235), .C(n_194), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_247), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_247), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_244), .A2(n_215), .B(n_235), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_243), .A2(n_220), .B1(n_222), .B2(n_204), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_243), .A2(n_206), .B1(n_233), .B2(n_224), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_247), .B(n_224), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_245), .A2(n_224), .B1(n_228), .B2(n_234), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_245), .A2(n_224), .B1(n_228), .B2(n_234), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_246), .B(n_232), .Y(n_280) );
OAI21x1_ASAP7_75t_SL g281 ( .A1(n_249), .A2(n_251), .B(n_248), .Y(n_281) );
OAI21xp33_ASAP7_75t_SL g282 ( .A1(n_251), .A2(n_221), .B(n_236), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_251), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_221), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_241), .A2(n_236), .B(n_229), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_228), .B1(n_234), .B2(n_203), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_257), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_260), .B(n_232), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_255), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_285), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_239), .Y(n_292) );
NAND2xp33_ASAP7_75t_R g293 ( .A(n_273), .B(n_8), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_270), .B(n_239), .Y(n_294) );
CKINVDCx14_ASAP7_75t_R g295 ( .A(n_270), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_290), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_254), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_277), .B(n_239), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
CKINVDCx8_ASAP7_75t_R g301 ( .A(n_281), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_269), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_288), .B(n_254), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_290), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_277), .B(n_249), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_277), .B(n_260), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_272), .B(n_265), .Y(n_308) );
BUFx4f_ASAP7_75t_L g309 ( .A(n_267), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_267), .B(n_261), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_296), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_291), .B(n_267), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_300), .Y(n_318) );
AOI211xp5_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_268), .B(n_283), .C(n_282), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
AOI33xp33_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_275), .A3(n_276), .B1(n_278), .B2(n_279), .B3(n_284), .Y(n_321) );
AOI211xp5_ASAP7_75t_SL g322 ( .A1(n_306), .A2(n_268), .B(n_283), .C(n_289), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_305), .B(n_284), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_312), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_284), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_302), .B(n_289), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_301), .B(n_281), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_298), .B(n_286), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_309), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_312), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_274), .B(n_286), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_311), .B(n_286), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_311), .B(n_282), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_292), .B(n_274), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
XNOR2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_242), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_309), .A2(n_264), .B1(n_271), .B2(n_287), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_306), .B(n_250), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_310), .B(n_266), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_303), .B(n_167), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_315), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_326), .B(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_326), .B(n_307), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_318), .B(n_306), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_336), .B(n_292), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_324), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_330), .B(n_310), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_341), .B(n_327), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_336), .B(n_294), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_323), .B(n_307), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_335), .B(n_310), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_322), .A2(n_293), .B(n_313), .C(n_308), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_333), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_314), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_333), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_325), .B(n_294), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_316), .B(n_313), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_321), .B(n_299), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_335), .B(n_299), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_328), .B(n_308), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
OAI222xp33_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_301), .B1(n_256), .B2(n_250), .C1(n_261), .C2(n_262), .Y(n_376) );
NOR3xp33_ASAP7_75t_SL g377 ( .A(n_339), .B(n_8), .C(n_9), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_341), .B(n_10), .Y(n_378) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_341), .B(n_84), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_84), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_331), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_342), .B(n_101), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_334), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_342), .B(n_101), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_334), .B(n_101), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_338), .B(n_11), .Y(n_386) );
AND2x2_ASAP7_75t_SL g387 ( .A(n_342), .B(n_258), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_338), .B(n_12), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_328), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_334), .B(n_101), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_368), .B(n_319), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_365), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_373), .B(n_332), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_373), .B(n_332), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_352), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_363), .A2(n_377), .B(n_378), .C(n_329), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_361), .B(n_332), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_361), .B(n_332), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_364), .B(n_337), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_347), .B(n_337), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_349), .B(n_319), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_345), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_374), .B(n_337), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_354), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_364), .B(n_340), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_360), .B(n_322), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_367), .B(n_340), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_351), .B(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_367), .B(n_343), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_358), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_357), .Y(n_417) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_387), .B(n_343), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_357), .Y(n_419) );
XNOR2xp5_ASAP7_75t_L g420 ( .A(n_387), .B(n_329), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_350), .B(n_101), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_357), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_371), .B(n_372), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_384), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_389), .B(n_339), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_389), .B(n_344), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_355), .B(n_329), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_362), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_362), .B(n_13), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_350), .B(n_109), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_350), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_363), .B(n_13), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_365), .B(n_14), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_366), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_366), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_369), .B(n_109), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_381), .B(n_14), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_386), .B(n_15), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_380), .B(n_15), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_388), .A2(n_113), .B1(n_109), .B2(n_266), .C(n_263), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_393), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_405), .B(n_380), .Y(n_446) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_415), .B(n_358), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_433), .A2(n_378), .B(n_379), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g452 ( .A(n_420), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_399), .A2(n_376), .B(n_109), .C(n_113), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_415), .B(n_358), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_424), .A2(n_113), .B1(n_109), .B2(n_390), .C(n_385), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_404), .B(n_385), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_390), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_416), .B(n_358), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_SL g459 ( .A1(n_399), .A2(n_16), .B(n_17), .C(n_263), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_442), .A2(n_113), .B1(n_266), .B2(n_16), .C(n_17), .Y(n_460) );
NAND2xp33_ASAP7_75t_L g461 ( .A(n_415), .B(n_113), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_414), .B(n_21), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_442), .A2(n_262), .B(n_258), .C(n_242), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_418), .A2(n_266), .B1(n_242), .B2(n_262), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_432), .B(n_241), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_409), .A2(n_262), .B1(n_258), .B2(n_242), .C(n_229), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_391), .B(n_259), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_421), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g472 ( .A(n_430), .B(n_256), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_403), .B(n_259), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_432), .B(n_23), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_421), .A2(n_258), .B1(n_236), .B2(n_229), .C(n_234), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_418), .A2(n_255), .B(n_256), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_426), .A2(n_256), .B1(n_250), .B2(n_228), .C(n_214), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_407), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_394), .B(n_26), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_406), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_443), .A2(n_29), .B(n_31), .C(n_32), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_431), .A2(n_237), .B1(n_216), .B2(n_203), .C(n_153), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_394), .B(n_396), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_406), .Y(n_487) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_408), .B(n_256), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g489 ( .A1(n_422), .A2(n_182), .B(n_39), .C(n_40), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_425), .A2(n_250), .B1(n_237), .B2(n_216), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_453), .A2(n_428), .B1(n_419), .B2(n_423), .C(n_417), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_481), .B(n_396), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_464), .Y(n_493) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_454), .B(n_410), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_452), .A2(n_400), .B1(n_401), .B2(n_439), .C(n_440), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_485), .B(n_401), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_461), .A2(n_438), .B(n_427), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_487), .B(n_400), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_486), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_445), .Y(n_502) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_454), .B(n_435), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_470), .A2(n_413), .B1(n_410), .B2(n_408), .Y(n_504) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_447), .B(n_438), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_448), .B(n_441), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
OAI32xp33_ASAP7_75t_L g508 ( .A1(n_470), .A2(n_427), .A3(n_413), .B1(n_436), .B2(n_437), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_471), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_462), .Y(n_510) );
OAI31xp33_ASAP7_75t_L g511 ( .A1(n_465), .A2(n_437), .A3(n_436), .B(n_392), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_478), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_479), .B(n_392), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_457), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_483), .Y(n_515) );
XOR2x2_ASAP7_75t_L g516 ( .A(n_472), .B(n_444), .Y(n_516) );
AOI22x1_ASAP7_75t_SL g517 ( .A1(n_459), .A2(n_34), .B1(n_41), .B2(n_43), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_488), .A2(n_476), .B1(n_489), .B2(n_446), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_466), .A2(n_250), .B1(n_237), .B2(n_216), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_468), .A2(n_184), .B1(n_176), .B2(n_150), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_510), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_508), .A2(n_460), .B1(n_450), .B2(n_477), .C(n_455), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_494), .A2(n_476), .B1(n_490), .B2(n_480), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_518), .A2(n_505), .B1(n_503), .B2(n_495), .Y(n_525) );
AOI211x1_ASAP7_75t_L g526 ( .A1(n_491), .A2(n_450), .B(n_474), .C(n_490), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_492), .B(n_467), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_519), .A2(n_469), .B1(n_463), .B2(n_482), .C(n_475), .Y(n_528) );
OAI21xp33_ASAP7_75t_L g529 ( .A1(n_504), .A2(n_473), .B(n_489), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_516), .A2(n_484), .B1(n_150), .B2(n_47), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_499), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_498), .A2(n_184), .B1(n_176), .B2(n_150), .Y(n_532) );
NOR4xp25_ASAP7_75t_L g533 ( .A(n_493), .B(n_45), .C(n_46), .D(n_48), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_506), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_506), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_501), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_497), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_511), .A2(n_53), .B(n_55), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
OAI221xp5_ASAP7_75t_SL g540 ( .A1(n_529), .A2(n_511), .B1(n_520), .B2(n_521), .C(n_500), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_525), .A2(n_500), .B1(n_514), .B2(n_496), .Y(n_541) );
OA211x2_ASAP7_75t_L g542 ( .A1(n_523), .A2(n_517), .B(n_513), .C(n_515), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_534), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_535), .B(n_512), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_531), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_524), .A2(n_507), .B(n_509), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_528), .A2(n_56), .B1(n_59), .B2(n_60), .Y(n_547) );
OA22x2_ASAP7_75t_SL g548 ( .A1(n_526), .A2(n_61), .B1(n_62), .B2(n_65), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_538), .A2(n_67), .B(n_68), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_540), .A2(n_522), .B(n_537), .C(n_530), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_541), .B(n_539), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_545), .Y(n_552) );
OAI22x1_ASAP7_75t_L g553 ( .A1(n_542), .A2(n_547), .B1(n_548), .B2(n_543), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_544), .B(n_536), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_554), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_550), .B(n_546), .C(n_537), .Y(n_556) );
AND4x1_ASAP7_75t_L g557 ( .A(n_551), .B(n_533), .C(n_549), .D(n_532), .Y(n_557) );
OAI21x1_ASAP7_75t_SL g558 ( .A1(n_555), .A2(n_552), .B(n_553), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_557), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_559), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_558), .Y(n_561) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_561), .A2(n_556), .B(n_527), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_562), .A2(n_560), .B(n_561), .Y(n_563) );
AOI322xp5_ASAP7_75t_L g564 ( .A1(n_563), .A2(n_533), .A3(n_73), .B1(n_75), .B2(n_76), .C1(n_69), .C2(n_78), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_564), .A2(n_77), .B(n_79), .Y(n_565) );
endmodule