module fake_netlist_5_646_n_774 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_774);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_774;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_753;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

BUFx10_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_65),
.B(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_53),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_R g165 ( 
.A(n_39),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_56),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_30),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_2),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_16),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_74),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_59),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_72),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_36),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_3),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_19),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_12),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_11),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_136),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_84),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_24),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_63),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_128),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_42),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_81),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_99),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_102),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_54),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_67),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_90),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_193),
.B(n_179),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_4),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_5),
.B(n_6),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_188),
.B(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_6),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_20),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_182),
.B(n_21),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_159),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_7),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_22),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_7),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_170),
.B(n_8),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_8),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_164),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_242),
.B(n_186),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_186),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_166),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_212),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

NOR2x1p5_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_173),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_206),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_174),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_177),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

NOR2x1p5_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_178),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_252),
.A2(n_202),
.B1(n_172),
.B2(n_160),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_183),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_187),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_227),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_257),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_225),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_190),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_234),
.A2(n_202),
.B1(n_172),
.B2(n_200),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_232),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_257),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_217),
.C(n_247),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_282),
.B(n_237),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_264),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_222),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_230),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_242),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_222),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_230),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_235),
.B1(n_254),
.B2(n_241),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_282),
.A2(n_248),
.B(n_216),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_222),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_222),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_230),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_230),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_248),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_248),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_269),
.B(n_237),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_294),
.B(n_237),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_225),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_225),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_267),
.A2(n_250),
.B(n_243),
.C(n_251),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_269),
.B(n_239),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_262),
.B(n_252),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_269),
.B(n_239),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_239),
.Y(n_353)
);

OR2x6_ASAP7_75t_L g354 ( 
.A(n_275),
.B(n_254),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_240),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_266),
.B(n_255),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_292),
.B(n_240),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_304),
.B(n_191),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_255),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_276),
.B(n_240),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_276),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_285),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_277),
.B(n_240),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_277),
.B(n_243),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_287),
.B(n_251),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_290),
.B(n_238),
.Y(n_372)
);

NOR2x1p5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_299),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_326),
.A2(n_216),
.B(n_236),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_334),
.A2(n_336),
.B(n_310),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_228),
.B1(n_223),
.B2(n_233),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_290),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_342),
.A2(n_236),
.B1(n_228),
.B2(n_232),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_310),
.A2(n_236),
.B1(n_192),
.B2(n_195),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_338),
.A2(n_199),
.B1(n_201),
.B2(n_197),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_236),
.B(n_228),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_323),
.A2(n_244),
.B(n_246),
.C(n_249),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_349),
.A2(n_291),
.B(n_305),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_352),
.A2(n_291),
.B(n_305),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_351),
.A2(n_236),
.B(n_228),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_298),
.B(n_293),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_306),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_316),
.B(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_327),
.B(n_293),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_223),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_330),
.A2(n_298),
.B(n_304),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_327),
.B(n_236),
.Y(n_393)
);

O2A1O1Ixp33_ASAP7_75t_SL g394 ( 
.A1(n_324),
.A2(n_233),
.B(n_224),
.C(n_231),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_328),
.A2(n_304),
.B(n_263),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_223),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_328),
.A2(n_304),
.B(n_263),
.Y(n_398)
);

OAI321xp33_ASAP7_75t_L g399 ( 
.A1(n_325),
.A2(n_215),
.A3(n_244),
.B1(n_249),
.B2(n_246),
.C(n_224),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_223),
.Y(n_400)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_308),
.B(n_165),
.Y(n_401)
);

O2A1O1Ixp5_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_249),
.B(n_246),
.C(n_231),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_363),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_355),
.A2(n_260),
.B(n_259),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_359),
.A2(n_260),
.B(n_259),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

O2A1O1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_325),
.A2(n_348),
.B(n_343),
.C(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_333),
.A2(n_232),
.B1(n_215),
.B2(n_236),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_322),
.B(n_9),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_361),
.A2(n_80),
.B(n_155),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_79),
.B(n_154),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_319),
.B(n_311),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_23),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_354),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_320),
.B(n_9),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_354),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_368),
.A2(n_82),
.B(n_153),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_313),
.A2(n_78),
.B1(n_151),
.B2(n_150),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_10),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_317),
.A2(n_76),
.B(n_149),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_354),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_318),
.A2(n_85),
.B1(n_148),
.B2(n_147),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g425 ( 
.A1(n_321),
.A2(n_75),
.B(n_142),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_337),
.A2(n_73),
.B(n_141),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_345),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_364),
.A2(n_71),
.B(n_139),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_339),
.A2(n_358),
.B(n_341),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_346),
.A2(n_70),
.B(n_137),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_347),
.A2(n_69),
.B(n_135),
.Y(n_431)
);

CKINVDCx8_ASAP7_75t_R g432 ( 
.A(n_369),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_362),
.A2(n_68),
.B(n_133),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_329),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

OAI321xp33_ASAP7_75t_L g437 ( 
.A1(n_369),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_332),
.A2(n_88),
.B(n_131),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_17),
.C(n_18),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_19),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_335),
.A2(n_356),
.B(n_350),
.Y(n_442)
);

OAI221xp5_ASAP7_75t_L g443 ( 
.A1(n_403),
.A2(n_366),
.B1(n_371),
.B2(n_364),
.C(n_309),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_388),
.A2(n_25),
.B(n_26),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_392),
.A2(n_309),
.B(n_28),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_384),
.B(n_385),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_375),
.A2(n_309),
.B(n_29),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_396),
.A2(n_309),
.B(n_31),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_387),
.A2(n_309),
.B(n_32),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_378),
.A2(n_309),
.B1(n_34),
.B2(n_35),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

AOI21x1_ASAP7_75t_L g453 ( 
.A1(n_395),
.A2(n_27),
.B(n_37),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_432),
.B(n_38),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_382),
.A2(n_40),
.B(n_43),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_374),
.A2(n_44),
.B(n_45),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_382),
.A2(n_46),
.B(n_47),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_391),
.B(n_49),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_386),
.A2(n_51),
.B(n_52),
.Y(n_460)
);

AO31x2_ASAP7_75t_L g461 ( 
.A1(n_376),
.A2(n_55),
.A3(n_57),
.B(n_58),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_389),
.B(n_60),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_374),
.A2(n_61),
.B(n_62),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_413),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_377),
.A2(n_64),
.B(n_66),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_381),
.B(n_87),
.Y(n_467)
);

AND2x6_ASAP7_75t_SL g468 ( 
.A(n_410),
.B(n_421),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_418),
.Y(n_469)
);

AOI211x1_ASAP7_75t_L g470 ( 
.A1(n_376),
.A2(n_89),
.B(n_91),
.C(n_92),
.Y(n_470)
);

AO31x2_ASAP7_75t_L g471 ( 
.A1(n_383),
.A2(n_93),
.A3(n_94),
.B(n_95),
.Y(n_471)
);

AND3x4_ASAP7_75t_L g472 ( 
.A(n_416),
.B(n_96),
.C(n_98),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_386),
.A2(n_100),
.B(n_103),
.Y(n_473)
);

AND3x4_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_107),
.C(n_108),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_390),
.B(n_109),
.Y(n_475)
);

AO31x2_ASAP7_75t_L g476 ( 
.A1(n_409),
.A2(n_110),
.A3(n_111),
.B(n_113),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_393),
.A2(n_114),
.B(n_115),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

NAND2x1_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_436),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_407),
.B(n_116),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_398),
.A2(n_117),
.B(n_118),
.Y(n_481)
);

AO31x2_ASAP7_75t_L g482 ( 
.A1(n_415),
.A2(n_119),
.A3(n_120),
.B(n_122),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_414),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_379),
.A2(n_124),
.B(n_125),
.C(n_126),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_433),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_442),
.A2(n_127),
.B(n_129),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_428),
.A2(n_157),
.B(n_405),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_404),
.A2(n_425),
.B(n_402),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_411),
.B(n_399),
.Y(n_490)
);

OA22x2_ASAP7_75t_L g491 ( 
.A1(n_423),
.A2(n_437),
.B1(n_417),
.B2(n_424),
.Y(n_491)
);

AO31x2_ASAP7_75t_L g492 ( 
.A1(n_380),
.A2(n_423),
.A3(n_422),
.B(n_430),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_440),
.A2(n_431),
.B(n_426),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_439),
.A2(n_434),
.B(n_412),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_435),
.B(n_420),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_373),
.B(n_419),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_438),
.A2(n_375),
.B(n_282),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_388),
.B(n_315),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_374),
.A2(n_310),
.B(n_375),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_381),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_392),
.A2(n_326),
.B(n_429),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_454),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_500),
.B(n_498),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_452),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_474),
.B1(n_495),
.B2(n_456),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_465),
.B(n_467),
.C(n_449),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

AOI21x1_ASAP7_75t_L g509 ( 
.A1(n_459),
.A2(n_475),
.B(n_497),
.Y(n_509)
);

AOI221x1_ASAP7_75t_L g510 ( 
.A1(n_499),
.A2(n_494),
.B1(n_490),
.B2(n_448),
.C(n_460),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_489),
.A2(n_473),
.B(n_447),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_454),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_458),
.A2(n_451),
.B1(n_444),
.B2(n_445),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_463),
.A2(n_462),
.B(n_481),
.C(n_477),
.Y(n_514)
);

AND2x6_ASAP7_75t_SL g515 ( 
.A(n_496),
.B(n_468),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_480),
.A2(n_501),
.B(n_457),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_484),
.A2(n_483),
.B(n_453),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_479),
.A2(n_487),
.B(n_466),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_486),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_455),
.B(n_485),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_472),
.A2(n_444),
.B1(n_493),
.B2(n_486),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_493),
.A2(n_470),
.B(n_443),
.Y(n_524)
);

AO31x2_ASAP7_75t_L g525 ( 
.A1(n_470),
.A2(n_461),
.A3(n_476),
.B(n_471),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_492),
.A2(n_444),
.B(n_471),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_492),
.A2(n_471),
.B(n_461),
.Y(n_527)
);

NOR2x1_ASAP7_75t_R g528 ( 
.A(n_482),
.B(n_461),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_465),
.B1(n_342),
.B2(n_310),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_476),
.A2(n_488),
.B(n_446),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_294),
.C(n_303),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_482),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_500),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_496),
.B(n_452),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_465),
.A2(n_342),
.B1(n_310),
.B2(n_495),
.Y(n_537)
);

AO31x2_ASAP7_75t_L g538 ( 
.A1(n_490),
.A2(n_376),
.A3(n_451),
.B(n_375),
.Y(n_538)
);

A2O1A1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_449),
.A2(n_342),
.B(n_458),
.C(n_456),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_454),
.Y(n_541)
);

NOR2x1_ASAP7_75t_SL g542 ( 
.A(n_478),
.B(n_310),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_488),
.A2(n_446),
.B(n_450),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_504),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_502),
.Y(n_548)
);

BUFx2_ASAP7_75t_SL g549 ( 
.A(n_506),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_506),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_505),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_535),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_540),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_540),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_505),
.B(n_507),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_544),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_544),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_539),
.A2(n_514),
.B(n_529),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_512),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_536),
.B(n_532),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_521),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_531),
.Y(n_567)
);

CKINVDCx11_ASAP7_75t_R g568 ( 
.A(n_515),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_522),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_539),
.B(n_510),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_520),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_523),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_509),
.A2(n_533),
.B(n_531),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_SL g578 ( 
.A1(n_513),
.A2(n_516),
.B(n_508),
.C(n_528),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_534),
.Y(n_579)
);

AOI221xp5_ASAP7_75t_L g580 ( 
.A1(n_513),
.A2(n_508),
.B1(n_538),
.B2(n_525),
.C(n_542),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_525),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_511),
.B(n_530),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_527),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_562),
.Y(n_588)
);

BUFx2_ASAP7_75t_SL g589 ( 
.A(n_562),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_579),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_560),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_525),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_569),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_553),
.B(n_558),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_562),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_560),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_551),
.B(n_525),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_517),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_551),
.B(n_524),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_573),
.B(n_530),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_567),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_574),
.B(n_518),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_546),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_549),
.B(n_518),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_543),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_548),
.B(n_554),
.Y(n_610)
);

AND2x4_ASAP7_75t_SL g611 ( 
.A(n_560),
.B(n_547),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_568),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_555),
.B(n_557),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_559),
.A2(n_571),
.B(n_578),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_573),
.B(n_552),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_561),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_556),
.B(n_563),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_561),
.B(n_563),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_564),
.B(n_584),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_564),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_560),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_577),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_586),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

CKINVDCx11_ASAP7_75t_R g628 ( 
.A(n_586),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_550),
.Y(n_629)
);

BUFx2_ASAP7_75t_SL g630 ( 
.A(n_550),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_583),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_627),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_583),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_627),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_604),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_580),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_572),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_604),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_617),
.B(n_575),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_593),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_606),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_594),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_587),
.B(n_552),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_602),
.B(n_601),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_587),
.B(n_572),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_606),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_603),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_590),
.B(n_618),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_625),
.B(n_582),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_588),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_626),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_609),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_618),
.B(n_582),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_552),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_614),
.B(n_585),
.Y(n_658)
);

INVx11_ASAP7_75t_L g659 ( 
.A(n_589),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_597),
.B(n_552),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_602),
.B(n_582),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_605),
.A2(n_628),
.B1(n_589),
.B2(n_598),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_634),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_646),
.B(n_609),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_634),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_661),
.B(n_654),
.Y(n_667)
);

NOR2x1_ASAP7_75t_L g668 ( 
.A(n_632),
.B(n_630),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_636),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_636),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_650),
.B(n_624),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_661),
.B(n_626),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_637),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_644),
.B(n_598),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_633),
.B(n_628),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_632),
.B(n_612),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_651),
.B(n_595),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_655),
.B(n_592),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_647),
.B(n_622),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_623),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_646),
.B(n_616),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_660),
.B(n_596),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_655),
.B(n_607),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_637),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_631),
.B(n_613),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_647),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_647),
.B(n_649),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_642),
.B(n_610),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_642),
.B(n_610),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_662),
.B(n_599),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_652),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_666),
.Y(n_694)
);

NOR2x1p5_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_612),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_664),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_687),
.B(n_688),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_666),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_669),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_687),
.B(n_647),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_663),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_667),
.B(n_631),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_663),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_669),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_670),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_670),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_691),
.A2(n_675),
.B1(n_638),
.B2(n_676),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_667),
.B(n_635),
.Y(n_708)
);

AND2x4_ASAP7_75t_SL g709 ( 
.A(n_679),
.B(n_645),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_673),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_635),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_690),
.B(n_641),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_673),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

AOI21xp33_ASAP7_75t_SL g715 ( 
.A1(n_707),
.A2(n_675),
.B(n_674),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_707),
.A2(n_679),
.B1(n_645),
.B2(n_688),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_R g717 ( 
.A(n_700),
.B(n_664),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_706),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_706),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_694),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_698),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_695),
.A2(n_679),
.B1(n_645),
.B2(n_688),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_712),
.B(n_665),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_711),
.B(n_665),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_696),
.A2(n_659),
.B1(n_668),
.B2(n_671),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_716),
.B(n_697),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_SL g727 ( 
.A(n_725),
.B(n_680),
.C(n_682),
.Y(n_727)
);

OAI222xp33_ASAP7_75t_L g728 ( 
.A1(n_725),
.A2(n_692),
.B1(n_696),
.B2(n_708),
.C1(n_702),
.C2(n_700),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_677),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_715),
.A2(n_709),
.B(n_700),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_718),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_SL g732 ( 
.A1(n_717),
.A2(n_714),
.B(n_713),
.C(n_710),
.Y(n_732)
);

AOI221x1_ASAP7_75t_SL g733 ( 
.A1(n_726),
.A2(n_720),
.B1(n_721),
.B2(n_719),
.C(n_704),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_730),
.A2(n_723),
.B1(n_724),
.B2(n_652),
.Y(n_734)
);

AOI222xp33_ASAP7_75t_L g735 ( 
.A1(n_728),
.A2(n_677),
.B1(n_678),
.B2(n_683),
.C1(n_699),
.C2(n_705),
.Y(n_735)
);

AOI311xp33_ASAP7_75t_L g736 ( 
.A1(n_732),
.A2(n_727),
.A3(n_684),
.B(n_693),
.C(n_653),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_726),
.B(n_681),
.Y(n_737)
);

AOI211xp5_ASAP7_75t_SL g738 ( 
.A1(n_729),
.A2(n_681),
.B(n_697),
.C(n_639),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_734),
.B(n_731),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_738),
.A2(n_697),
.B(n_709),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_733),
.B(n_678),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_737),
.Y(n_742)
);

NOR3xp33_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_736),
.C(n_629),
.Y(n_743)
);

AOI211xp5_ASAP7_75t_L g744 ( 
.A1(n_741),
.A2(n_735),
.B(n_703),
.C(n_701),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_743),
.B(n_742),
.C(n_740),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_744),
.Y(n_746)
);

NAND4xp75_ASAP7_75t_L g747 ( 
.A(n_743),
.B(n_608),
.C(n_629),
.D(n_659),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_746),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_745),
.B(n_685),
.Y(n_749)
);

XNOR2xp5_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_611),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_746),
.B(n_703),
.Y(n_751)
);

XNOR2xp5_ASAP7_75t_L g752 ( 
.A(n_745),
.B(n_611),
.Y(n_752)
);

NAND2x1_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_701),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_753),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_748),
.A2(n_683),
.B1(n_686),
.B2(n_653),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_752),
.Y(n_756)
);

OAI221xp5_ASAP7_75t_L g757 ( 
.A1(n_750),
.A2(n_658),
.B1(n_686),
.B2(n_648),
.C(n_643),
.Y(n_757)
);

OAI222xp33_ASAP7_75t_L g758 ( 
.A1(n_749),
.A2(n_658),
.B1(n_621),
.B2(n_599),
.C1(n_591),
.C2(n_648),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_751),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_759),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_754),
.Y(n_761)
);

OAI22x1_ASAP7_75t_L g762 ( 
.A1(n_756),
.A2(n_591),
.B1(n_621),
.B2(n_599),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_755),
.B(n_685),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_761),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_757),
.B1(n_758),
.B2(n_658),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_763),
.B(n_672),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_762),
.B(n_640),
.Y(n_767)
);

XOR2x1_ASAP7_75t_L g768 ( 
.A(n_766),
.B(n_549),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_765),
.B(n_672),
.Y(n_769)
);

XNOR2xp5_ASAP7_75t_L g770 ( 
.A(n_768),
.B(n_630),
.Y(n_770)
);

OAI221xp5_ASAP7_75t_L g771 ( 
.A1(n_769),
.A2(n_591),
.B1(n_599),
.B2(n_621),
.C(n_658),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_767),
.B(n_643),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_772),
.B(n_771),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_615),
.B1(n_621),
.B2(n_599),
.Y(n_774)
);


endmodule