module fake_jpeg_8070_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_17),
.B1(n_15),
.B2(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_40),
.B1(n_25),
.B2(n_13),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_29),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_12),
.B1(n_19),
.B2(n_11),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_36),
.C(n_31),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.C(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_47),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_22),
.B(n_13),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_11),
.B2(n_4),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_13),
.Y(n_50)
);

XOR2x1_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_21),
.B1(n_5),
.B2(n_3),
.Y(n_68)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_70),
.C(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_21),
.A3(n_37),
.B1(n_7),
.B2(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_51),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_47),
.B(n_48),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_81),
.B(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_60),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_45),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.C(n_66),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_67),
.B(n_63),
.C(n_62),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_79),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_87),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_80),
.A2(n_41),
.B1(n_56),
.B2(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_59),
.B1(n_64),
.B2(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_78),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_83),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_78),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_84),
.B(n_85),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_100),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.C(n_101),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_7),
.B(n_5),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_107),
.Y(n_109)
);


endmodule