module fake_jpeg_21072_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_1),
.C(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_31),
.Y(n_52)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_16),
.B1(n_33),
.B2(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_49),
.A2(n_29),
.B1(n_28),
.B2(n_0),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_51),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_20),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_23),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_68),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_19),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_30),
.B1(n_18),
.B2(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_65),
.B1(n_8),
.B2(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_27),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_24),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_75),
.B1(n_55),
.B2(n_48),
.Y(n_116)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_108),
.B1(n_93),
.B2(n_62),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_106),
.B1(n_56),
.B2(n_55),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_8),
.B1(n_2),
.B2(n_4),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_58),
.B1(n_66),
.B2(n_48),
.Y(n_118)
);

AO22x2_ASAP7_75t_SL g108 ( 
.A1(n_49),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_78),
.B1(n_80),
.B2(n_53),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_114),
.B1(n_120),
.B2(n_135),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_78),
.B1(n_53),
.B2(n_75),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_95),
.C(n_92),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_138),
.B1(n_93),
.B2(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_75),
.B1(n_62),
.B2(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_130),
.Y(n_157)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_128),
.B(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_73),
.B1(n_72),
.B2(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_50),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_61),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_59),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_97),
.B(n_6),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_150),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_100),
.C(n_94),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_90),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_156),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_85),
.B1(n_82),
.B2(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_158),
.B1(n_133),
.B2(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_60),
.B1(n_67),
.B2(n_10),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_124),
.B1(n_123),
.B2(n_138),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_137),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_178),
.B1(n_160),
.B2(n_142),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_143),
.B(n_163),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_124),
.B(n_120),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_177),
.B(n_179),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_127),
.B(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_118),
.B1(n_114),
.B2(n_110),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_125),
.B(n_131),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_136),
.B(n_9),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_157),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_189),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_150),
.C(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_195),
.C(n_141),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_162),
.B(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

OAI321xp33_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_166),
.A3(n_173),
.B1(n_176),
.B2(n_167),
.C(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_167),
.B1(n_178),
.B2(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_174),
.B1(n_141),
.B2(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_151),
.C(n_154),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_177),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_206),
.C(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_165),
.C(n_161),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_192),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_192),
.B(n_188),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_186),
.A3(n_184),
.B(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_204),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_224),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_225),
.B(n_213),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_216),
.B(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_203),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_220),
.C(n_222),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_233),
.B(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_202),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_234),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_199),
.B(n_191),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_237),
.B(n_7),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_185),
.C(n_9),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);


endmodule