module fake_jpeg_12617_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_33),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_38),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_26),
.B1(n_20),
.B2(n_30),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_80),
.A2(n_82),
.B(n_89),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_30),
.B1(n_23),
.B2(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_36),
.B1(n_23),
.B2(n_30),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_43),
.B1(n_42),
.B2(n_24),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_26),
.C(n_17),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_29),
.B1(n_27),
.B2(n_34),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_51),
.B1(n_27),
.B2(n_17),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_31),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_31),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_59),
.Y(n_131)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_71),
.B1(n_72),
.B2(n_49),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_75),
.B1(n_89),
.B2(n_80),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_102),
.B1(n_110),
.B2(n_94),
.Y(n_164)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_123),
.Y(n_180)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_64),
.B1(n_55),
.B2(n_73),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_126),
.A2(n_127),
.B1(n_147),
.B2(n_155),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_44),
.B1(n_24),
.B2(n_17),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_63),
.B1(n_58),
.B2(n_53),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_139),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_41),
.B1(n_50),
.B2(n_48),
.Y(n_133)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_102),
.B1(n_74),
.B2(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_76),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_59),
.B1(n_24),
.B2(n_37),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_81),
.B(n_19),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_1),
.Y(n_171)
);

AND2x4_ASAP7_75t_SL g151 ( 
.A(n_79),
.B(n_85),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_106),
.C(n_37),
.Y(n_188)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_19),
.A3(n_104),
.B1(n_96),
.B2(n_78),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_134),
.B(n_116),
.C(n_149),
.D(n_123),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_162),
.B1(n_173),
.B2(n_190),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_112),
.B1(n_74),
.B2(n_94),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_117),
.B1(n_129),
.B2(n_131),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_171),
.B(n_2),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_106),
.B1(n_99),
.B2(n_98),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_37),
.C(n_19),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_179),
.C(n_35),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_37),
.Y(n_179)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_136),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_140),
.A2(n_98),
.B1(n_88),
.B2(n_35),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_19),
.B(n_35),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_156),
.B(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_141),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_194),
.B(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_146),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_196),
.B(n_204),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_222),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_192),
.B1(n_187),
.B2(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_203),
.B1(n_209),
.B2(n_210),
.Y(n_238)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_144),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_191),
.C(n_170),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_118),
.B1(n_130),
.B2(n_133),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_135),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_124),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_151),
.B1(n_152),
.B2(n_147),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_212),
.B1(n_215),
.B2(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_151),
.B1(n_147),
.B2(n_120),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_147),
.B1(n_151),
.B2(n_128),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_216),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_137),
.B1(n_125),
.B2(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_214),
.A2(n_221),
.B(n_225),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_153),
.B1(n_123),
.B2(n_155),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_219),
.Y(n_247)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_115),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_223),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_157),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_230),
.B1(n_180),
.B2(n_169),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_172),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_174),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_156),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_9),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_264),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_182),
.B1(n_183),
.B2(n_180),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_248),
.B1(n_218),
.B2(n_207),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_191),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_241),
.A2(n_257),
.B1(n_231),
.B2(n_207),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_246),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_200),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_183),
.B1(n_172),
.B2(n_167),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_250),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_214),
.B(n_202),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_251),
.A2(n_10),
.B(n_11),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_170),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_169),
.B(n_167),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_185),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_259),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_198),
.A2(n_184),
.B1(n_7),
.B2(n_8),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_212),
.B(n_184),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_221),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_263),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_195),
.B(n_6),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_286),
.B1(n_291),
.B2(n_265),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_274),
.C(n_276),
.Y(n_305)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_208),
.C(n_213),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_233),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_223),
.C(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_224),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_284),
.C(n_294),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_203),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_232),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_238),
.A2(n_199),
.B1(n_230),
.B2(n_227),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_290),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_199),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_295),
.B(n_266),
.Y(n_300)
);

AO22x2_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_264),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_10),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_238),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_302),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_266),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_297),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_300),
.A2(n_304),
.B(n_290),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_301),
.B(n_288),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_266),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_266),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_267),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_240),
.B(n_257),
.C(n_242),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_260),
.B1(n_232),
.B2(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_260),
.B1(n_252),
.B2(n_247),
.Y(n_309)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_256),
.C(n_240),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_292),
.C(n_283),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_284),
.B(n_289),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_317),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_SL g317 ( 
.A(n_274),
.B(n_241),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_279),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_320),
.B1(n_319),
.B2(n_316),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_330),
.C(n_333),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_292),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_328),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_340),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_267),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_294),
.C(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_306),
.B(n_250),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_308),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_282),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_282),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_311),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_287),
.C(n_278),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_317),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_297),
.B(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_338),
.A2(n_313),
.B1(n_297),
.B2(n_300),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_343),
.A2(n_353),
.B1(n_357),
.B2(n_304),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_341),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_346),
.B(n_352),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_339),
.A2(n_313),
.B1(n_332),
.B2(n_321),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_348),
.A2(n_355),
.B1(n_326),
.B2(n_337),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_354),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_336),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_310),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_356),
.A2(n_330),
.B(n_315),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_318),
.B1(n_304),
.B2(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_323),
.C(n_325),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_362),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_367),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_323),
.C(n_340),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_342),
.B1(n_324),
.B2(n_304),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_334),
.C(n_333),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_347),
.C(n_362),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_366),
.B(n_370),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_327),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_327),
.B1(n_262),
.B2(n_245),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_351),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_357),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_360),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_368),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_378),
.B(n_368),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_361),
.A2(n_356),
.B(n_347),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_380),
.A2(n_381),
.B(n_370),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_350),
.B(n_245),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_382),
.B(n_384),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_385),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_358),
.Y(n_384)
);

OAI321xp33_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_366),
.A3(n_359),
.B1(n_258),
.B2(n_236),
.C(n_290),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_372),
.C(n_377),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_379),
.B(n_258),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_388),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_373),
.A2(n_236),
.B1(n_263),
.B2(n_246),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_376),
.A2(n_367),
.B1(n_243),
.B2(n_244),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_244),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_394),
.B(n_390),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_382),
.A2(n_377),
.B(n_243),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_384),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_397),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_398),
.A2(n_399),
.B(n_400),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_243),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_243),
.B(n_290),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_393),
.Y(n_403)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_403),
.A2(n_401),
.B(n_394),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_290),
.C(n_13),
.Y(n_405)
);

AOI31xp33_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_13),
.B(n_260),
.Y(n_407)
);


endmodule