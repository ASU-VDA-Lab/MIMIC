module fake_jpeg_17878_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_47),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_1),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_23),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_16),
.B1(n_34),
.B2(n_32),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_16),
.B1(n_23),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_76),
.B1(n_4),
.B2(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_77),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_32),
.B1(n_25),
.B2(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_28),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_31),
.C(n_27),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_28),
.B(n_31),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_12),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_105),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_93),
.Y(n_118)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_98),
.Y(n_119)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_58),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_79),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_124),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_70),
.B1(n_71),
.B2(n_68),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_111),
.B(n_114),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_99),
.B1(n_94),
.B2(n_63),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_95),
.B(n_85),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_64),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_80),
.C(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_75),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_65),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_105),
.B1(n_74),
.B2(n_63),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_136),
.B1(n_119),
.B2(n_121),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_138),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_53),
.B(n_69),
.C(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_90),
.B1(n_103),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_140),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_135),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_54),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_121),
.C(n_124),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_152),
.B1(n_132),
.B2(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_127),
.C(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_127),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_164),
.C(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_153),
.B1(n_123),
.B2(n_151),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_144),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_163),
.B(n_161),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_146),
.B1(n_156),
.B2(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_173),
.C(n_159),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_158),
.B(n_157),
.Y(n_184)
);

OAI31xp33_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_178),
.A3(n_171),
.B(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_180),
.C(n_140),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_176),
.A3(n_160),
.B1(n_157),
.B2(n_164),
.C1(n_161),
.C2(n_54),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_185),
.B(n_181),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_13),
.B(n_14),
.Y(n_190)
);


endmodule