module fake_jpeg_9394_n_114 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_23),
.B1(n_22),
.B2(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_48),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_40),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_23),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_65),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_61),
.B(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_39),
.B1(n_29),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_47),
.B1(n_39),
.B2(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_53),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_42),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_36),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_13),
.C(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_71),
.B(n_73),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_45),
.B1(n_24),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_75),
.B1(n_63),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_44),
.B1(n_43),
.B2(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_57),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_18),
.B1(n_12),
.B2(n_27),
.C(n_30),
.Y(n_82)
);

OAI322xp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_9),
.A3(n_3),
.B1(n_4),
.B2(n_7),
.C1(n_8),
.C2(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_71),
.A3(n_74),
.B1(n_77),
.B2(n_73),
.C1(n_31),
.C2(n_27),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_78),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_8),
.A3(n_9),
.B1(n_2),
.B2(n_0),
.C(n_1),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_83),
.C(n_94),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.C(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_49),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_91),
.B1(n_62),
.B2(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_96),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_107),
.C(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_102),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_2),
.Y(n_112)
);

OAI21x1_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_2),
.B(n_110),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_28),
.Y(n_114)
);


endmodule