module fake_jpeg_28502_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_59),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_70),
.B1(n_54),
.B2(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_80),
.B1(n_64),
.B2(n_24),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_65),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_6),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_49),
.B1(n_56),
.B2(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_66),
.B(n_51),
.C(n_50),
.Y(n_91)
);

NOR2x1_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_66),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_26),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_60),
.B1(n_48),
.B2(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_100),
.B1(n_79),
.B2(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_101),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_4),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_9),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_111),
.B1(n_118),
.B2(n_121),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_7),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_112),
.B1(n_113),
.B2(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_30),
.C(n_44),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_10),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NOR4xp25_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_25),
.C(n_43),
.D(n_41),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_14),
.B(n_18),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_140),
.B1(n_136),
.B2(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_147),
.B1(n_23),
.B2(n_31),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_19),
.B(n_21),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_132),
.C(n_34),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_128),
.C(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_150),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_137),
.B1(n_129),
.B2(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_149),
.C(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_146),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_142),
.B(n_152),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_146),
.A3(n_145),
.B1(n_141),
.B2(n_153),
.C(n_32),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_36),
.CI(n_38),
.CON(n_162),
.SN(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_40),
.Y(n_163)
);


endmodule