module fake_jpeg_19011_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_0),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_1),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_47),
.B1(n_49),
.B2(n_60),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_63),
.B1(n_39),
.B2(n_61),
.Y(n_80)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_68),
.B1(n_56),
.B2(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_51),
.B1(n_62),
.B2(n_40),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_79),
.B1(n_48),
.B2(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_51),
.B1(n_44),
.B2(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_54),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_88),
.B(n_10),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_23),
.B1(n_34),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_58),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_74),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_103),
.B(n_30),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_101),
.B1(n_28),
.B2(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_14),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_93),
.B1(n_97),
.B2(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_108),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_97),
.C(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_110),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_109),
.Y(n_129)
);


endmodule