module fake_jpeg_27698_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_55),
.B1(n_23),
.B2(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_16),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_0),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_69),
.B1(n_22),
.B2(n_33),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_32),
.B1(n_24),
.B2(n_23),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_0),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_74),
.Y(n_108)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_76),
.Y(n_128)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_83),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_102),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_90),
.B1(n_93),
.B2(n_19),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_76),
.B1(n_77),
.B2(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_98),
.B1(n_19),
.B2(n_20),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_33),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_64),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_68),
.B1(n_70),
.B2(n_57),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_118),
.B1(n_119),
.B2(n_127),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_61),
.B1(n_53),
.B2(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_74),
.B1(n_71),
.B2(n_99),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_56),
.B1(n_63),
.B2(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_125),
.B1(n_132),
.B2(n_101),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_53),
.B1(n_50),
.B2(n_49),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_33),
.B1(n_26),
.B2(n_20),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_0),
.B(n_1),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_26),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_96),
.B1(n_84),
.B2(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_81),
.C(n_73),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_143),
.C(n_155),
.Y(n_168)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_161),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_100),
.B(n_103),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_165),
.B(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_85),
.C(n_104),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_78),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_141),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_151),
.B1(n_25),
.B2(n_18),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_98),
.B(n_88),
.C(n_79),
.D(n_74),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_149),
.B(n_25),
.C(n_14),
.Y(n_195)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_105),
.B1(n_125),
.B2(n_115),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_79),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_97),
.C(n_92),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_163),
.Y(n_197)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_164),
.B1(n_127),
.B2(n_119),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_71),
.B1(n_25),
.B2(n_18),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_112),
.B1(n_121),
.B2(n_113),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_107),
.C(n_131),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_182),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_191),
.B1(n_166),
.B2(n_148),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_186),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_196),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_116),
.B1(n_114),
.B2(n_121),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_192),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_157),
.A2(n_113),
.B1(n_107),
.B2(n_109),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_106),
.B1(n_123),
.B2(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_130),
.C(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_177),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_178),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_140),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_194),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_25),
.B1(n_18),
.B2(n_97),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_198),
.B1(n_199),
.B2(n_134),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_97),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_200),
.C(n_2),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_25),
.B1(n_14),
.B2(n_13),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_136),
.A2(n_142),
.B1(n_138),
.B2(n_141),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_12),
.C(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_209),
.B1(n_221),
.B2(n_188),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_165),
.B(n_138),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_216),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_215),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_230),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_158),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_3),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_4),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_199),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_168),
.C(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_249),
.C(n_219),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_214),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_235),
.B(n_209),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_168),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_245),
.B1(n_252),
.B2(n_229),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_182),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_243),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_169),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_191),
.B1(n_193),
.B2(n_171),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_187),
.C(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_173),
.B1(n_5),
.B2(n_6),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_259),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_211),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_215),
.C(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_272),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_263),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_213),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_205),
.B1(n_245),
.B2(n_233),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_217),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_275),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_210),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_203),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_274),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_227),
.C(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_217),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_218),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_243),
.C(n_240),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_286),
.C(n_264),
.Y(n_292)
);

OAI322xp33_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_246),
.A3(n_249),
.B1(n_251),
.B2(n_248),
.C1(n_238),
.C2(n_247),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_222),
.B(n_273),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_236),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_260),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_254),
.C(n_202),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_259),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_252),
.B1(n_211),
.B2(n_221),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_228),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_299),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_297),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_264),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_300),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_260),
.C(n_228),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.C(n_277),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_4),
.C(n_5),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_284),
.A2(n_5),
.B(n_6),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_6),
.B(n_7),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_5),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_276),
.B(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_285),
.CI(n_277),
.CON(n_308),
.SN(n_308)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_301),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_303),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_296),
.B(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_317),
.B(n_323),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_324),
.B(n_312),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_328),
.C(n_321),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g327 ( 
.A(n_319),
.B(n_290),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_299),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_318),
.C(n_311),
.Y(n_333)
);

AOI321xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_315),
.C(n_327),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_8),
.B(n_9),
.Y(n_336)
);


endmodule