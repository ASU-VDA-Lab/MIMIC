module fake_jpeg_2090_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_58),
.B1(n_53),
.B2(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_79),
.B1(n_51),
.B2(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_53),
.B1(n_61),
.B2(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_82),
.B1(n_69),
.B2(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_54),
.B1(n_49),
.B2(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_46),
.B1(n_55),
.B2(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_86),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_49),
.B(n_57),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_98),
.B(n_81),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_83),
.B1(n_81),
.B2(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_57),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_35),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_7),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_83),
.B1(n_44),
.B2(n_41),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_121),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_36),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_128),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_97),
.B(n_34),
.C(n_32),
.D(n_31),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_133),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_6),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_29),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_R g148 ( 
.A(n_134),
.B(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_7),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_140),
.B(n_110),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_18),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_9),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_110),
.B(n_114),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_112),
.C(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_134),
.C(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_115),
.A3(n_110),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_9),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_154),
.A3(n_153),
.B1(n_126),
.B2(n_144),
.C1(n_155),
.C2(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_128),
.C(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_140),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_122),
.B(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_160),
.B1(n_151),
.B2(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_157),
.B1(n_127),
.B2(n_12),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_166),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_147),
.C(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_163),
.C(n_165),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_10),
.B(n_11),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_10),
.B(n_13),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_14),
.B(n_15),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_16),
.Y(n_175)
);


endmodule