module real_jpeg_143_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_40),
.B1(n_69),
.B2(n_70),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_1),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_69),
.B1(n_70),
.B2(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_164),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_2),
.A2(n_34),
.B1(n_41),
.B2(n_164),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_69),
.B1(n_70),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_34),
.B1(n_41),
.B2(n_80),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_34),
.B1(n_41),
.B2(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_6),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_46),
.B1(n_48),
.B2(n_74),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_74),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_8),
.A2(n_69),
.B1(n_70),
.B2(n_130),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_8),
.A2(n_46),
.B1(n_48),
.B2(n_130),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_8),
.A2(n_34),
.B1(n_41),
.B2(n_130),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_69),
.B1(n_70),
.B2(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_46),
.B1(n_48),
.B2(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_9),
.A2(n_34),
.B1(n_41),
.B2(n_184),
.Y(n_263)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_10),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_45),
.B1(n_69),
.B2(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_11),
.A2(n_45),
.B1(n_62),
.B2(n_63),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_11),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_329),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_15),
.B(n_330),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_16),
.A2(n_62),
.B1(n_63),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_16),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_16),
.A2(n_46),
.B1(n_48),
.B2(n_72),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_16),
.A2(n_34),
.B1(n_41),
.B2(n_72),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_18),
.B(n_62),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_18),
.B(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_18),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_18),
.A2(n_62),
.B(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_18),
.B(n_83),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_18),
.A2(n_70),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_18),
.B(n_34),
.C(n_51),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_18),
.A2(n_46),
.B1(n_48),
.B2(n_210),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_18),
.B(n_37),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_18),
.B(n_56),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_324),
.B(n_327),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_316),
.B(n_320),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_303),
.B(n_315),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_144),
.B(n_300),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_131),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_104),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_27),
.B(n_104),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_75),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_90),
.C(n_102),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_57),
.B(n_58),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_29),
.A2(n_30),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_31),
.A2(n_57),
.B1(n_58),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_31),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_38),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_32),
.A2(n_36),
.B1(n_118),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_32),
.A2(n_36),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_32),
.A2(n_36),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_37),
.B1(n_39),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_33),
.A2(n_37),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_33),
.A2(n_37),
.B1(n_177),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_33),
.A2(n_37),
.B1(n_214),
.B2(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_33),
.A2(n_37),
.B1(n_210),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_33),
.A2(n_37),
.B1(n_263),
.B2(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_34),
.B(n_261),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_44),
.A2(n_49),
.B1(n_56),
.B2(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AO22x2_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_48),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_46),
.A2(n_70),
.A3(n_84),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_46),
.B(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_48),
.B(n_85),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_56),
.B(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_49),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_49),
.A2(n_56),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_49),
.A2(n_56),
.B1(n_206),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_49),
.A2(n_56),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_49),
.A2(n_56),
.B1(n_233),
.B2(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_53),
.A2(n_122),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_53),
.A2(n_157),
.B1(n_205),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_68),
.B1(n_73),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_68),
.B1(n_71),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_59),
.A2(n_68),
.B1(n_93),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_59),
.A2(n_68),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_59),
.A2(n_68),
.B1(n_183),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_129),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_60),
.A2(n_165),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_60),
.A2(n_165),
.B1(n_311),
.B2(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_60),
.A2(n_165),
.B(n_318),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_63),
.A2(n_67),
.A3(n_70),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_65),
.B(n_69),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_69),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_70),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_69),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_90),
.B1(n_102),
.B2(n_103),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_77),
.B(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_83),
.B2(n_87),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_79),
.A2(n_82),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_83),
.B1(n_87),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_81),
.A2(n_83),
.B1(n_125),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_81),
.A2(n_83),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_82),
.A2(n_100),
.B1(n_126),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_82),
.A2(n_126),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_82),
.A2(n_126),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_82),
.A2(n_126),
.B1(n_180),
.B2(n_196),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_82),
.A2(n_126),
.B1(n_195),
.B2(n_242),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_92),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_96),
.C(n_98),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_92),
.B(n_135),
.C(n_142),
.Y(n_304)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_101),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_101),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_96),
.B(n_138),
.C(n_140),
.Y(n_314)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_112),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.C(n_127),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_114),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_127),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_131),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_143),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_132),
.B(n_143),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_139),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_166),
.B(n_299),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_146),
.B(n_148),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.C(n_162),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_155),
.B(n_158),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_189),
.B(n_298),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_187),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_168),
.B(n_187),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_186),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_169),
.B(n_186),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_171),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.C(n_182),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_172),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_176),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_179),
.B(n_182),
.Y(n_289)
);

AOI31xp33_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_283),
.A3(n_292),
.B(n_295),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_228),
.B(n_282),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_216),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_216),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.C(n_207),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_198),
.C(n_202),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_203),
.B(n_207),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_212),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_216),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_216),
.B(n_293),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.CI(n_219),
.CON(n_216),
.SN(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_220),
.B(n_223),
.C(n_227),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_277),
.B(n_281),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_246),
.B(n_276),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_238),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_235),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_241),
.C(n_244),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_257),
.B(n_275),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_269),
.B(n_274),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_264),
.B(n_268),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_287),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_314),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_312),
.C(n_314),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_326),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule