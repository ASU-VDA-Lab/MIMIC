module fake_netlist_6_2708_n_1349 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1349);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1349;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_934;
wire n_482;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_367;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_924;
wire n_475;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g314 ( 
.A(n_115),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_203),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_309),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_299),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_304),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_128),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_93),
.Y(n_320)
);

INVxp33_ASAP7_75t_R g321 ( 
.A(n_188),
.Y(n_321)
);

BUFx8_ASAP7_75t_SL g322 ( 
.A(n_118),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_3),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_207),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_254),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_6),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_25),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_303),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_164),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_31),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_236),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_112),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_154),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_87),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_42),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_91),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_51),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_72),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_177),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_217),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_256),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_313),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_119),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_121),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_278),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_34),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_284),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_101),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_148),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_182),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_184),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_262),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_127),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_25),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_2),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_135),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_116),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_263),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_73),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_28),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_186),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_194),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_287),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_21),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_51),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_168),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_84),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_10),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_155),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_296),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_32),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_69),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_291),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_143),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_125),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_52),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_80),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_179),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_159),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_132),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_24),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_28),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_131),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_150),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_153),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_61),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_208),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_221),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_123),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_114),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_266),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_139),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_204),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_76),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_307),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_152),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_48),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_3),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_250),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_124),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_41),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_103),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_228),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_292),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_122),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_27),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_197),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_231),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_218),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_26),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_175),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_180),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_88),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_9),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_35),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_170),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_295),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_7),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_202),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_297),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_183),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_270),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_11),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_141),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_288),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_172),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_289),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_308),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_41),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_243),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_16),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_29),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_126),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_239),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_36),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_100),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_86),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_78),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_310),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_17),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_111),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_42),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_268),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_162),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_94),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_57),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_96),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_196),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_166),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_260),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_201),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_290),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_20),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_301),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_20),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_233),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_157),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_265),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_209),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_7),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_187),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_32),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_113),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_271),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_235),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_220),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_305),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_189),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_130),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_225),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_158),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_190),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_258),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_181),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_302),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_108),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_229),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_275),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_264),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_95),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_133),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_63),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_312),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_322),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_405),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_356),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_331),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_315),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_384),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_359),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_395),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_359),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_360),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_323),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_0),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_316),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_363),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_317),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_359),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_448),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_397),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_368),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_327),
.B(n_0),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_360),
.Y(n_515)
);

INVxp33_ASAP7_75t_SL g516 ( 
.A(n_326),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_371),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_371),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_314),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_359),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_353),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_318),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_319),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_400),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_333),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_320),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_372),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_346),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_364),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_365),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_324),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_376),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_325),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_328),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_377),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_382),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_468),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_329),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_447),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_386),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_431),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_348),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_332),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g544 ( 
.A(n_327),
.B(n_1),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_334),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_375),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_336),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_339),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_391),
.B(n_1),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_393),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_340),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_335),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_401),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_359),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_380),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_379),
.B(n_2),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_416),
.B(n_4),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_331),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_413),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_342),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_424),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_338),
.B(n_4),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_450),
.B(n_5),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_338),
.B(n_5),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_344),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_345),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_389),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_347),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_349),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_357),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_350),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_341),
.B(n_6),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_351),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_474),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_369),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_354),
.B(n_8),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_352),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_355),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_477),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_495),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_519),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_505),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_542),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_560),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_574),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_337),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_507),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_525),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_539),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_542),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_528),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_529),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_510),
.B(n_406),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_362),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_557),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_504),
.B(n_388),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_504),
.B(n_388),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_522),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_496),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_535),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_574),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_574),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_506),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_536),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_502),
.B(n_337),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_523),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_540),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_558),
.B(n_388),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_526),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_531),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_533),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_498),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_534),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_502),
.B(n_343),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_538),
.B(n_429),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_553),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_555),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_500),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_561),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_558),
.B(n_412),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_500),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_509),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_543),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_508),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_508),
.A2(n_452),
.B(n_412),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_545),
.B(n_441),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_548),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_563),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_565),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_551),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_583),
.A2(n_330),
.B1(n_402),
.B2(n_385),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_343),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_564),
.B(n_478),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_572),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_573),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_516),
.B(n_480),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_512),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_521),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_585),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_588),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_559),
.B(n_392),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_580),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_513),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_524),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_586),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_515),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_490),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_520),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_554),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_489),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_537),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_671),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_625),
.B(n_554),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_672),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_590),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_593),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_552),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_617),
.B(n_628),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_595),
.B(n_511),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_589),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_651),
.B(n_527),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_605),
.B(n_560),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_597),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_625),
.B(n_517),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_594),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_600),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_636),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_671),
.Y(n_691)
);

INVx8_ASAP7_75t_L g692 ( 
.A(n_669),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_668),
.B(n_518),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_594),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_604),
.B(n_546),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_671),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_671),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_632),
.B(n_359),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_603),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_591),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_606),
.B(n_494),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_604),
.B(n_499),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_642),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_659),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_620),
.B(n_492),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_629),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_613),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_612),
.Y(n_711)
);

INVxp33_ASAP7_75t_L g712 ( 
.A(n_650),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_607),
.B(n_501),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_619),
.Y(n_715)
);

INVx6_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_621),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_604),
.B(n_452),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_596),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_620),
.B(n_547),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_514),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_659),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_637),
.B(n_549),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_631),
.B(n_389),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_633),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_653),
.B(n_571),
.Y(n_726)
);

AND2x2_ASAP7_75t_SL g727 ( 
.A(n_637),
.B(n_559),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_613),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_666),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_644),
.B(n_549),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_635),
.B(n_544),
.Y(n_731)
);

CKINVDCx11_ASAP7_75t_R g732 ( 
.A(n_592),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_614),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_614),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_643),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_607),
.B(n_579),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_632),
.B(n_359),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_608),
.B(n_584),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_567),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_663),
.B(n_321),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_646),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_634),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_647),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_648),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_663),
.B(n_575),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_609),
.B(n_576),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_652),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_634),
.B(n_484),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_618),
.B(n_578),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_622),
.B(n_587),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_655),
.B(n_486),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_602),
.A2(n_567),
.B1(n_583),
.B2(n_411),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_623),
.B(n_392),
.Y(n_753)
);

INVx6_ASAP7_75t_L g754 ( 
.A(n_598),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_660),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_662),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_638),
.B(n_487),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_642),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_666),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_638),
.B(n_389),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_602),
.B(n_403),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_624),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_742),
.Y(n_764)
);

NAND2x1_ASAP7_75t_L g765 ( 
.A(n_674),
.B(n_641),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_747),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_708),
.A2(n_569),
.B(n_566),
.C(n_658),
.Y(n_767)
);

OAI221xp5_ASAP7_75t_L g768 ( 
.A1(n_723),
.A2(n_419),
.B1(n_406),
.B2(n_658),
.C(n_420),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_692),
.B(n_716),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_688),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_727),
.A2(n_419),
.B1(n_423),
.B2(n_415),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_719),
.B(n_627),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_730),
.B(n_641),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_685),
.B(n_640),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_736),
.A2(n_670),
.B1(n_656),
.B2(n_426),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_718),
.B(n_656),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_696),
.B(n_645),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_718),
.B(n_670),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_695),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_677),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_707),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_680),
.A2(n_654),
.B1(n_664),
.B2(n_649),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_678),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_709),
.B(n_681),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_686),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_675),
.A2(n_426),
.B(n_389),
.Y(n_786)
);

NOR3x1_ASAP7_75t_L g787 ( 
.A(n_682),
.B(n_493),
.C(n_434),
.Y(n_787)
);

AND2x4_ASAP7_75t_SL g788 ( 
.A(n_719),
.B(n_610),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_707),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_718),
.B(n_667),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_718),
.B(n_358),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_738),
.B(n_361),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_759),
.B(n_366),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_703),
.B(n_739),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_684),
.B(n_673),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_675),
.B(n_426),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_705),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_712),
.A2(n_426),
.B1(n_432),
.B2(n_392),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_716),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_743),
.B(n_367),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_710),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_748),
.B(n_432),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_762),
.B(n_493),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_747),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_734),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_763),
.B(n_370),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_748),
.B(n_432),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_693),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_714),
.A2(n_758),
.B(n_694),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_758),
.B(n_432),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_687),
.B(n_373),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_687),
.B(n_374),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_700),
.B(n_378),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_713),
.B(n_381),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_721),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_741),
.B(n_673),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_689),
.B(n_383),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_683),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_720),
.B(n_610),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_715),
.B(n_390),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_725),
.B(n_394),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_744),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_755),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_756),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_745),
.A2(n_398),
.B1(n_399),
.B2(n_396),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_757),
.B(n_408),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_721),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_676),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_674),
.B(n_691),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_735),
.B(n_409),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_691),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_698),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_702),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_706),
.B(n_428),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_711),
.B(n_626),
.Y(n_836)
);

AND2x6_ASAP7_75t_SL g837 ( 
.A(n_740),
.B(n_592),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_735),
.B(n_410),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_717),
.B(n_626),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_743),
.B(n_414),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_740),
.A2(n_639),
.B1(n_599),
.B2(n_445),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_735),
.A2(n_460),
.B1(n_465),
.B2(n_437),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_747),
.B(n_417),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_726),
.B(n_751),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_702),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_731),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_698),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_752),
.A2(n_467),
.B1(n_421),
.B2(n_488),
.C(n_485),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_731),
.Y(n_849)
);

AND2x6_ASAP7_75t_SL g850 ( 
.A(n_740),
.B(n_599),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_699),
.B(n_737),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_679),
.B(n_639),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_752),
.A2(n_425),
.B1(n_427),
.B2(n_422),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_699),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_737),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_754),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_698),
.B(n_430),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_704),
.B(n_433),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_SL g859 ( 
.A(n_774),
.B(n_763),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_819),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_SL g861 ( 
.A(n_790),
.B(n_701),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_805),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_800),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_780),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_854),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_764),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_777),
.B(n_749),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_769),
.B(n_692),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_856),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_805),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_769),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_SL g874 ( 
.A(n_841),
.B(n_753),
.C(n_746),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_R g875 ( 
.A(n_804),
.B(n_732),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_793),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_784),
.B(n_706),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_796),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_785),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_773),
.A2(n_750),
.B1(n_704),
.B2(n_754),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_823),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_809),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_795),
.B(n_722),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_825),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_SL g885 ( 
.A(n_771),
.B(n_439),
.C(n_438),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_773),
.B(n_810),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_810),
.A2(n_761),
.B(n_692),
.C(n_760),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_834),
.B(n_704),
.Y(n_888)
);

OAI21xp33_ASAP7_75t_L g889 ( 
.A1(n_771),
.A2(n_760),
.B(n_722),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_855),
.B(n_707),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_770),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_851),
.B(n_728),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_820),
.B(n_729),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_SL g894 ( 
.A(n_817),
.B(n_768),
.C(n_848),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_769),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_766),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_818),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_851),
.B(n_728),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_833),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_852),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_779),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_798),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_802),
.Y(n_903)
);

BUFx5_ASAP7_75t_L g904 ( 
.A(n_824),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_806),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_832),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_835),
.B(n_792),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_844),
.A2(n_761),
.B(n_443),
.C(n_444),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_829),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_788),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_845),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_816),
.B(n_728),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_831),
.A2(n_446),
.B1(n_449),
.B2(n_442),
.Y(n_913)
);

INVx6_ASAP7_75t_L g914 ( 
.A(n_837),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_812),
.B(n_733),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_836),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_847),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_828),
.B(n_733),
.Y(n_918)
);

OR2x2_ASAP7_75t_SL g919 ( 
.A(n_849),
.B(n_850),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_781),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_846),
.B(n_733),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_799),
.A2(n_454),
.B(n_453),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_782),
.B(n_697),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_830),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_812),
.B(n_697),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_818),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_864),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_876),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_865),
.Y(n_929)
);

BUFx12f_ASAP7_75t_L g930 ( 
.A(n_860),
.Y(n_930)
);

AOI31xp67_ASAP7_75t_L g931 ( 
.A1(n_886),
.A2(n_797),
.A3(n_808),
.B(n_803),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_878),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_866),
.B(n_813),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_892),
.A2(n_778),
.B(n_776),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_866),
.B(n_898),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_890),
.A2(n_778),
.B(n_776),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_883),
.B(n_813),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_915),
.A2(n_789),
.B(n_781),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_867),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_894),
.A2(n_831),
.B1(n_838),
.B2(n_853),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_923),
.A2(n_842),
.B(n_767),
.C(n_838),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_924),
.A2(n_789),
.B(n_765),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_924),
.A2(n_797),
.B(n_803),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_867),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_925),
.A2(n_896),
.B(n_766),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_896),
.A2(n_791),
.B(n_857),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_920),
.A2(n_811),
.B(n_808),
.Y(n_947)
);

CKINVDCx11_ASAP7_75t_R g948 ( 
.A(n_870),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_866),
.B(n_772),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_866),
.B(n_807),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_868),
.Y(n_951)
);

NAND2x1_ASAP7_75t_L g952 ( 
.A(n_862),
.B(n_811),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_907),
.B(n_839),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_879),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_920),
.A2(n_857),
.B(n_786),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_887),
.A2(n_775),
.B(n_794),
.Y(n_956)
);

AO31x2_ASAP7_75t_L g957 ( 
.A1(n_913),
.A2(n_853),
.A3(n_815),
.B(n_821),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_896),
.A2(n_840),
.B(n_801),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_881),
.A2(n_822),
.B(n_814),
.Y(n_959)
);

OAI22x1_ASAP7_75t_L g960 ( 
.A1(n_877),
.A2(n_826),
.B1(n_787),
.B2(n_843),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_866),
.B(n_827),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_904),
.B(n_909),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_874),
.B(n_858),
.C(n_456),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_906),
.A2(n_56),
.B(n_55),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_900),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_911),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_904),
.B(n_455),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_904),
.B(n_457),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_906),
.A2(n_59),
.B(n_58),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_917),
.A2(n_62),
.B(n_60),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_885),
.A2(n_459),
.B1(n_462),
.B2(n_463),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_863),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_869),
.B(n_464),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_902),
.A2(n_65),
.B(n_64),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_902),
.A2(n_67),
.B(n_66),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_908),
.A2(n_470),
.B(n_466),
.Y(n_976)
);

INVx5_ASAP7_75t_L g977 ( 
.A(n_870),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_891),
.A2(n_70),
.B(n_68),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_901),
.A2(n_74),
.B(n_71),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_893),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_904),
.B(n_882),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_884),
.Y(n_982)
);

AO21x2_ASAP7_75t_L g983 ( 
.A1(n_956),
.A2(n_880),
.B(n_889),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_965),
.Y(n_984)
);

AO21x2_ASAP7_75t_L g985 ( 
.A1(n_956),
.A2(n_905),
.B(n_903),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_897),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_929),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_937),
.B(n_904),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_933),
.A2(n_918),
.B(n_912),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_953),
.A2(n_922),
.B1(n_916),
.B2(n_926),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_977),
.B(n_873),
.Y(n_991)
);

OAI211xp5_ASAP7_75t_L g992 ( 
.A1(n_940),
.A2(n_875),
.B(n_910),
.C(n_859),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_940),
.A2(n_918),
.B(n_912),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_939),
.Y(n_994)
);

OA21x2_ASAP7_75t_L g995 ( 
.A1(n_943),
.A2(n_921),
.B(n_472),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_942),
.A2(n_861),
.B(n_862),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_951),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_954),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_933),
.A2(n_872),
.B(n_921),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_935),
.A2(n_961),
.B(n_950),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_932),
.A2(n_895),
.B1(n_871),
.B2(n_888),
.C(n_475),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_927),
.Y(n_1002)
);

AOI221x1_ASAP7_75t_L g1003 ( 
.A1(n_941),
.A2(n_899),
.B1(n_863),
.B2(n_872),
.C(n_888),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_938),
.A2(n_899),
.B(n_863),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_966),
.Y(n_1005)
);

OA21x2_ASAP7_75t_L g1006 ( 
.A1(n_947),
.A2(n_473),
.B(n_471),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_932),
.B(n_919),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_944),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_973),
.B(n_899),
.Y(n_1009)
);

BUFx10_ASAP7_75t_L g1010 ( 
.A(n_972),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_SL g1011 ( 
.A1(n_962),
.A2(n_914),
.B(n_77),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_982),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_955),
.A2(n_724),
.B(n_79),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_962),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_934),
.A2(n_936),
.B(n_978),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_935),
.A2(n_724),
.B(n_481),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_957),
.B(n_479),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_981),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_963),
.A2(n_914),
.B1(n_483),
.B2(n_482),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_979),
.A2(n_724),
.B(n_81),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_964),
.A2(n_724),
.B(n_82),
.Y(n_1021)
);

AO21x2_ASAP7_75t_L g1022 ( 
.A1(n_967),
.A2(n_83),
.B(n_75),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_959),
.B(n_85),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_969),
.A2(n_90),
.B(n_89),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_928),
.B(n_8),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_974),
.A2(n_97),
.B(n_92),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_975),
.A2(n_99),
.B(n_98),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_972),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_972),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_931),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_963),
.B(n_959),
.C(n_971),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_970),
.A2(n_104),
.B(n_102),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_971),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1033)
);

OAI221xp5_ASAP7_75t_SL g1034 ( 
.A1(n_949),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_977),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_952),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_946),
.A2(n_106),
.B(n_105),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_987),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_1031),
.A2(n_960),
.B(n_967),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_994),
.Y(n_1040)
);

OAI211xp5_ASAP7_75t_L g1041 ( 
.A1(n_1033),
.A2(n_948),
.B(n_977),
.C(n_976),
.Y(n_1041)
);

CKINVDCx11_ASAP7_75t_R g1042 ( 
.A(n_1002),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1023),
.A2(n_930),
.B1(n_968),
.B2(n_958),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_990),
.B(n_957),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_1002),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1023),
.A2(n_945),
.B1(n_957),
.B2(n_14),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1034),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1014),
.B(n_16),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_1010),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_991),
.B(n_107),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_994),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_993),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_984),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_1029),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_997),
.Y(n_1055)
);

CKINVDCx6p67_ASAP7_75t_R g1056 ( 
.A(n_991),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_991),
.B(n_109),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_988),
.B(n_110),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1015),
.A2(n_120),
.B(n_117),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_998),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1005),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1025),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.C(n_22),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1009),
.B(n_22),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1007),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1007),
.B(n_23),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1000),
.A2(n_27),
.A3(n_29),
.B(n_30),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1028),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1008),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1012),
.B(n_30),
.Y(n_1069)
);

CKINVDCx8_ASAP7_75t_R g1070 ( 
.A(n_995),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1019),
.B(n_31),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_988),
.B(n_33),
.Y(n_1072)
);

OAI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1003),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_992),
.B(n_129),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1018),
.Y(n_1075)
);

INVx6_ASAP7_75t_L g1076 ( 
.A(n_1010),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_1035),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1001),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1078)
);

OAI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1017),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_986),
.B(n_39),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1029),
.B(n_40),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_999),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_983),
.B(n_43),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1029),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_983),
.B(n_44),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_983),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_985),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_989),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_1011),
.B(n_134),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1017),
.B(n_136),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_1010),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1003),
.A2(n_226),
.B(n_306),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_989),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_985),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1011),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1030),
.A2(n_1036),
.B1(n_995),
.B2(n_1006),
.Y(n_1097)
);

XOR2x2_ASAP7_75t_L g1098 ( 
.A(n_1065),
.B(n_45),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1075),
.B(n_1000),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1067),
.Y(n_1100)
);

OAI22x1_ASAP7_75t_L g1101 ( 
.A1(n_1086),
.A2(n_1006),
.B1(n_995),
.B2(n_1036),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1047),
.A2(n_1078),
.B1(n_1071),
.B2(n_1062),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1072),
.B(n_1022),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1061),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1053),
.B(n_1022),
.Y(n_1105)
);

OAI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1047),
.A2(n_1006),
.B1(n_1030),
.B2(n_1022),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_1073),
.A2(n_1016),
.B(n_1037),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1086),
.A2(n_1052),
.B1(n_1078),
.B2(n_1064),
.Y(n_1108)
);

OAI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_1043),
.A2(n_1037),
.B1(n_1032),
.B2(n_1027),
.C(n_1026),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_1038),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1064),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1111)
);

OAI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1079),
.A2(n_1027),
.B(n_1026),
.C(n_1024),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1040),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1042),
.Y(n_1114)
);

INVx4_ASAP7_75t_SL g1115 ( 
.A(n_1090),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1082),
.A2(n_1016),
.B1(n_50),
.B2(n_52),
.C(n_53),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1041),
.A2(n_1032),
.B1(n_1024),
.B2(n_1021),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1051),
.Y(n_1118)
);

OAI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1043),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1054),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1091),
.A2(n_1016),
.B1(n_996),
.B2(n_1021),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1039),
.B(n_49),
.C(n_54),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1077),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1093),
.A2(n_1039),
.B(n_1046),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1082),
.A2(n_54),
.B1(n_996),
.B2(n_1020),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1081),
.B(n_137),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1044),
.A2(n_1020),
.B1(n_1013),
.B2(n_1015),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1068),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1048),
.A2(n_1004),
.B1(n_1013),
.B2(n_142),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_L g1130 ( 
.A(n_1056),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1080),
.B(n_138),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1048),
.B(n_1004),
.Y(n_1132)
);

OAI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1074),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.C(n_146),
.Y(n_1133)
);

AOI222xp33_ASAP7_75t_L g1134 ( 
.A1(n_1063),
.A2(n_147),
.B1(n_149),
.B2(n_151),
.C1(n_156),
.C2(n_160),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1090),
.B(n_161),
.C(n_163),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1090),
.A2(n_1057),
.B1(n_1050),
.B2(n_1096),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1050),
.A2(n_165),
.B1(n_167),
.B2(n_169),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1057),
.A2(n_1058),
.B1(n_1083),
.B2(n_1085),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1058),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1045),
.A2(n_176),
.B1(n_178),
.B2(n_185),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1069),
.B(n_191),
.C(n_192),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1055),
.A2(n_193),
.B1(n_195),
.B2(n_198),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1045),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1060),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1084),
.B(n_212),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1059),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1049),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1066),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1097),
.A2(n_216),
.B1(n_219),
.B2(n_222),
.C(n_223),
.Y(n_1149)
);

OAI221xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1089),
.A2(n_224),
.B1(n_227),
.B2(n_230),
.C(n_232),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1092),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1049),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1103),
.B(n_1095),
.Y(n_1153)
);

OAI33xp33_ASAP7_75t_L g1154 ( 
.A1(n_1111),
.A2(n_1097),
.A3(n_1066),
.B1(n_1088),
.B2(n_1087),
.B3(n_1070),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1100),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1110),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1115),
.B(n_1094),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1110),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1108),
.A2(n_1119),
.B1(n_1136),
.B2(n_1122),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1128),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1115),
.B(n_1094),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1104),
.Y(n_1162)
);

INVx4_ASAP7_75t_SL g1163 ( 
.A(n_1125),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1099),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1113),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1118),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1148),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_1107),
.A2(n_1054),
.B(n_1076),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1132),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1147),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1105),
.B(n_240),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1138),
.B(n_1076),
.Y(n_1172)
);

INVxp33_ASAP7_75t_L g1173 ( 
.A(n_1123),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1115),
.B(n_241),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1101),
.B(n_242),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1152),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1127),
.B(n_244),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1120),
.B(n_245),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1129),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1106),
.B(n_246),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1124),
.B(n_247),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1129),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1109),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1120),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1135),
.B(n_248),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1112),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1111),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1121),
.B(n_249),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1107),
.B(n_251),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1145),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1131),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1126),
.B(n_252),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1117),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1141),
.B(n_255),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1108),
.B(n_1116),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1130),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1159),
.A2(n_1133),
.B1(n_1149),
.B2(n_1114),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1156),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1162),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1155),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1195),
.A2(n_1102),
.B1(n_1150),
.B2(n_1144),
.C(n_1151),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1174),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1167),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1158),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1195),
.A2(n_1134),
.B(n_1098),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1160),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1186),
.A2(n_1139),
.B(n_1142),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1153),
.B(n_1114),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1168),
.A2(n_1134),
.B(n_1146),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_SL g1210 ( 
.A1(n_1185),
.A2(n_1174),
.B(n_1194),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1168),
.A2(n_1186),
.B(n_1183),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1196),
.B(n_1114),
.Y(n_1212)
);

NAND4xp25_ASAP7_75t_SL g1213 ( 
.A(n_1193),
.B(n_1137),
.C(n_1140),
.D(n_1143),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1162),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1153),
.B(n_257),
.Y(n_1215)
);

AOI32xp33_ASAP7_75t_L g1216 ( 
.A1(n_1181),
.A2(n_1130),
.A3(n_261),
.B1(n_267),
.B2(n_269),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1167),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1163),
.A2(n_259),
.B1(n_272),
.B2(n_273),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1217),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1217),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1208),
.B(n_1155),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1212),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1198),
.B(n_1169),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1199),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1200),
.B(n_1169),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1203),
.B(n_1157),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1203),
.B(n_1157),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1199),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1214),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1208),
.B(n_1170),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1211),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1214),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1206),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1204),
.B(n_1164),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1211),
.B(n_1170),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1222),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1219),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1233),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1230),
.B(n_1173),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1225),
.B(n_1211),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1219),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1221),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1230),
.B(n_1202),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1225),
.B(n_1183),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1221),
.B(n_1215),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1223),
.B(n_1215),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1226),
.B(n_1184),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1243),
.B(n_1247),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1238),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1236),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1247),
.B(n_1242),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1239),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1244),
.B(n_1234),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1245),
.B(n_1235),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1246),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1240),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1237),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1241),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1237),
.B(n_1235),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1236),
.B(n_1205),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1238),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1260),
.A2(n_1216),
.B(n_1201),
.C(n_1179),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1250),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_1260),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1249),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1261),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1248),
.B(n_1226),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1248),
.B(n_1226),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1257),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1255),
.A2(n_1197),
.B1(n_1182),
.B2(n_1213),
.C(n_1210),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1267),
.B(n_1251),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1269),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1265),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1266),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1263),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1264),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1276),
.B(n_1264),
.Y(n_1277)
);

NOR2x1_ASAP7_75t_SL g1278 ( 
.A(n_1275),
.B(n_1268),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1271),
.B(n_1252),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1272),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1271),
.B(n_1270),
.Y(n_1281)
);

NOR4xp25_ASAP7_75t_SL g1282 ( 
.A(n_1273),
.B(n_1270),
.C(n_1262),
.D(n_1190),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_L g1283 ( 
.A(n_1277),
.B(n_1274),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1279),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_L g1285 ( 
.A(n_1282),
.B(n_1181),
.C(n_1218),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1279),
.B(n_1251),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1278),
.B(n_1254),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1281),
.A2(n_1258),
.B1(n_1256),
.B2(n_1193),
.Y(n_1288)
);

NAND4xp25_ASAP7_75t_L g1289 ( 
.A(n_1280),
.B(n_1210),
.C(n_1196),
.D(n_1172),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1279),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1290),
.A2(n_1283),
.B(n_1288),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1284),
.Y(n_1292)
);

OAI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1285),
.A2(n_1196),
.B1(n_1253),
.B2(n_1202),
.C(n_1171),
.Y(n_1293)
);

AOI211x1_ASAP7_75t_SL g1294 ( 
.A1(n_1286),
.A2(n_1220),
.B(n_1191),
.C(n_1163),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1289),
.A2(n_1287),
.B1(n_1259),
.B2(n_1254),
.C(n_1175),
.Y(n_1295)
);

AOI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1288),
.A2(n_1209),
.B1(n_1231),
.B2(n_1259),
.C(n_1154),
.Y(n_1296)
);

OAI221xp5_ASAP7_75t_L g1297 ( 
.A1(n_1285),
.A2(n_1171),
.B1(n_1180),
.B2(n_1189),
.C(n_1207),
.Y(n_1297)
);

AOI211xp5_ASAP7_75t_L g1298 ( 
.A1(n_1291),
.A2(n_1292),
.B(n_1297),
.C(n_1293),
.Y(n_1298)
);

XOR2xp5_ASAP7_75t_L g1299 ( 
.A(n_1294),
.B(n_1192),
.Y(n_1299)
);

XNOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1296),
.B(n_1185),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1295),
.B(n_1227),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1292),
.Y(n_1302)
);

NAND4xp25_ASAP7_75t_SL g1303 ( 
.A(n_1295),
.B(n_1163),
.C(n_1180),
.D(n_1175),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1292),
.B(n_1228),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1292),
.B(n_1227),
.Y(n_1305)
);

AOI222xp33_ASAP7_75t_L g1306 ( 
.A1(n_1300),
.A2(n_1163),
.B1(n_1185),
.B2(n_1194),
.C1(n_1189),
.C2(n_1188),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1302),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1305),
.B(n_1192),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1304),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_L g1310 ( 
.A(n_1303),
.B(n_1174),
.Y(n_1310)
);

NAND4xp75_ASAP7_75t_L g1311 ( 
.A(n_1301),
.B(n_1298),
.C(n_1299),
.D(n_1188),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1298),
.A2(n_1177),
.B1(n_1187),
.B2(n_1232),
.C(n_1229),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1302),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_L g1314 ( 
.A(n_1302),
.B(n_1192),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_SL g1315 ( 
.A(n_1307),
.B(n_1177),
.C(n_1190),
.Y(n_1315)
);

XOR2xp5_ASAP7_75t_L g1316 ( 
.A(n_1311),
.B(n_1194),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1313),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1309),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1314),
.B(n_1227),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1308),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1310),
.A2(n_1209),
.B1(n_1178),
.B2(n_1207),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1312),
.A2(n_1209),
.B1(n_1178),
.B2(n_1207),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1306),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1307),
.B(n_1224),
.Y(n_1324)
);

NAND4xp25_ASAP7_75t_L g1325 ( 
.A(n_1307),
.B(n_1178),
.C(n_1191),
.D(n_1157),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1317),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1318),
.B(n_1232),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1323),
.Y(n_1328)
);

NOR3xp33_ASAP7_75t_L g1329 ( 
.A(n_1320),
.B(n_1176),
.C(n_1161),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1316),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1324),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1319),
.B(n_1224),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1315),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1326),
.B(n_1325),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1333),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1330),
.Y(n_1336)
);

XNOR2xp5_ASAP7_75t_L g1337 ( 
.A(n_1328),
.B(n_1321),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1335),
.B(n_1331),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1336),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1338),
.B(n_1337),
.C(n_1339),
.Y(n_1340)
);

AOI21xp33_ASAP7_75t_L g1341 ( 
.A1(n_1338),
.A2(n_1334),
.B(n_1327),
.Y(n_1341)
);

AOI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1341),
.A2(n_1332),
.B(n_1322),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1340),
.Y(n_1343)
);

AOI222xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1340),
.A2(n_1329),
.B1(n_1224),
.B2(n_1229),
.C1(n_1220),
.C2(n_282),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1343),
.B(n_1168),
.Y(n_1345)
);

AOI222xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1344),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.C1(n_281),
.C2(n_283),
.Y(n_1346)
);

AOI322xp5_ASAP7_75t_L g1347 ( 
.A1(n_1346),
.A2(n_1342),
.A3(n_1345),
.B1(n_1161),
.B2(n_1166),
.C1(n_1165),
.C2(n_298),
.Y(n_1347)
);

OAI221xp5_ASAP7_75t_R g1348 ( 
.A1(n_1347),
.A2(n_285),
.B1(n_286),
.B2(n_293),
.C(n_294),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1348),
.A2(n_1161),
.B1(n_1165),
.B2(n_1166),
.Y(n_1349)
);


endmodule