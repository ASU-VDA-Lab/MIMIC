module fake_jpeg_11680_n_441 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_3),
.B(n_9),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_57),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_72),
.Y(n_113)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_92),
.Y(n_134)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_86),
.Y(n_124)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_10),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_10),
.B(n_1),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_93),
.A2(n_39),
.B(n_30),
.C(n_4),
.Y(n_153)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_95),
.B(n_109),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_102),
.Y(n_129)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_95),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_112),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_117),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_24),
.B1(n_28),
.B2(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_118),
.A2(n_128),
.B1(n_130),
.B2(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_29),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_6),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_28),
.B1(n_35),
.B2(n_52),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_35),
.B1(n_34),
.B2(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_21),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_131),
.B(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_43),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_170),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_60),
.A2(n_49),
.B1(n_38),
.B2(n_30),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_137),
.A2(n_165),
.B1(n_173),
.B2(n_175),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_38),
.B1(n_49),
.B2(n_45),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_147),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_65),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_108),
.B(n_7),
.C(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_162),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_90),
.A2(n_39),
.B1(n_43),
.B2(n_27),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_101),
.A2(n_50),
.B1(n_33),
.B2(n_31),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_50),
.B1(n_33),
.B2(n_31),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_68),
.B(n_26),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_25),
.B1(n_27),
.B2(n_4),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_87),
.B(n_25),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_9),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_75),
.A2(n_25),
.B1(n_2),
.B2(n_5),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_110),
.B1(n_91),
.B2(n_100),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_99),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_99),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_179),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_186),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_181),
.A2(n_198),
.B(n_202),
.C(n_212),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_57),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_182),
.B(n_206),
.C(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_129),
.Y(n_186)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_194),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_10),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_116),
.B(n_76),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_203),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_134),
.A2(n_79),
.B(n_64),
.C(n_69),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_200),
.A2(n_163),
.B1(n_178),
.B2(n_217),
.Y(n_270)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_70),
.B1(n_83),
.B2(n_170),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_132),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_133),
.B(n_140),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_120),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_113),
.B(n_124),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_208),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_123),
.B(n_127),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_214),
.Y(n_269)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

OR2x4_ASAP7_75t_L g212 ( 
.A(n_122),
.B(n_125),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_143),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_144),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_225),
.Y(n_272)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

AOI22x1_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_151),
.B1(n_139),
.B2(n_121),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_224),
.A2(n_177),
.B1(n_178),
.B2(n_163),
.Y(n_268)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_122),
.B(n_142),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_125),
.B(n_142),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_231),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_167),
.B(n_146),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_121),
.A2(n_159),
.B1(n_114),
.B2(n_146),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_114),
.B1(n_150),
.B2(n_157),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_164),
.B(n_141),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_234),
.Y(n_247)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_187),
.A2(n_150),
.B1(n_157),
.B2(n_177),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_258),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_250),
.A2(n_278),
.B1(n_267),
.B2(n_244),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_197),
.B1(n_194),
.B2(n_187),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_268),
.B1(n_273),
.B2(n_182),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_221),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_270),
.A2(n_246),
.B1(n_257),
.B2(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_189),
.B(n_182),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_232),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_219),
.A2(n_224),
.B1(n_215),
.B2(n_192),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_184),
.A2(n_195),
.B1(n_217),
.B2(n_202),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_281),
.A2(n_286),
.B1(n_293),
.B2(n_310),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_282),
.B(n_289),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_287),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_224),
.B1(n_202),
.B2(n_198),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_249),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_181),
.B1(n_202),
.B2(n_206),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_270),
.A2(n_208),
.B1(n_190),
.B2(n_212),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_292),
.A2(n_294),
.B1(n_302),
.B2(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_206),
.B1(n_210),
.B2(n_204),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_222),
.B(n_216),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_295),
.A2(n_261),
.B(n_262),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_220),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_307),
.C(n_242),
.Y(n_332)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_241),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_299),
.B(n_303),
.Y(n_337)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_243),
.A2(n_235),
.B1(n_211),
.B2(n_201),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_185),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_238),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_213),
.C(n_179),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_238),
.A2(n_179),
.B1(n_252),
.B2(n_239),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_265),
.B1(n_245),
.B2(n_278),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_255),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_247),
.A2(n_259),
.B1(n_251),
.B2(n_240),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_240),
.B1(n_251),
.B2(n_248),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_314),
.B1(n_262),
.B2(n_267),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_269),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_248),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_256),
.C(n_261),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_333),
.B(n_297),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_291),
.B(n_288),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_324),
.B(n_331),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_339),
.Y(n_345)
);

AO22x1_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_245),
.B1(n_265),
.B2(n_256),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_279),
.B(n_276),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_334),
.C(n_295),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_279),
.B(n_276),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_275),
.C(n_254),
.Y(n_334)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_281),
.A2(n_280),
.B1(n_254),
.B2(n_242),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_294),
.A2(n_292),
.B1(n_285),
.B2(n_299),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_340),
.A2(n_307),
.B1(n_313),
.B2(n_309),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_324),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_343),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_325),
.B(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_325),
.B(n_296),
.Y(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_355),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_340),
.A2(n_286),
.B1(n_285),
.B2(n_293),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_353),
.B1(n_357),
.B2(n_358),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_323),
.A2(n_282),
.B1(n_310),
.B2(n_311),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_317),
.C(n_335),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_330),
.C(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_326),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_329),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_360),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_323),
.A2(n_307),
.B1(n_312),
.B2(n_289),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_284),
.B1(n_298),
.B2(n_290),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_362),
.B1(n_321),
.B2(n_320),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_338),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_335),
.A2(n_283),
.B1(n_302),
.B2(n_301),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_338),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_363),
.B(n_350),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_351),
.A2(n_327),
.B1(n_320),
.B2(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_376),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_381),
.C(n_341),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_316),
.B1(n_319),
.B2(n_331),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_319),
.C(n_316),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_358),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g376 ( 
.A1(n_355),
.A2(n_322),
.A3(n_324),
.B1(n_339),
.B2(n_306),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_345),
.B1(n_360),
.B2(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_344),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_364),
.A2(n_366),
.B1(n_345),
.B2(n_379),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_368),
.A2(n_351),
.B1(n_347),
.B2(n_354),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_385),
.A2(n_392),
.B1(n_378),
.B2(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_341),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_396),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_373),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_391),
.C(n_370),
.Y(n_398)
);

AO21x1_ASAP7_75t_L g389 ( 
.A1(n_368),
.A2(n_352),
.B(n_353),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_376),
.B(n_372),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_354),
.C(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_393),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_349),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_380),
.Y(n_403)
);

AO22x1_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_333),
.B1(n_342),
.B2(n_361),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_397),
.A2(n_402),
.B1(n_405),
.B2(n_392),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_406),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_385),
.B(n_348),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_407),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_373),
.B1(n_371),
.B2(n_380),
.Y(n_402)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_362),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_388),
.B(n_322),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_386),
.C(n_383),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_411),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_383),
.C(n_389),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_396),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_401),
.Y(n_422)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_408),
.A2(n_384),
.B1(n_390),
.B2(n_396),
.Y(n_417)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_417),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_417),
.A2(n_408),
.B(n_384),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_422),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_399),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_420),
.A2(n_394),
.B(n_397),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_402),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_424),
.B(n_414),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_425),
.B(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_428),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_410),
.C(n_416),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_421),
.A2(n_390),
.B1(n_411),
.B2(n_372),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_412),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_430),
.B(n_346),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_420),
.C(n_419),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_434),
.Y(n_436)
);

AO221x1_ASAP7_75t_L g435 ( 
.A1(n_432),
.A2(n_427),
.B1(n_346),
.B2(n_336),
.C(n_304),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_433),
.B(n_427),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_436),
.B(n_263),
.Y(n_438)
);

BUFx24_ASAP7_75t_SL g439 ( 
.A(n_438),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_263),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_440),
.B(n_275),
.Y(n_441)
);


endmodule