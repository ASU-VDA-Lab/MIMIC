module fake_jpeg_13250_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_12),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_51),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g141 ( 
.A(n_50),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_52),
.Y(n_115)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_54),
.B(n_79),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_61),
.B(n_66),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_20),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_69),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_98),
.B1(n_47),
.B2(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_71),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_81),
.Y(n_121)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_10),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_84),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_33),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_91),
.Y(n_134)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_97),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_37),
.B(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_26),
.B1(n_45),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_104),
.B1(n_107),
.B2(n_111),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_43),
.B1(n_41),
.B2(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_45),
.B1(n_26),
.B2(n_36),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_105),
.A2(n_147),
.B1(n_68),
.B2(n_64),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_45),
.B1(n_36),
.B2(n_35),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_118),
.B(n_143),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_65),
.B1(n_96),
.B2(n_89),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_35),
.B1(n_25),
.B2(n_39),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_38),
.B1(n_1),
.B2(n_0),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_114),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_1),
.B1(n_12),
.B2(n_13),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_1),
.B1(n_14),
.B2(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_14),
.B1(n_75),
.B2(n_60),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_53),
.A2(n_74),
.B1(n_52),
.B2(n_62),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_88),
.A2(n_59),
.B1(n_81),
.B2(n_92),
.Y(n_147)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_179),
.B1(n_181),
.B2(n_146),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_69),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_154),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_155),
.Y(n_187)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_81),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

OA22x2_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_50),
.B1(n_58),
.B2(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_58),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_115),
.C(n_127),
.Y(n_205)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_164),
.Y(n_186)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_119),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_173),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_103),
.B(n_113),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_176),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_109),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_106),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_108),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_207),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_118),
.B(n_143),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_197),
.B(n_158),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_105),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_149),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_127),
.B(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_171),
.B1(n_152),
.B2(n_178),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_210),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_169),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_160),
.B(n_179),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_224),
.B(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_189),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_168),
.B1(n_159),
.B2(n_133),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_221),
.B1(n_229),
.B2(n_195),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_187),
.A2(n_168),
.B1(n_133),
.B2(n_136),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_160),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_199),
.C(n_205),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_166),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_136),
.B1(n_110),
.B2(n_158),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_247),
.C(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_237),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_232),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_218),
.B(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_183),
.B1(n_199),
.B2(n_202),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_243),
.B1(n_245),
.B2(n_217),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_202),
.B1(n_190),
.B2(n_184),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_184),
.B1(n_203),
.B2(n_167),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_215),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_188),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_219),
.B(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_251),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_212),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_218),
.B(n_211),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_254),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_209),
.B1(n_214),
.B2(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_228),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_235),
.C(n_247),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_270),
.C(n_274),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_244),
.B(n_246),
.C(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_267),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_254),
.B(n_261),
.C(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_259),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_241),
.C(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_243),
.C(n_222),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_260),
.A3(n_257),
.B1(n_249),
.B2(n_252),
.C1(n_255),
.C2(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_266),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_285),
.B1(n_273),
.B2(n_271),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_256),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_245),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_284),
.C(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_295),
.B1(n_129),
.B2(n_116),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_265),
.B1(n_203),
.B2(n_185),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_194),
.B1(n_185),
.B2(n_201),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_201),
.B1(n_185),
.B2(n_170),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_297),
.B1(n_301),
.B2(n_302),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_281),
.C(n_286),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_300),
.C(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_286),
.C(n_181),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_194),
.B1(n_153),
.B2(n_156),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_194),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_308),
.C(n_163),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_290),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_308),
.A3(n_305),
.B1(n_194),
.B2(n_148),
.C1(n_137),
.C2(n_116),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_117),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_125),
.A3(n_101),
.B1(n_165),
.B2(n_161),
.C1(n_139),
.C2(n_144),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_101),
.A3(n_125),
.B1(n_139),
.B2(n_144),
.C1(n_122),
.C2(n_117),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.C(n_122),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_313),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_135),
.B(n_312),
.Y(n_320)
);


endmodule