module fake_jpeg_20986_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_20),
.B(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_53),
.C(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_80),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_41),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_41),
.B1(n_49),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_47),
.B1(n_62),
.B2(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_58),
.B1(n_52),
.B2(n_57),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_42),
.C(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_0),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_89),
.B1(n_96),
.B2(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_92),
.Y(n_109)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_93),
.B1(n_5),
.B2(n_6),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_40),
.B1(n_46),
.B2(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_60),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_59),
.B1(n_54),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_99),
.B1(n_110),
.B2(n_7),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_104),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_44),
.B(n_2),
.C(n_4),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_0),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_2),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_21),
.B(n_37),
.C(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_5),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_23),
.C(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_117),
.Y(n_122)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_104),
.C(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_107),
.B(n_110),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_114),
.B(n_10),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.C(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_116),
.B1(n_118),
.B2(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_122),
.C(n_113),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_9),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_28),
.B(n_33),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_25),
.Y(n_137)
);


endmodule