module real_aes_5727_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g130 ( .A(n_0), .B(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_1), .Y(n_177) );
OA22x2_ASAP7_75t_L g118 ( .A1(n_2), .A2(n_119), .B1(n_120), .B2(n_121), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_2), .Y(n_119) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_3), .A2(n_172), .B(n_204), .C(n_205), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g143 ( .A1(n_4), .A2(n_84), .B1(n_138), .B2(n_144), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_5), .A2(n_31), .B1(n_603), .B2(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
BUFx2_ASAP7_75t_L g943 ( .A(n_6), .Y(n_943) );
INVx1_ASAP7_75t_L g950 ( .A(n_6), .Y(n_950) );
OAI22x1_ASAP7_75t_R g525 ( .A1(n_7), .A2(n_83), .B1(n_526), .B2(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_7), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_8), .A2(n_91), .B1(n_645), .B2(n_646), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_9), .A2(n_59), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_9), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_10), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_11), .A2(n_70), .B1(n_144), .B2(n_159), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_12), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_13), .A2(n_32), .B1(n_590), .B2(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g575 ( .A(n_14), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_15), .A2(n_64), .B1(n_138), .B2(n_178), .Y(n_240) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_16), .A2(n_69), .B(n_134), .Y(n_133) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_16), .A2(n_69), .B(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_17), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g573 ( .A(n_18), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_19), .B(n_181), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_20), .Y(n_270) );
BUFx3_ASAP7_75t_L g540 ( .A(n_21), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_22), .A2(n_145), .B(n_210), .C(n_211), .Y(n_209) );
OAI22xp33_ASAP7_75t_SL g137 ( .A1(n_23), .A2(n_49), .B1(n_138), .B2(n_139), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_24), .A2(n_30), .B1(n_139), .B2(n_155), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g597 ( .A1(n_25), .A2(n_598), .B(n_601), .C(n_604), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_26), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_27), .B(n_535), .Y(n_534) );
O2A1O1Ixp5_ASAP7_75t_L g221 ( .A1(n_28), .A2(n_172), .B(n_222), .C(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g117 ( .A(n_29), .Y(n_117) );
AND2x2_ASAP7_75t_L g962 ( .A(n_33), .B(n_963), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_34), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_35), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_36), .A2(n_40), .B1(n_648), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_37), .A2(n_68), .B1(n_610), .B2(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_38), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g681 ( .A(n_39), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_41), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_42), .B(n_163), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_43), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_44), .A2(n_145), .B(n_571), .C(n_572), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_45), .A2(n_548), .B1(n_549), .B2(n_552), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_45), .Y(n_552) );
INVx1_ASAP7_75t_L g718 ( .A(n_46), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_47), .Y(n_946) );
INVx2_ASAP7_75t_L g612 ( .A(n_48), .Y(n_612) );
INVx1_ASAP7_75t_L g134 ( .A(n_50), .Y(n_134) );
AND2x4_ASAP7_75t_L g147 ( .A(n_51), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g215 ( .A(n_51), .B(n_148), .Y(n_215) );
INVx2_ASAP7_75t_L g674 ( .A(n_52), .Y(n_674) );
INVxp67_ASAP7_75t_SL g200 ( .A(n_53), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_53), .B(n_166), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_53), .A2(n_67), .B1(n_166), .B2(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_55), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_56), .Y(n_231) );
INVx2_ASAP7_75t_L g198 ( .A(n_57), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_58), .A2(n_172), .B(n_272), .C(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g550 ( .A(n_59), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_60), .Y(n_174) );
INVx1_ASAP7_75t_SL g602 ( .A(n_61), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_62), .B(n_181), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_63), .A2(n_79), .B1(n_158), .B2(n_160), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_65), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_66), .Y(n_179) );
NAND2xp33_ASAP7_75t_R g244 ( .A(n_67), .B(n_190), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_71), .A2(n_145), .B(n_603), .C(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g964 ( .A(n_72), .B(n_965), .Y(n_964) );
OR2x6_ASAP7_75t_L g114 ( .A(n_73), .B(n_115), .Y(n_114) );
AND3x1_ASAP7_75t_L g961 ( .A(n_73), .B(n_943), .C(n_962), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_74), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g704 ( .A(n_75), .Y(n_704) );
INVx1_ASAP7_75t_L g714 ( .A(n_76), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_77), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_78), .B(n_590), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g567 ( .A(n_80), .B(n_222), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_81), .A2(n_172), .B(n_671), .C(n_673), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_81), .A2(n_172), .B(n_671), .C(n_673), .Y(n_697) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_82), .B(n_117), .Y(n_960) );
INVx1_ASAP7_75t_L g526 ( .A(n_83), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_85), .A2(n_96), .B1(n_634), .B2(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g963 ( .A(n_86), .Y(n_963) );
BUFx5_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g156 ( .A(n_87), .Y(n_156) );
INVx2_ASAP7_75t_L g217 ( .A(n_88), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_89), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g276 ( .A(n_90), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_92), .Y(n_212) );
INVx2_ASAP7_75t_SL g148 ( .A(n_93), .Y(n_148) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_94), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_94), .Y(n_545) );
INVx1_ASAP7_75t_L g229 ( .A(n_95), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_97), .B(n_190), .Y(n_715) );
INVx1_ASAP7_75t_SL g665 ( .A(n_98), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_99), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g234 ( .A(n_100), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_101), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_SL g531 ( .A(n_101), .Y(n_531) );
AND2x2_ASAP7_75t_L g638 ( .A(n_101), .B(n_189), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g268 ( .A1(n_102), .A2(n_138), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g611 ( .A(n_103), .Y(n_611) );
AOI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_955), .B(n_964), .Y(n_104) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_536), .B(n_541), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_118), .B(n_529), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp67_ASAP7_75t_R g530 ( .A(n_109), .B(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_SL g535 ( .A(n_110), .Y(n_535) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx8_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_114), .A2(n_543), .B(n_945), .Y(n_542) );
OR2x6_ASAP7_75t_L g949 ( .A(n_114), .B(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AOI21x1_ASAP7_75t_L g529 ( .A1(n_118), .A2(n_530), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI22x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_525), .B2(n_528), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g944 ( .A(n_123), .Y(n_944) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_416), .Y(n_123) );
NAND4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_313), .C(n_353), .D(n_387), .Y(n_124) );
AOI211xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_183), .B(n_245), .C(n_304), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_149), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_127), .A2(n_290), .B1(n_400), .B2(n_402), .Y(n_399) );
BUFx3_ASAP7_75t_L g413 ( .A(n_127), .Y(n_413) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g262 ( .A(n_128), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_128), .B(n_317), .Y(n_343) );
AND2x4_ASAP7_75t_L g385 ( .A(n_128), .B(n_307), .Y(n_385) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g290 ( .A(n_129), .Y(n_290) );
AND2x2_ASAP7_75t_L g310 ( .A(n_129), .B(n_307), .Y(n_310) );
INVx2_ASAP7_75t_L g328 ( .A(n_129), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_129), .B(n_263), .Y(n_338) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_129), .Y(n_370) );
NAND2xp33_ASAP7_75t_R g466 ( .A(n_129), .B(n_263), .Y(n_466) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
INVx2_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_131), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_132), .B(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_132), .B(n_217), .Y(n_216) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx2_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_142), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_137), .B(n_141), .Y(n_136) );
AOI22xp33_ASAP7_75t_SL g173 ( .A1(n_138), .A2(n_139), .B1(n_174), .B2(n_175), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_138), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_138), .A2(n_139), .B1(n_193), .B2(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_138), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_138), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_138), .B(n_270), .Y(n_269) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_138), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g585 ( .A(n_138), .Y(n_585) );
INVx2_ASAP7_75t_L g590 ( .A(n_138), .Y(n_590) );
INVx2_ASAP7_75t_L g636 ( .A(n_138), .Y(n_636) );
INVx2_ASAP7_75t_L g645 ( .A(n_138), .Y(n_645) );
INVx1_ASAP7_75t_L g672 ( .A(n_138), .Y(n_672) );
INVx2_ASAP7_75t_SL g160 ( .A(n_139), .Y(n_160) );
INVx2_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
INVx1_ASAP7_75t_L g588 ( .A(n_139), .Y(n_588) );
INVx2_ASAP7_75t_L g600 ( .A(n_139), .Y(n_600) );
INVx1_ASAP7_75t_L g707 ( .A(n_139), .Y(n_707) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g144 ( .A(n_140), .Y(n_144) );
INVx2_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
INVx3_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
INVx3_ASAP7_75t_L g145 ( .A(n_141), .Y(n_145) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx1_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
INVx4_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_141), .B(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_L g607 ( .A(n_141), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_146), .Y(n_142) );
INVx2_ASAP7_75t_L g610 ( .A(n_144), .Y(n_610) );
INVx1_ASAP7_75t_L g709 ( .A(n_144), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g171 ( .A1(n_145), .A2(n_147), .B1(n_172), .B2(n_173), .C(n_176), .Y(n_171) );
INVx3_ASAP7_75t_L g631 ( .A(n_145), .Y(n_631) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g243 ( .A(n_147), .Y(n_243) );
INVx3_ASAP7_75t_L g592 ( .A(n_147), .Y(n_592) );
AND2x2_ASAP7_75t_L g637 ( .A(n_147), .B(n_162), .Y(n_637) );
INVx2_ASAP7_75t_L g367 ( .A(n_149), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_149), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
AND2x2_ASAP7_75t_L g521 ( .A(n_149), .B(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_167), .Y(n_149) );
OR2x2_ASAP7_75t_L g337 ( .A(n_150), .B(n_307), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_162), .B(n_164), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_152), .A2(n_165), .B(n_280), .Y(n_279) );
OA22x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_157), .B2(n_161), .Y(n_152) );
INVx4_ASAP7_75t_L g604 ( .A(n_153), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_155), .A2(n_178), .B1(n_197), .B2(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_155), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_155), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g635 ( .A(n_155), .Y(n_635) );
INVx2_ASAP7_75t_L g648 ( .A(n_155), .Y(n_648) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g159 ( .A(n_156), .Y(n_159) );
INVx1_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
INVx3_ASAP7_75t_L g603 ( .A(n_158), .Y(n_603) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_162), .B(n_187), .Y(n_667) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_163), .B(n_243), .Y(n_613) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g641 ( .A(n_166), .Y(n_641) );
AND2x4_ASAP7_75t_L g327 ( .A(n_167), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_168), .B(n_263), .Y(n_291) );
INVx2_ASAP7_75t_L g372 ( .A(n_168), .Y(n_372) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_180), .Y(n_168) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_169), .A2(n_171), .B(n_180), .Y(n_307) );
NOR2x1_ASAP7_75t_SL g562 ( .A(n_169), .B(n_214), .Y(n_562) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g199 ( .A(n_170), .B(n_200), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B1(n_195), .B2(n_196), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_172), .A2(n_195), .B1(n_240), .B2(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
INVx1_ASAP7_75t_L g568 ( .A(n_172), .Y(n_568) );
INVx2_ASAP7_75t_SL g649 ( .A(n_172), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_172), .B(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_172), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_178), .Y(n_571) );
INVx2_ASAP7_75t_L g630 ( .A(n_178), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_181), .B(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx3_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_182), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_182), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_218), .Y(n_183) );
AND2x2_ASAP7_75t_L g312 ( .A(n_184), .B(n_257), .Y(n_312) );
INVx2_ASAP7_75t_SL g320 ( .A(n_184), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_184), .A2(n_322), .B1(n_329), .B2(n_334), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_184), .B(n_218), .Y(n_340) );
AND2x2_ASAP7_75t_L g396 ( .A(n_184), .B(n_391), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_184), .B(n_283), .Y(n_516) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_201), .Y(n_184) );
INVx1_ASAP7_75t_L g404 ( .A(n_185), .Y(n_404) );
AND2x2_ASAP7_75t_L g481 ( .A(n_185), .B(n_237), .Y(n_481) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_191), .B(n_199), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_187), .B(n_643), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_188), .B(n_215), .Y(n_280) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
INVx1_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
INVx2_ASAP7_75t_L g302 ( .A(n_190), .Y(n_302) );
INVx1_ASAP7_75t_L g621 ( .A(n_190), .Y(n_621) );
INVx1_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_227), .B1(n_228), .B2(n_230), .Y(n_226) );
INVx2_ASAP7_75t_L g253 ( .A(n_195), .Y(n_253) );
O2A1O1Ixp5_ASAP7_75t_SL g703 ( .A1(n_195), .A2(n_704), .B(n_705), .C(n_708), .Y(n_703) );
INVx1_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
AND2x2_ASAP7_75t_L g248 ( .A(n_201), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g286 ( .A(n_201), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_201), .B(n_219), .Y(n_303) );
INVx2_ASAP7_75t_L g333 ( .A(n_201), .Y(n_333) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_201), .Y(n_352) );
INVx1_ASAP7_75t_L g386 ( .A(n_201), .Y(n_386) );
OR2x2_ASAP7_75t_L g432 ( .A(n_201), .B(n_249), .Y(n_432) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_201), .Y(n_449) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_208), .A3(n_213), .B(n_216), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_206), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_210), .A2(n_609), .B1(n_611), .B2(n_612), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_214), .B(n_221), .C(n_226), .Y(n_220) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_214), .A2(n_253), .B1(n_254), .B2(n_255), .C(n_256), .Y(n_252) );
NOR4xp25_ASAP7_75t_L g696 ( .A(n_214), .B(n_615), .C(n_676), .D(n_697), .Y(n_696) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g265 ( .A(n_215), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g362 ( .A(n_218), .B(n_248), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_218), .B(n_285), .Y(n_373) );
AND2x4_ASAP7_75t_L g430 ( .A(n_218), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_236), .Y(n_218) );
INVx2_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
AND2x2_ASAP7_75t_L g332 ( .A(n_219), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_R g350 ( .A(n_219), .Y(n_350) );
INVx2_ASAP7_75t_L g392 ( .A(n_219), .Y(n_392) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_219), .Y(n_409) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_232), .B(n_233), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g227 ( .A(n_223), .Y(n_227) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
INVx2_ASAP7_75t_L g583 ( .A(n_223), .Y(n_583) );
INVx2_ASAP7_75t_L g646 ( .A(n_223), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_232), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g579 ( .A(n_232), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_237), .Y(n_284) );
AND2x2_ASAP7_75t_L g391 ( .A(n_237), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AND2x2_ASAP7_75t_L g299 ( .A(n_238), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
OAI221xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_260), .B1(n_281), .B2(n_287), .C(n_292), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_257), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_248), .B(n_350), .Y(n_428) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_248), .Y(n_491) );
AND2x2_ASAP7_75t_L g285 ( .A(n_249), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_249), .B(n_258), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_249), .B(n_439), .Y(n_504) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g298 ( .A(n_251), .B(n_299), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_253), .A2(n_268), .B(n_271), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_253), .A2(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g434 ( .A(n_257), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g494 ( .A(n_257), .B(n_365), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_257), .B(n_351), .Y(n_524) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g458 ( .A(n_258), .B(n_317), .Y(n_458) );
AND2x2_ASAP7_75t_L g379 ( .A(n_259), .B(n_333), .Y(n_379) );
INVx1_ASAP7_75t_SL g401 ( .A(n_259), .Y(n_401) );
INVx1_ASAP7_75t_L g440 ( .A(n_259), .Y(n_440) );
BUFx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_261), .B(n_383), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_277), .Y(n_261) );
INVx2_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
INVx2_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
INVx2_ASAP7_75t_L g326 ( .A(n_263), .Y(n_326) );
INVx1_ASAP7_75t_L g366 ( .A(n_263), .Y(n_366) );
AND2x2_ASAP7_75t_L g406 ( .A(n_263), .B(n_372), .Y(n_406) );
OR2x2_ASAP7_75t_L g477 ( .A(n_263), .B(n_328), .Y(n_477) );
BUFx2_ASAP7_75t_L g484 ( .A(n_263), .Y(n_484) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_275), .Y(n_264) );
AND2x4_ASAP7_75t_L g384 ( .A(n_277), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_277), .B(n_341), .Y(n_397) );
INVx3_ASAP7_75t_L g407 ( .A(n_277), .Y(n_407) );
AND2x2_ASAP7_75t_L g441 ( .A(n_277), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g518 ( .A(n_277), .B(n_338), .Y(n_518) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g308 ( .A(n_278), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_278), .B(n_307), .Y(n_318) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g346 ( .A(n_279), .Y(n_346) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_282), .B(n_384), .Y(n_444) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
OR2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_320), .Y(n_319) );
NOR4xp25_ASAP7_75t_L g382 ( .A(n_283), .B(n_359), .C(n_383), .D(n_386), .Y(n_382) );
OR2x2_ASAP7_75t_L g469 ( .A(n_283), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g509 ( .A(n_286), .B(n_448), .Y(n_509) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_289), .B(n_345), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g451 ( .A(n_290), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_SL g354 ( .A1(n_293), .A2(n_355), .B(n_357), .C(n_361), .Y(n_354) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g462 ( .A(n_294), .B(n_336), .Y(n_462) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_295), .A2(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_303), .Y(n_296) );
OR2x2_ASAP7_75t_L g330 ( .A(n_297), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g459 ( .A(n_297), .Y(n_459) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g415 ( .A(n_298), .B(n_392), .Y(n_415) );
INVx1_ASAP7_75t_L g448 ( .A(n_298), .Y(n_448) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g615 ( .A(n_302), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_302), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g500 ( .A(n_303), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_309), .B(n_311), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g339 ( .A1(n_306), .A2(n_340), .A3(n_341), .B1(n_344), .B2(n_347), .Y(n_339) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g479 ( .A(n_309), .Y(n_479) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g442 ( .A(n_310), .B(n_326), .Y(n_442) );
OAI322xp33_ASAP7_75t_L g519 ( .A1(n_311), .A2(n_372), .A3(n_377), .B1(n_474), .B2(n_484), .C1(n_520), .C2(n_523), .Y(n_519) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_339), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_319), .B(n_321), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx2_ASAP7_75t_L g497 ( .A(n_324), .Y(n_497) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
AND2x2_ASAP7_75t_L g465 ( .A(n_326), .B(n_346), .Y(n_465) );
AND2x2_ASAP7_75t_L g505 ( .A(n_327), .B(n_407), .Y(n_505) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g480 ( .A(n_332), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g390 ( .A(n_333), .Y(n_390) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g356 ( .A(n_337), .Y(n_356) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g377 ( .A(n_343), .B(n_346), .Y(n_377) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_346), .B(n_370), .Y(n_496) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g437 ( .A(n_352), .B(n_438), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_363), .C(n_374), .D(n_382), .Y(n_353) );
INVx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_358), .A2(n_425), .B1(n_426), .B2(n_429), .C(n_433), .Y(n_424) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_360), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_368), .B(n_373), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_366), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_379), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g503 ( .A(n_379), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g470 ( .A(n_381), .B(n_390), .Y(n_470) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_407), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_385), .B(n_407), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_385), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_385), .B(n_484), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_385), .B(n_464), .Y(n_502) );
INVx1_ASAP7_75t_SL g510 ( .A(n_385), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_386), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g435 ( .A(n_386), .Y(n_435) );
INVx1_ASAP7_75t_L g492 ( .A(n_386), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B(n_394), .C(n_410), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g487 ( .A(n_391), .Y(n_487) );
INVx1_ASAP7_75t_L g439 ( .A(n_392), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_405), .C(n_407), .D(n_408), .Y(n_398) );
OR2x2_ASAP7_75t_L g402 ( .A(n_401), .B(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_403), .Y(n_423) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g450 ( .A(n_406), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g476 ( .A(n_407), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_432), .Y(n_474) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g490 ( .A(n_411), .Y(n_490) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_413), .B(n_468), .Y(n_467) );
AOI21xp33_ASAP7_75t_SL g463 ( .A1(n_414), .A2(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_452), .C(n_506), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_424), .C(n_443), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_429), .A2(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g486 ( .A(n_432), .B(n_487), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B(n_441), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_436), .A2(n_502), .B1(n_503), .B2(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_471), .C(n_488), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_467), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_459), .B1(n_460), .B2(n_461), .C(n_463), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g513 ( .A(n_470), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_478), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_482), .B2(n_485), .Y(n_478) );
AND2x4_ASAP7_75t_L g499 ( .A(n_481), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_493), .B1(n_495), .B2(n_498), .C(n_501), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .C(n_519), .Y(n_506) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_514), .B(n_517), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_525), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_533), .A2(n_542), .B(n_951), .Y(n_541) );
BUFx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
CKINVDCx6p67_ASAP7_75t_R g954 ( .A(n_540), .Y(n_954) );
XOR2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .Y(n_543) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_941), .B1(n_942), .B2(n_944), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_831), .Y(n_554) );
NOR4xp75_ASAP7_75t_SL g555 ( .A(n_556), .B(n_749), .C(n_795), .D(n_815), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_720), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_616), .B(n_622), .C(n_682), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g896 ( .A1(n_558), .A2(n_863), .B1(n_897), .B2(n_900), .C1(n_904), .C2(n_910), .Y(n_896) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_576), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g684 ( .A(n_560), .B(n_594), .Y(n_684) );
INVx1_ASAP7_75t_L g732 ( .A(n_560), .Y(n_732) );
INVx1_ASAP7_75t_L g861 ( .A(n_560), .Y(n_861) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g700 ( .A(n_561), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g723 ( .A(n_561), .Y(n_723) );
OR2x2_ASAP7_75t_L g755 ( .A(n_561), .B(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g798 ( .A(n_561), .B(n_701), .Y(n_798) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_561), .Y(n_805) );
AND2x2_ASAP7_75t_L g865 ( .A(n_561), .B(n_756), .Y(n_865) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .A3(n_569), .B(n_574), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_567), .B(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_568), .A2(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g760 ( .A(n_576), .Y(n_760) );
INVx1_ASAP7_75t_L g940 ( .A(n_576), .Y(n_940) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_594), .Y(n_576) );
AND2x2_ASAP7_75t_L g685 ( .A(n_577), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g807 ( .A(n_577), .B(n_702), .Y(n_807) );
INVx2_ASAP7_75t_L g812 ( .A(n_577), .Y(n_812) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B(n_593), .Y(n_578) );
OAI21x1_ASAP7_75t_L g719 ( .A1(n_579), .A2(n_592), .B(n_715), .Y(n_719) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_580), .A2(n_593), .B(n_620), .Y(n_619) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_586), .B(n_591), .Y(n_580) );
INVx1_ASAP7_75t_L g659 ( .A(n_583), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_585), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_591), .B(n_641), .Y(n_663) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g778 ( .A(n_594), .B(n_619), .Y(n_778) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g618 ( .A(n_595), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_595), .B(n_861), .Y(n_860) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g686 ( .A(n_596), .Y(n_686) );
INVx1_ASAP7_75t_L g745 ( .A(n_596), .Y(n_745) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_605), .B(n_614), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_604), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_604), .B(n_658), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_608), .B(n_613), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_606), .A2(n_644), .B1(n_647), .B2(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_610), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_610), .B(n_678), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_616), .A2(n_853), .B(n_854), .Y(n_852) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp67_ASAP7_75t_L g783 ( .A(n_617), .B(n_700), .Y(n_783) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g724 ( .A(n_618), .Y(n_724) );
AND2x2_ASAP7_75t_L g733 ( .A(n_619), .B(n_702), .Y(n_733) );
BUFx2_ASAP7_75t_L g830 ( .A(n_619), .Y(n_830) );
OR2x2_ASAP7_75t_L g875 ( .A(n_619), .B(n_755), .Y(n_875) );
OA21x2_ASAP7_75t_L g691 ( .A1(n_620), .A2(n_651), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_621), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_652), .Y(n_623) );
INVx1_ASAP7_75t_L g872 ( .A(n_624), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_639), .Y(n_624) );
AND2x4_ASAP7_75t_L g694 ( .A(n_625), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g728 ( .A(n_625), .B(n_666), .Y(n_728) );
BUFx2_ASAP7_75t_SL g736 ( .A(n_625), .Y(n_736) );
INVx1_ASAP7_75t_L g748 ( .A(n_625), .Y(n_748) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2x1_ASAP7_75t_L g767 ( .A(n_626), .B(n_727), .Y(n_767) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g786 ( .A(n_627), .Y(n_786) );
AO31x2_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_632), .A3(n_637), .B(n_638), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_631), .A2(n_661), .B(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g712 ( .A(n_636), .Y(n_712) );
AND2x2_ASAP7_75t_L g814 ( .A(n_639), .B(n_743), .Y(n_814) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g726 ( .A(n_640), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g851 ( .A(n_640), .B(n_654), .Y(n_851) );
AOI21x1_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_650), .Y(n_640) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2x1_ASAP7_75t_L g834 ( .A(n_652), .B(n_835), .Y(n_834) );
OR2x2_ASAP7_75t_L g889 ( .A(n_652), .B(n_736), .Y(n_889) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_653), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g792 ( .A(n_653), .B(n_736), .Y(n_792) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_666), .Y(n_653) );
AND2x2_ASAP7_75t_L g738 ( .A(n_654), .B(n_691), .Y(n_738) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g743 ( .A(n_655), .Y(n_743) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g727 ( .A(n_656), .Y(n_727) );
AOI21x1_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B(n_664), .Y(n_656) );
NOR2x1_ASAP7_75t_L g873 ( .A(n_666), .B(n_727), .Y(n_873) );
OA21x2_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B(n_679), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g695 ( .A(n_680), .B(n_696), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_693), .B2(n_698), .Y(n_682) );
NOR2xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_684), .B(n_794), .Y(n_931) );
AND2x2_ASAP7_75t_L g699 ( .A(n_685), .B(n_700), .Y(n_699) );
NAND2x1_ASAP7_75t_SL g817 ( .A(n_685), .B(n_805), .Y(n_817) );
INVx2_ASAP7_75t_SL g754 ( .A(n_686), .Y(n_754) );
AND2x2_ASAP7_75t_L g887 ( .A(n_686), .B(n_701), .Y(n_887) );
BUFx2_ASAP7_75t_L g934 ( .A(n_686), .Y(n_934) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_688), .A2(n_826), .B(n_827), .C(n_829), .Y(n_825) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2x1p5_ASAP7_75t_L g766 ( .A(n_690), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g782 ( .A(n_690), .Y(n_782) );
INVx2_ASAP7_75t_L g907 ( .A(n_690), .Y(n_907) );
INVx1_ASAP7_75t_L g911 ( .A(n_690), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_690), .B(n_901), .Y(n_924) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g774 ( .A(n_691), .Y(n_774) );
INVx1_ASAP7_75t_L g836 ( .A(n_691), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_691), .B(n_786), .Y(n_856) );
OR2x2_ASAP7_75t_L g898 ( .A(n_693), .B(n_899), .Y(n_898) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g770 ( .A(n_694), .B(n_726), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_694), .B(n_821), .Y(n_820) );
AND2x4_ASAP7_75t_L g880 ( .A(n_694), .B(n_850), .Y(n_880) );
AND2x2_ASAP7_75t_L g915 ( .A(n_694), .B(n_742), .Y(n_915) );
INVx1_ASAP7_75t_L g764 ( .A(n_695), .Y(n_764) );
NOR2x1_ASAP7_75t_L g773 ( .A(n_695), .B(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g785 ( .A(n_695), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_695), .B(n_929), .Y(n_928) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g853 ( .A(n_700), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_701), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI21x1_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_710), .B(n_719), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_703), .A2(n_710), .B(n_719), .Y(n_756) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_706), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND3x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .C(n_716), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_725), .B1(n_729), .B2(n_734), .C(n_739), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_722), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx2_ASAP7_75t_SL g777 ( .A(n_723), .Y(n_777) );
AND2x4_ASAP7_75t_L g842 ( .A(n_723), .B(n_733), .Y(n_842) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_723), .Y(n_901) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
AND2x2_ASAP7_75t_L g803 ( .A(n_726), .B(n_736), .Y(n_803) );
AND2x2_ASAP7_75t_L g933 ( .A(n_726), .B(n_934), .Y(n_933) );
AND2x6_ASAP7_75t_SL g937 ( .A(n_726), .B(n_824), .Y(n_937) );
INVx1_ASAP7_75t_L g828 ( .A(n_727), .Y(n_828) );
AND2x2_ASAP7_75t_L g781 ( .A(n_728), .B(n_782), .Y(n_781) );
AND2x4_ASAP7_75t_L g849 ( .A(n_728), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g936 ( .A(n_728), .Y(n_936) );
NOR4xp25_ASAP7_75t_L g739 ( .A(n_730), .B(n_740), .C(n_744), .D(n_746), .Y(n_739) );
INVx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g883 ( .A(n_731), .B(n_844), .Y(n_883) );
AND2x4_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_733), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g794 ( .A(n_733), .Y(n_794) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g784 ( .A(n_738), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g899 ( .A(n_738), .Y(n_899) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_741), .B(n_746), .Y(n_923) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g821 ( .A(n_743), .Y(n_821) );
INVx1_ASAP7_75t_L g929 ( .A(n_743), .Y(n_929) );
OR2x2_ASAP7_75t_L g854 ( .A(n_744), .B(n_798), .Y(n_854) );
AND2x2_ASAP7_75t_L g891 ( .A(n_744), .B(n_892), .Y(n_891) );
INVx2_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g789 ( .A(n_745), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_746), .A2(n_755), .B1(n_759), .B2(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g813 ( .A(n_748), .B(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_750), .B(n_779), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_757), .B(n_761), .C(n_768), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
AND2x2_ASAP7_75t_L g848 ( .A(n_753), .B(n_807), .Y(n_848) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g806 ( .A(n_754), .B(n_807), .Y(n_806) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_754), .Y(n_839) );
INVx1_ASAP7_75t_L g867 ( .A(n_754), .Y(n_867) );
OR2x2_ASAP7_75t_L g939 ( .A(n_755), .B(n_940), .Y(n_939) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_756), .Y(n_759) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx2_ASAP7_75t_L g826 ( .A(n_759), .Y(n_826) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
AND2x2_ASAP7_75t_L g791 ( .A(n_763), .B(n_766), .Y(n_791) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_764), .B(n_824), .Y(n_847) );
AND2x2_ASAP7_75t_L g920 ( .A(n_764), .B(n_821), .Y(n_920) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g771 ( .A(n_767), .B(n_772), .Y(n_771) );
AOI21xp33_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_771), .B(n_775), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_769), .A2(n_856), .B1(n_857), .B2(n_862), .Y(n_855) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_770), .A2(n_865), .B1(n_866), .B2(n_870), .C(n_874), .Y(n_864) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g823 ( .A(n_773), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
OR2x2_ASAP7_75t_L g810 ( .A(n_777), .B(n_811), .Y(n_810) );
OR2x6_ASAP7_75t_L g868 ( .A(n_777), .B(n_869), .Y(n_868) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_778), .Y(n_878) );
INVx1_ASAP7_75t_L g903 ( .A(n_778), .Y(n_903) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_790), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B1(n_784), .B2(n_787), .Y(n_780) );
INVx1_ASAP7_75t_L g840 ( .A(n_781), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_785), .B(n_821), .Y(n_838) );
AND2x2_ASAP7_75t_L g910 ( .A(n_785), .B(n_911), .Y(n_910) );
BUFx3_ASAP7_75t_L g824 ( .A(n_786), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_787), .A2(n_834), .B(n_837), .Y(n_833) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g800 ( .A(n_791), .Y(n_800) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_808), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_799), .B1(n_801), .B2(n_804), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_797), .A2(n_910), .B1(n_915), .B2(n_916), .Y(n_914) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVxp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI21xp5_ASAP7_75t_SL g808 ( .A1(n_804), .A2(n_809), .B(n_813), .Y(n_808) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx2_ASAP7_75t_L g859 ( .A(n_807), .Y(n_859) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g892 ( .A(n_811), .Y(n_892) );
BUFx2_ASAP7_75t_SL g869 ( .A(n_812), .Y(n_869) );
INVx1_ASAP7_75t_L g886 ( .A(n_812), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_818), .B(n_825), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g827 ( .A(n_823), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_824), .B(n_873), .Y(n_909) );
INVx1_ASAP7_75t_L g916 ( .A(n_826), .Y(n_916) );
INVxp67_ASAP7_75t_L g845 ( .A(n_828), .Y(n_845) );
AOI21xp33_ASAP7_75t_L g922 ( .A1(n_829), .A2(n_923), .B(n_924), .Y(n_922) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_830), .A2(n_919), .B(n_921), .Y(n_918) );
NOR3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_881), .C(n_912), .Y(n_831) );
NAND3xp33_ASAP7_75t_SL g832 ( .A(n_833), .B(n_843), .C(n_864), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2x1_ASAP7_75t_L g894 ( .A(n_836), .B(n_895), .Y(n_894) );
O2A1O1Ixp33_ASAP7_75t_SL g837 ( .A1(n_838), .A2(n_839), .B(n_840), .C(n_841), .Y(n_837) );
INVx1_ASAP7_75t_L g913 ( .A(n_839), .Y(n_913) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_848), .B1(n_849), .B2(n_852), .C(n_855), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g926 ( .A(n_856), .Y(n_926) );
INVx2_ASAP7_75t_SL g857 ( .A(n_858), .Y(n_857) );
NOR2x1_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g863 ( .A(n_859), .Y(n_863) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g877 ( .A(n_865), .Y(n_877) );
NOR2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B(n_879), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_890), .C(n_896), .Y(n_881) );
NOR2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NOR2x1_ASAP7_75t_L g884 ( .A(n_885), .B(n_888), .Y(n_884) );
NAND2x1p5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g921 ( .A(n_887), .Y(n_921) );
BUFx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g895 ( .A(n_889), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
AND2x4_ASAP7_75t_L g904 ( .A(n_905), .B(n_908), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI211xp5_ASAP7_75t_SL g912 ( .A1(n_913), .A2(n_914), .B(n_917), .C(n_932), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_922), .B1(n_925), .B2(n_930), .Y(n_917) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AND2x2_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVxp33_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_935), .B1(n_937), .B2(n_938), .Y(n_932) );
INVxp67_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
BUFx8_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_952), .Y(n_951) );
BUFx8_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_956), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_957), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_957), .Y(n_965) );
BUFx8_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
BUFx5_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
endmodule