module real_jpeg_19699_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_0),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_0),
.A2(n_46),
.B1(n_48),
.B2(n_124),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_124),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_124),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_57),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_34),
.B1(n_46),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_2),
.A2(n_34),
.B1(n_64),
.B2(n_65),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_119),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_119),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_119),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_4),
.A2(n_22),
.B1(n_64),
.B2(n_65),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_4),
.A2(n_22),
.B1(n_46),
.B2(n_48),
.Y(n_284)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_6),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_88),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_46),
.B1(n_48),
.B2(n_88),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_88),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_7),
.A2(n_48),
.B(n_60),
.C(n_104),
.D(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_45),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_7),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_125),
.B(n_127),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_31),
.B(n_42),
.C(n_164),
.D(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_7),
.B(n_31),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_7),
.B(n_35),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_7),
.A2(n_32),
.B(n_204),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_143),
.Y(n_221)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_10),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_12),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_107),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_107),
.Y(n_224)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_338),
.B(n_341),
.Y(n_17)
);

OAI21x1_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_74),
.B(n_337),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_20),
.B(n_36),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_20),
.B(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_20),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_23),
.A2(n_28),
.B(n_143),
.C(n_203),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_26),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_26),
.B(n_224),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_340)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_27),
.A2(n_30),
.B1(n_232),
.B2(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_27),
.A2(n_223),
.B(n_261),
.Y(n_279)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_30),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_30),
.A2(n_87),
.B(n_233),
.Y(n_303)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_35),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_69),
.C(n_71),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_38),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_41),
.A2(n_50),
.B1(n_183),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_41),
.A2(n_218),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_45),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_42),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_42),
.A2(n_45),
.B1(n_258),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_42),
.A2(n_45),
.B1(n_93),
.B2(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_44),
.Y(n_172)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_46),
.B(n_47),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_48),
.A2(n_164),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_50),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_50),
.A2(n_184),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_53),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_58),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_59),
.A2(n_67),
.B1(n_118),
.B2(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_59),
.A2(n_162),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_59),
.A2(n_67),
.B1(n_215),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_59),
.A2(n_67),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_59),
.A2(n_67),
.B1(n_252),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_60),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_60),
.A2(n_63),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_64),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g125 ( 
.A(n_64),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_67),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_67),
.A2(n_120),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_94),
.B(n_336),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_76),
.B(n_80),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.C(n_89),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_86),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_86),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_89),
.B(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_319),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_345),
.Y(n_94)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_269),
.A3(n_307),
.B1(n_313),
.B2(n_318),
.C(n_346),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_226),
.C(n_265),
.Y(n_96)
);

AOI21x1_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_196),
.B(n_225),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_177),
.B(n_195),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_156),
.B(n_176),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_131),
.B(n_155),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_102),
.B(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_108),
.B1(n_109),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_105),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_117),
.C(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_125),
.B(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_125),
.A2(n_126),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_125),
.A2(n_152),
.B1(n_208),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_125),
.A2(n_145),
.B1(n_241),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_125),
.A2(n_126),
.B(n_250),
.Y(n_282)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_147),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_130),
.A2(n_136),
.B1(n_174),
.B2(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_140),
.B(n_154),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_148),
.B(n_153),
.Y(n_140)
);

NOR2x1_ASAP7_75t_R g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_158),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_169),
.B2(n_175),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_168),
.C(n_175),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_191),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_192),
.C(n_193),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_186),
.B2(n_190),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_187),
.C(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_198),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_212),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_211),
.C(n_212),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_220),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_227),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_245),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_228),
.B(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_239),
.C(n_244),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_242),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_263),
.B2(n_264),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_253),
.C(n_264),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_259),
.C(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_267),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_287),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_270),
.B(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.C(n_286),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_271),
.A2(n_272),
.B1(n_280),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_282),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_299),
.B(n_303),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_283),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_305),
.B2(n_306),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_298),
.C(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B(n_296),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_296),
.A2(n_321),
.B1(n_325),
.B2(n_333),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule