module fake_jpeg_1539_n_109 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_37),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_31),
.B(n_37),
.C(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_32),
.B1(n_38),
.B2(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_41),
.B1(n_33),
.B2(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_1),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_43),
.B(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_56),
.B1(n_50),
.B2(n_43),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_12),
.B1(n_25),
.B2(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_2),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_75),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_62),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_88),
.C(n_89),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_14),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_27),
.B(n_20),
.C(n_17),
.D(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_3),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_3),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_4),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_11),
.C(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_98),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_82),
.B(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_93),
.B1(n_95),
.B2(n_92),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_93),
.C(n_99),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_97),
.C(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_8),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.C(n_9),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_10),
.CI(n_84),
.CON(n_109),
.SN(n_109)
);


endmodule