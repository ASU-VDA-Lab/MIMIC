module fake_jpeg_25411_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_26),
.Y(n_45)
);

BUFx2_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_26),
.C(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_50),
.B1(n_55),
.B2(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_33),
.B1(n_38),
.B2(n_19),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_26),
.C(n_22),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_23),
.B1(n_16),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_23),
.B1(n_16),
.B2(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_19),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_17),
.B(n_28),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_78),
.B1(n_50),
.B2(n_58),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_65),
.B1(n_69),
.B2(n_58),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_21),
.B1(n_33),
.B2(n_40),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_72),
.B1(n_81),
.B2(n_44),
.Y(n_107)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_71),
.Y(n_88)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_31),
.B1(n_19),
.B2(n_28),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_28),
.B1(n_38),
.B2(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_38),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_45),
.B(n_0),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_90),
.B(n_108),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_41),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_70),
.B1(n_42),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_99),
.B1(n_65),
.B2(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_100),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_50),
.C(n_47),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_110),
.C(n_39),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_107),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_22),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_57),
.B1(n_56),
.B2(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_44),
.B1(n_57),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_77),
.B1(n_56),
.B2(n_43),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_1),
.B(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_34),
.C(n_39),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_130),
.B1(n_105),
.B2(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_116),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_25),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_34),
.Y(n_119)
);

NAND2xp67_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_34),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_128),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_131),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_83),
.B(n_37),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_25),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_134),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_89),
.B(n_22),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_67),
.B1(n_30),
.B2(n_37),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_153),
.Y(n_175)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_158),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_107),
.B1(n_106),
.B2(n_100),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_103),
.B1(n_64),
.B2(n_85),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_161),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_95),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_101),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_121),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_98),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_110),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_124),
.B(n_120),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_180),
.B(n_140),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_124),
.B1(n_115),
.B2(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_183),
.C(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_115),
.B1(n_130),
.B2(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_184),
.B2(n_187),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_115),
.B1(n_112),
.B2(n_108),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_129),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_102),
.B(n_109),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_67),
.B1(n_30),
.B2(n_48),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_140),
.B1(n_138),
.B2(n_146),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_67),
.B1(n_30),
.B2(n_18),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_25),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_160),
.C(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_148),
.B1(n_145),
.B2(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_150),
.B(n_138),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_210),
.B(n_154),
.Y(n_214)
);

NOR4xp25_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_162),
.C(n_157),
.D(n_161),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_187),
.B1(n_179),
.B2(n_188),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_137),
.B1(n_151),
.B2(n_142),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_9),
.B1(n_2),
.B2(n_4),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_170),
.B1(n_176),
.B2(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_207),
.B1(n_174),
.B2(n_185),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

BUFx4f_ASAP7_75t_SL g209 ( 
.A(n_185),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_180),
.B(n_173),
.C(n_186),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_157),
.B(n_177),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_224),
.B1(n_195),
.B2(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_191),
.B1(n_194),
.B2(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_168),
.C(n_147),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_222),
.C(n_223),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_197),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_147),
.C(n_30),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_9),
.C(n_2),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_196),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_204),
.C(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_237),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_210),
.C(n_197),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_194),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_238),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_215),
.B1(n_224),
.B2(n_221),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_220),
.B(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_236),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_221),
.B(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_10),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_243),
.Y(n_261)
);

NAND4xp25_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_237),
.C(n_213),
.D(n_231),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_246),
.A3(n_248),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_256),
.B(n_13),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_209),
.B1(n_2),
.B2(n_5),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_10),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_12),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_15),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_257)
);

NAND2x1_ASAP7_75t_SL g258 ( 
.A(n_257),
.B(n_13),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_252),
.B1(n_6),
.B2(n_11),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_259),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_267),
.B(n_262),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_264),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_248),
.B(n_14),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_14),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_1),
.B1(n_15),
.B2(n_262),
.Y(n_273)
);


endmodule