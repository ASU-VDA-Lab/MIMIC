module real_jpeg_11837_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_69),
.B1(n_71),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_3),
.A2(n_50),
.B1(n_54),
.B2(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_89),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_5),
.A2(n_50),
.B1(n_54),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_69),
.B1(n_71),
.B2(n_77),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_50),
.B1(n_54),
.B2(n_57),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_7),
.A2(n_57),
.B1(n_69),
.B2(n_71),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_9),
.A2(n_44),
.B1(n_69),
.B2(n_71),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_69),
.B1(n_71),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_10),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_10),
.A2(n_50),
.B1(n_54),
.B2(n_91),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_91),
.Y(n_306)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_30),
.B(n_36),
.C(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_12),
.B(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_31),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_12),
.A2(n_31),
.B(n_142),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_65),
.C(n_71),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_41),
.B1(n_50),
.B2(n_54),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_85),
.B1(n_86),
.B2(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_12),
.B(n_113),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_13),
.A2(n_50),
.B1(n_54),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_74),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_13),
.A2(n_69),
.B1(n_71),
.B2(n_74),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_74),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_14),
.A2(n_50),
.B1(n_54),
.B2(n_59),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_59),
.B1(n_69),
.B2(n_71),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_59),
.Y(n_223)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_322),
.C(n_326),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_320),
.B(n_324),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_313),
.B(n_319),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_279),
.B(n_310),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_257),
.B(n_278),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_230),
.B(n_256),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_125),
.B(n_206),
.C(n_229),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_104),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_24),
.B(n_104),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_80),
.C(n_95),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_25),
.B(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_60),
.C(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_27),
.B(n_275),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_27),
.A2(n_45),
.B(n_252),
.Y(n_326)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_28),
.A2(n_29),
.B1(n_43),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_28),
.A2(n_29),
.B1(n_108),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_28),
.A2(n_223),
.B(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_28),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_28),
.A2(n_29),
.B1(n_291),
.B2(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_28),
.A2(n_274),
.B(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_29),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_32),
.B1(n_52),
.B2(n_53),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_31),
.A2(n_34),
.B(n_41),
.Y(n_94)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_SL g143 ( 
.A(n_32),
.B(n_52),
.C(n_54),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_41),
.B(n_86),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_41),
.B(n_68),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_45),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_45),
.B(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_60),
.B1(n_61),
.B2(n_79),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_48),
.A2(n_58),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_48),
.A2(n_49),
.B1(n_103),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_48),
.A2(n_112),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_48),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_48),
.A2(n_225),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_49),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_50),
.A2(n_53),
.B(n_141),
.C(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_72),
.B(n_75),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_62),
.A2(n_68),
.B(n_72),
.Y(n_288)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_63),
.A2(n_78),
.B1(n_136),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_63),
.A2(n_78),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_63),
.A2(n_78),
.B1(n_159),
.B2(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_63),
.A2(n_78),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_63),
.A2(n_216),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_69),
.B(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_78),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_75),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_81),
.B1(n_95),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_84),
.A2(n_123),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_84),
.A2(n_87),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_85),
.A2(n_86),
.B1(n_172),
.B2(n_180),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_85),
.A2(n_174),
.B(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_85),
.A2(n_86),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_99),
.Y(n_123)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_88),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_87),
.B(n_146),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_98),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_105),
.B(n_116),
.C(n_124),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_114),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_109),
.C(n_114),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_110),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_111),
.A2(n_113),
.B(n_249),
.Y(n_316)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_113),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_113),
.A2(n_249),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_117),
.B(n_120),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_118),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_119),
.B(n_137),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_204),
.B(n_205),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_147),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_131),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_138),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_160),
.B(n_203),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_152),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_197),
.B(n_202),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_186),
.B(n_196),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_175),
.B(n_185),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_170),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_167),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_184),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_188),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_192),
.C(n_195),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_201),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_228),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_228),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_210),
.C(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_217),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_221),
.C(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_227),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_255),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_241),
.B1(n_253),
.B2(n_254),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_254),
.C(n_255),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_236),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_238),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_236),
.A2(n_269),
.B(n_271),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_246),
.C(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_292),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_277),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_277),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_276),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_262),
.C(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_266),
.B(n_267),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_282),
.C(n_294),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_282),
.CI(n_294),
.CON(n_309),
.SN(n_309)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_307),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_295),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_295),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_290),
.B2(n_293),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_289),
.C(n_290),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_289),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_302),
.C(n_304),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_293),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_296),
.C(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_309),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_315),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_322),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.CI(n_318),
.CON(n_315),
.SN(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule