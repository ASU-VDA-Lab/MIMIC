module fake_jpeg_5823_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_16),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_47),
.B1(n_50),
.B2(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_18),
.B1(n_17),
.B2(n_21),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_15),
.Y(n_51)
);

AOI32xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_39),
.A3(n_31),
.B1(n_15),
.B2(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_39),
.B1(n_33),
.B2(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_63),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_48),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_20),
.B(n_22),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_44),
.B(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_43),
.C(n_49),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_73),
.C(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_48),
.B1(n_56),
.B2(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_15),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_40),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_46),
.C(n_31),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_64),
.B1(n_62),
.B2(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_79),
.B1(n_12),
.B2(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_56),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_15),
.B(n_12),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_67),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_89),
.B(n_85),
.C(n_90),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_29),
.B1(n_38),
.B2(n_36),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_76),
.B1(n_38),
.B2(n_36),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_87),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_91),
.B(n_92),
.C(n_7),
.D(n_5),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_7),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_2),
.C2(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_99),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_3),
.C(n_6),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_3),
.C(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_40),
.B(n_6),
.Y(n_108)
);


endmodule