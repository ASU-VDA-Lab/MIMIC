module fake_netlist_1_5960_n_460 (n_117, n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_124, n_120, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_122, n_126, n_118, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_460);
input n_117;
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_120;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_122;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_460;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_457;
wire n_223;
wire n_453;
wire n_372;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g128 ( .A(n_61), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_109), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_79), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_25), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
INVxp67_ASAP7_75t_SL g133 ( .A(n_113), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_66), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_38), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_99), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_14), .B(n_47), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_120), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_101), .Y(n_144) );
CKINVDCx14_ASAP7_75t_R g145 ( .A(n_27), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_2), .Y(n_147) );
INVx1_ASAP7_75t_SL g148 ( .A(n_112), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_110), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_80), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_54), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_78), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_58), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_76), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_0), .B(n_90), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_60), .Y(n_158) );
INVxp67_ASAP7_75t_SL g159 ( .A(n_98), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_65), .Y(n_160) );
INVxp67_ASAP7_75t_SL g161 ( .A(n_40), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_62), .Y(n_162) );
INVxp67_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_26), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_82), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g166 ( .A(n_127), .Y(n_166) );
CKINVDCx14_ASAP7_75t_R g167 ( .A(n_36), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_83), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_53), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_10), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_37), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_67), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_20), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_105), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_69), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_11), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_81), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_73), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_126), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_21), .Y(n_180) );
NOR2xp67_ASAP7_75t_L g181 ( .A(n_122), .B(n_86), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_30), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_97), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_125), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_121), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_102), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_19), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_4), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_35), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_41), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_117), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_119), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_123), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_4), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_72), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_115), .Y(n_197) );
INVxp33_ASAP7_75t_SL g198 ( .A(n_44), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_45), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_0), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_55), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_70), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_59), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_75), .B(n_107), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_71), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_13), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_118), .Y(n_207) );
NOR2xp67_ASAP7_75t_L g208 ( .A(n_84), .B(n_49), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_2), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_100), .Y(n_210) );
INVxp67_ASAP7_75t_SL g211 ( .A(n_42), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_103), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_91), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_77), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_185), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_200), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_170), .B(n_1), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_206), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_147), .B(n_1), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_195), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_134), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_185), .B(n_209), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_166), .B(n_3), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_137), .B(n_3), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_142), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_143), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_152), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_146), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_162), .B(n_5), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_233), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_233), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_235), .B(n_214), .Y(n_238) );
NOR2x1p5_ASAP7_75t_L g239 ( .A(n_219), .B(n_133), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_221), .B(n_153), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_223), .B(n_175), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_217), .B(n_191), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_229), .B(n_213), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_216), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_224), .B(n_128), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_218), .B(n_163), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_230), .B(n_145), .Y(n_249) );
CKINVDCx11_ASAP7_75t_R g250 ( .A(n_240), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_240), .B(n_226), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_249), .A2(n_225), .B(n_227), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_238), .B(n_231), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_244), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_241), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_244), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_236), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_245), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_248), .B(n_220), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_243), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_242), .B(n_232), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_255), .B(n_248), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_239), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_260), .B(n_131), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_261), .B(n_238), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_251), .B(n_238), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_252), .A2(n_247), .B(n_235), .C(n_234), .Y(n_268) );
CKINVDCx8_ASAP7_75t_R g269 ( .A(n_250), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_256), .B(n_246), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_254), .B(n_198), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_259), .A2(n_161), .B(n_159), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_258), .B(n_138), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_264), .B(n_189), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_268), .A2(n_157), .B(n_154), .C(n_155), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_270), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_263), .B(n_129), .Y(n_278) );
AO22x2_ASAP7_75t_L g279 ( .A1(n_269), .A2(n_160), .B1(n_148), .B2(n_211), .Y(n_279) );
OAI22x1_ASAP7_75t_L g280 ( .A1(n_265), .A2(n_193), .B1(n_160), .B2(n_148), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_271), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_273), .A2(n_204), .B(n_257), .Y(n_282) );
AOI21xp33_ASAP7_75t_L g283 ( .A1(n_267), .A2(n_262), .B(n_179), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_272), .A2(n_186), .A3(n_158), .B(n_212), .Y(n_284) );
AO31x2_ASAP7_75t_L g285 ( .A1(n_274), .A2(n_182), .A3(n_171), .B(n_164), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_270), .Y(n_286) );
BUFx4_ASAP7_75t_SL g287 ( .A(n_269), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_268), .A2(n_169), .B(n_168), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_266), .A2(n_178), .B(n_172), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_264), .B(n_188), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_277), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_286), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_282), .A2(n_208), .B(n_181), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_289), .A2(n_192), .B(n_183), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_276), .A2(n_199), .B(n_194), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_288), .A2(n_202), .B(n_180), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_281), .B(n_201), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_284), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_284), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_203), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_280), .B(n_5), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_275), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_287), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_207), .B(n_140), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_288), .A2(n_228), .B(n_215), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_282), .A2(n_130), .B(n_139), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_141), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_277), .B(n_167), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_289), .A2(n_156), .B(n_228), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_290), .A2(n_174), .B1(n_210), .B2(n_205), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_289), .A2(n_197), .B(n_196), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_292), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_293), .A2(n_190), .B(n_187), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_313), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_302), .A2(n_184), .B(n_177), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_308), .A2(n_176), .B(n_173), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_314), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_6), .B(n_7), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_307), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_304), .B(n_8), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_301), .B(n_12), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_319), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_311), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_305), .B(n_144), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_165), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_149), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_295), .B(n_151), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_315), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_317), .B(n_18), .Y(n_345) );
INVxp33_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_291), .Y(n_349) );
AOI21xp5_ASAP7_75t_SL g350 ( .A1(n_296), .A2(n_22), .B(n_23), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_306), .B(n_24), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_292), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_292), .Y(n_353) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_293), .A2(n_28), .B(n_29), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_291), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_292), .B(n_31), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_335), .A2(n_32), .B(n_33), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_349), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_320), .B(n_34), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_332), .B(n_39), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_356), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_353), .B(n_43), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_348), .B(n_46), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_335), .A2(n_48), .B(n_50), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_322), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_323), .B(n_51), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_355), .B(n_52), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_357), .B(n_56), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_358), .B(n_57), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_331), .B(n_351), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_327), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_321), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_343), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_344), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_337), .B(n_63), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_354), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_321), .B(n_64), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_371), .B(n_340), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_362), .B(n_346), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_366), .B(n_324), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_373), .B(n_339), .Y(n_398) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_382), .B(n_350), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_363), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_377), .B(n_347), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_360), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_364), .B(n_347), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_384), .B(n_379), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_387), .B(n_345), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_384), .B(n_325), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_396), .B(n_386), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_403), .B(n_369), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_406), .B(n_388), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_409), .B(n_374), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_410), .B(n_374), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_416), .B(n_381), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_411), .B(n_389), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_392), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_395), .B(n_376), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_405), .Y(n_427) );
INVx3_ASAP7_75t_SL g428 ( .A(n_413), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_415), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_417), .B(n_407), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_429), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_428), .B(n_400), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_421), .B(n_402), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_418), .B(n_394), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_422), .B(n_401), .Y(n_435) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_420), .B(n_370), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_433), .A2(n_423), .B1(n_414), .B2(n_399), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_431), .B(n_426), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_431), .B(n_426), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_432), .B(n_424), .Y(n_440) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_433), .B(n_427), .Y(n_441) );
XOR2x2_ASAP7_75t_L g442 ( .A(n_434), .B(n_398), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g443 ( .A1(n_440), .A2(n_436), .A3(n_435), .B(n_430), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g444 ( .A1(n_441), .A2(n_391), .B(n_365), .C(n_425), .Y(n_444) );
OAI21xp33_ASAP7_75t_SL g445 ( .A1(n_437), .A2(n_419), .B(n_397), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_438), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g447 ( .A1(n_439), .A2(n_404), .A3(n_408), .B(n_412), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_442), .A2(n_404), .B(n_415), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_448), .B(n_446), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_443), .B(n_447), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_450), .A2(n_445), .B1(n_444), .B2(n_385), .Y(n_451) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_449), .B(n_359), .Y(n_452) );
XOR2x1_ASAP7_75t_L g453 ( .A(n_451), .B(n_341), .Y(n_453) );
XOR2xp5_ASAP7_75t_L g454 ( .A(n_453), .B(n_452), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_454), .B(n_342), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g456 ( .A1(n_455), .A2(n_390), .B1(n_372), .B2(n_359), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_456), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_457), .A2(n_68), .B(n_74), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_458), .A2(n_85), .B1(n_87), .B2(n_92), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_459), .A2(n_93), .B1(n_94), .B2(n_96), .Y(n_460) );
endmodule