module fake_jpeg_19037_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_2),
.B(n_24),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_97),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_71),
.B(n_47),
.C(n_46),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_66),
.B1(n_69),
.B2(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_105),
.B1(n_75),
.B2(n_61),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_58),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_65),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_56),
.B1(n_54),
.B2(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_52),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_119),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_117),
.Y(n_130)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_63),
.B1(n_6),
.B2(n_5),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_84),
.B1(n_52),
.B2(n_58),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_118),
.B1(n_55),
.B2(n_2),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_48),
.B1(n_73),
.B2(n_49),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_65),
.B1(n_60),
.B2(n_53),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_9),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_50),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_131),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_134),
.Y(n_138)
);

BUFx4f_ASAP7_75t_SL g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_127),
.B1(n_124),
.B2(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_143),
.B1(n_128),
.B2(n_134),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_116),
.B1(n_12),
.B2(n_15),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_142),
.C(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_138),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_143),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_11),
.C(n_19),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_28),
.B(n_29),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_31),
.C(n_34),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_36),
.B(n_38),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_40),
.Y(n_158)
);


endmodule