module fake_jpeg_2044_n_636 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_636);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_636;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_585;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_62),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_67),
.Y(n_182)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_126),
.Y(n_140)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_74),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_42),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_78),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_81),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_89),
.Y(n_142)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_36),
.B(n_9),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_54),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_20),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_123),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_207)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_10),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_22),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_145),
.B(n_149),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_54),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_26),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_156),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_26),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_157),
.B(n_161),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_46),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_46),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_162),
.B(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_168),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_73),
.B(n_45),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_73),
.B(n_30),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_174),
.B(n_176),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_67),
.B(n_47),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_175),
.B(n_202),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_45),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_178),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_106),
.B(n_52),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_197),
.C(n_208),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_110),
.A2(n_27),
.B1(n_51),
.B2(n_104),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_188),
.A2(n_193),
.B1(n_210),
.B2(n_213),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_114),
.B(n_47),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_200),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_104),
.A2(n_27),
.B1(n_51),
.B2(n_39),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_90),
.A2(n_48),
.B1(n_58),
.B2(n_30),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_207),
.B1(n_19),
.B2(n_8),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_98),
.B(n_51),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_103),
.B(n_48),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_91),
.B(n_58),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_93),
.B(n_31),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_108),
.A2(n_51),
.B1(n_59),
.B2(n_55),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_95),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_116),
.B(n_52),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_4),
.Y(n_273)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_39),
.B1(n_55),
.B2(n_59),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_142),
.B(n_53),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_228),
.B(n_244),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_100),
.C(n_96),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_229),
.B(n_196),
.Y(n_359)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_55),
.B1(n_59),
.B2(n_53),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_231),
.Y(n_344)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_165),
.A2(n_53),
.B1(n_72),
.B2(n_79),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_233),
.A2(n_237),
.B1(n_292),
.B2(n_299),
.Y(n_328)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_234),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_165),
.A2(n_77),
.B1(n_76),
.B2(n_71),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_199),
.A2(n_97),
.B1(n_78),
.B2(n_66),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_239),
.A2(n_256),
.B1(n_286),
.B2(n_300),
.Y(n_361)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_241),
.B(n_262),
.Y(n_336)
);

BUFx2_ASAP7_75t_SL g243 ( 
.A(n_171),
.Y(n_243)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_130),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_246),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_65),
.B1(n_115),
.B2(n_127),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_247),
.A2(n_286),
.B1(n_300),
.B2(n_301),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_119),
.B(n_22),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_251),
.A2(n_259),
.B(n_265),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_195),
.A2(n_121),
.B1(n_120),
.B2(n_117),
.Y(n_252)
);

AOI22x1_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_224),
.B1(n_216),
.B2(n_222),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_57),
.B(n_10),
.C(n_11),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_253),
.A2(n_260),
.B(n_295),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_254),
.A2(n_164),
.B1(n_219),
.B2(n_203),
.Y(n_343)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_143),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_256)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_258),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_215),
.A2(n_154),
.B1(n_148),
.B2(n_186),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_167),
.A2(n_6),
.B(n_15),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_201),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_217),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_153),
.Y(n_266)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_217),
.A2(n_5),
.B1(n_14),
.B2(n_13),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_268),
.A2(n_185),
.B(n_221),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_137),
.B(n_0),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_271),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_141),
.B(n_0),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_272),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_273),
.B(n_282),
.Y(n_309)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_274),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_275),
.Y(n_360)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_147),
.B(n_158),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_278),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_182),
.Y(n_279)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_184),
.Y(n_281)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_4),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_285),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_132),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_134),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_288),
.Y(n_331)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_146),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_289),
.Y(n_313)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_187),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_291),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_173),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_144),
.A2(n_5),
.B1(n_12),
.B2(n_11),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_297),
.Y(n_321)
);

INVx3_ASAP7_75t_SL g294 ( 
.A(n_181),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_294),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_135),
.A2(n_3),
.B(n_5),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_182),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_209),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_0),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g348 ( 
.A1(n_298),
.A2(n_304),
.B(n_305),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_144),
.A2(n_3),
.B1(n_12),
.B2(n_19),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_209),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_163),
.A2(n_2),
.B1(n_3),
.B2(n_194),
.Y(n_301)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_302),
.Y(n_342)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_159),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_181),
.Y(n_335)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_160),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_180),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_311),
.A2(n_334),
.B1(n_361),
.B2(n_229),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_254),
.A2(n_220),
.B1(n_194),
.B2(n_163),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_322),
.A2(n_329),
.B1(n_343),
.B2(n_239),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_170),
.B1(n_166),
.B2(n_133),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_261),
.B(n_223),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_330),
.B(n_341),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_250),
.A2(n_159),
.B1(n_164),
.B2(n_203),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_347),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_228),
.B(n_204),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_262),
.B(n_238),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_244),
.B(n_220),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_271),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_235),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_230),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_253),
.A2(n_180),
.B(n_166),
.C(n_170),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_247),
.B(n_298),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_298),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_259),
.A2(n_196),
.B1(n_219),
.B2(n_133),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_362),
.A2(n_294),
.B1(n_246),
.B2(n_263),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

AO21x2_ASAP7_75t_L g367 ( 
.A1(n_340),
.A2(n_251),
.B(n_302),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_367),
.A2(n_372),
.B1(n_388),
.B2(n_404),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_316),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_270),
.B1(n_249),
.B2(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_280),
.B1(n_272),
.B2(n_257),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_374),
.A2(n_375),
.B1(n_378),
.B2(n_409),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_272),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_385),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_377),
.A2(n_393),
.B1(n_394),
.B2(n_398),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_342),
.A2(n_269),
.B1(n_271),
.B2(n_265),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_402),
.Y(n_420)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

BUFx4f_ASAP7_75t_SL g384 ( 
.A(n_307),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_278),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_278),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_386),
.B(n_390),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_336),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_392),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_288),
.B1(n_297),
.B2(n_266),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_338),
.B(n_267),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_SL g438 ( 
.A(n_396),
.B(n_400),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_341),
.A2(n_268),
.B1(n_234),
.B2(n_242),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_399),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_281),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_401),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_287),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_330),
.B(n_285),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_403),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_322),
.A2(n_240),
.B1(n_232),
.B2(n_226),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_405),
.Y(n_421)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_406),
.A2(n_408),
.B(n_320),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_245),
.C(n_255),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_410),
.C(n_248),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_336),
.B(n_242),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_339),
.A2(n_284),
.B1(n_277),
.B2(n_276),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_339),
.B(n_248),
.C(n_263),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_411),
.A2(n_311),
.B1(n_318),
.B2(n_360),
.Y(n_423)
);

AO22x1_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_356),
.B1(n_344),
.B2(n_358),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_369),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_423),
.A2(n_409),
.B1(n_401),
.B2(n_394),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_405),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_311),
.B1(n_344),
.B2(n_328),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_406),
.B1(n_393),
.B2(n_384),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_317),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_320),
.C(n_325),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_447),
.C(n_407),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_367),
.A2(n_358),
.B1(n_315),
.B2(n_329),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_430),
.A2(n_431),
.B1(n_436),
.B2(n_439),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_367),
.A2(n_315),
.B1(n_318),
.B2(n_337),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_367),
.A2(n_312),
.B1(n_321),
.B2(n_313),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_375),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_437),
.A2(n_446),
.B1(n_404),
.B2(n_386),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_372),
.A2(n_354),
.B1(n_325),
.B2(n_323),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_371),
.A2(n_323),
.B1(n_352),
.B2(n_303),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_440),
.A2(n_389),
.B1(n_391),
.B2(n_373),
.Y(n_466)
);

A2O1A1O1Ixp25_ASAP7_75t_L g443 ( 
.A1(n_376),
.A2(n_323),
.B(n_310),
.C(n_309),
.D(n_319),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_443),
.A2(n_396),
.B(n_385),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_375),
.A2(n_319),
.B1(n_352),
.B2(n_324),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_380),
.B(n_236),
.C(n_274),
.Y(n_447)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_397),
.C(n_402),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_447),
.C(n_444),
.Y(n_513)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_453),
.A2(n_454),
.B(n_456),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_413),
.A2(n_400),
.B(n_390),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_437),
.A2(n_436),
.B(n_446),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_395),
.B(n_410),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_457),
.A2(n_467),
.B(n_481),
.Y(n_486)
);

OAI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_429),
.A2(n_388),
.B1(n_403),
.B2(n_395),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_459),
.A2(n_465),
.B1(n_473),
.B2(n_480),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_460),
.A2(n_412),
.B1(n_443),
.B2(n_445),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_461),
.B(n_483),
.Y(n_503)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_463),
.A2(n_412),
.B1(n_439),
.B2(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_429),
.A2(n_381),
.B1(n_378),
.B2(n_365),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_425),
.A2(n_379),
.B1(n_366),
.B2(n_392),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_420),
.B(n_353),
.C(n_305),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_472),
.C(n_427),
.Y(n_504)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_442),
.A2(n_368),
.B1(n_382),
.B2(n_383),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_425),
.A2(n_413),
.B1(n_431),
.B2(n_419),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_474),
.A2(n_475),
.B1(n_477),
.B2(n_478),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_419),
.A2(n_384),
.B1(n_353),
.B2(n_350),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_422),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_484),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_440),
.A2(n_294),
.B1(n_346),
.B2(n_290),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_426),
.A2(n_346),
.B1(n_363),
.B2(n_316),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_449),
.A2(n_307),
.B(n_363),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_416),
.B(n_424),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_417),
.A2(n_421),
.B1(n_445),
.B2(n_449),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_443),
.A2(n_326),
.B(n_317),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_482),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_326),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_416),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_487),
.A2(n_497),
.B1(n_513),
.B2(n_514),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_480),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_490),
.B(n_496),
.Y(n_544)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_491),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_479),
.Y(n_496)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_506),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_415),
.Y(n_505)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_433),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_475),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_507),
.Y(n_522)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_457),
.B(n_433),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_470),
.C(n_453),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_472),
.B(n_428),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_483),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_474),
.A2(n_418),
.B1(n_415),
.B2(n_438),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_516),
.B1(n_458),
.B2(n_459),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_418),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_451),
.C(n_471),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_456),
.A2(n_430),
.B1(n_423),
.B2(n_448),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_463),
.A2(n_448),
.B1(n_434),
.B2(n_444),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_515),
.A2(n_466),
.B1(n_478),
.B2(n_482),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_458),
.A2(n_468),
.B1(n_467),
.B2(n_460),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_521),
.A2(n_531),
.B1(n_539),
.B2(n_489),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_517),
.A2(n_481),
.B(n_488),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_524),
.A2(n_486),
.B(n_496),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_525),
.B(n_534),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_532),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_528),
.A2(n_535),
.B1(n_520),
.B2(n_522),
.Y(n_563)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_529),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_454),
.C(n_473),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_540),
.C(n_543),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_454),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_505),
.B(n_441),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_533),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_469),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_489),
.A2(n_477),
.B1(n_464),
.B2(n_462),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_535),
.A2(n_498),
.B1(n_507),
.B2(n_490),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_511),
.B(n_441),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_538),
.Y(n_552)
);

FAx1_ASAP7_75t_SL g538 ( 
.A(n_509),
.B(n_435),
.CI(n_450),
.CON(n_538),
.SN(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_516),
.A2(n_452),
.B1(n_435),
.B2(n_316),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_504),
.B(n_296),
.C(n_357),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_500),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_541),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_357),
.C(n_293),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_497),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_545),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_554),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_549),
.A2(n_551),
.B1(n_558),
.B2(n_566),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_521),
.A2(n_487),
.B1(n_514),
.B2(n_515),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_486),
.C(n_517),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_561),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g556 ( 
.A(n_530),
.B(n_508),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_556),
.B(n_499),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_520),
.A2(n_502),
.B1(n_501),
.B2(n_499),
.Y(n_558)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_523),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_523),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_562),
.B(n_564),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_565),
.Y(n_572)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_542),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_544),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_566),
.A2(n_528),
.B1(n_538),
.B2(n_518),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_501),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_550),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_568),
.B(n_583),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_540),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_571),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_525),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_548),
.B(n_534),
.C(n_543),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_527),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_576),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_532),
.C(n_519),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_577),
.C(n_579),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_536),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_556),
.B(n_544),
.C(n_524),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_518),
.C(n_539),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_580),
.A2(n_585),
.B1(n_563),
.B2(n_557),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_559),
.A2(n_538),
.B(n_485),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_581),
.A2(n_562),
.B(n_564),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_554),
.B(n_493),
.C(n_485),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_547),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_577),
.A2(n_559),
.B1(n_551),
.B2(n_557),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_587),
.A2(n_593),
.B1(n_495),
.B2(n_494),
.Y(n_611)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_584),
.Y(n_588)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_588),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_590),
.B(n_595),
.Y(n_601)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_582),
.Y(n_591)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_570),
.Y(n_592)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_572),
.A2(n_546),
.B1(n_565),
.B2(n_552),
.Y(n_593)
);

BUFx24_ASAP7_75t_SL g596 ( 
.A(n_578),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_579),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_585),
.A2(n_546),
.B1(n_555),
.B2(n_561),
.Y(n_597)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_597),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_598),
.A2(n_572),
.B(n_580),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_602),
.A2(n_604),
.B(n_607),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_573),
.C(n_575),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_603),
.B(n_608),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_599),
.A2(n_578),
.B(n_558),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_583),
.C(n_493),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_594),
.B(n_495),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_611),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_612),
.A2(n_593),
.B1(n_597),
.B2(n_590),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_613),
.B(n_614),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_595),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_608),
.B(n_586),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_617),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_601),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_619),
.B(n_620),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_594),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_605),
.B(n_589),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_621),
.B(n_306),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_619),
.A2(n_610),
.B1(n_601),
.B2(n_609),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_623),
.B(n_625),
.Y(n_630)
);

A2O1A1O1Ixp25_ASAP7_75t_L g625 ( 
.A1(n_616),
.A2(n_589),
.B(n_494),
.C(n_306),
.D(n_283),
.Y(n_625)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_627),
.Y(n_628)
);

NOR2x1_ASAP7_75t_R g629 ( 
.A(n_624),
.B(n_615),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_629),
.B(n_622),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_631),
.A2(n_632),
.B1(n_628),
.B2(n_279),
.Y(n_633)
);

AOI31xp33_ASAP7_75t_L g632 ( 
.A1(n_630),
.A2(n_618),
.A3(n_626),
.B(n_617),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_275),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_634),
.A2(n_258),
.B(n_351),
.Y(n_635)
);

XNOR2x2_ASAP7_75t_SL g636 ( 
.A(n_635),
.B(n_351),
.Y(n_636)
);


endmodule