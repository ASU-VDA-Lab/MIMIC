module fake_netlist_5_1739_n_760 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_760);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_760;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_685;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_35),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_24),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_8),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_31),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_69),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_48),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_30),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_106),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_39),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_36),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_71),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_51),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_14),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_85),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_41),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_73),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_40),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_34),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_0),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_18),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_0),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_1),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_1),
.B(n_2),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_3),
.B(n_4),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_20),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_153),
.Y(n_228)
);

CKINVDCx6p67_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_148),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_152),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_213),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_190),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_R g253 ( 
.A(n_212),
.B(n_150),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_210),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

BUFx16f_ASAP7_75t_R g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_204),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_214),
.B(n_150),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_204),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_R g271 ( 
.A(n_203),
.B(n_147),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_217),
.A2(n_220),
.B(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_226),
.B(n_162),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_234),
.B(n_193),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_226),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_157),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_205),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_239),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

NOR2x1p5_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_261),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_226),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_248),
.B(n_206),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_206),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_205),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_255),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_205),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_205),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_242),
.B(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_239),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_232),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_232),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_250),
.B(n_205),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_262),
.B(n_238),
.C(n_223),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_267),
.B(n_185),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_232),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_230),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_209),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_230),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_237),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_271),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_253),
.B(n_237),
.C(n_184),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_259),
.B(n_237),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_264),
.B(n_271),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_246),
.B(n_237),
.Y(n_339)
);

OR2x6_ASAP7_75t_L g340 ( 
.A(n_240),
.B(n_225),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_247),
.B(n_237),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_241),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_277),
.A2(n_225),
.B(n_216),
.C(n_220),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_244),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_245),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_282),
.B(n_187),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_256),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_244),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_322),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_345),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_289),
.B(n_221),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_349),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_179),
.B1(n_163),
.B2(n_164),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_216),
.B1(n_198),
.B2(n_221),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_348),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_178),
.B1(n_166),
.B2(n_167),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_221),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_159),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_6),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_338),
.A2(n_168),
.B1(n_173),
.B2(n_176),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_288),
.A2(n_196),
.B1(n_195),
.B2(n_186),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_293),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_342),
.Y(n_374)
);

OR2x6_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_200),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_307),
.B(n_182),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_336),
.B(n_200),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_207),
.B1(n_200),
.B2(n_80),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_319),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_207),
.B1(n_9),
.B2(n_10),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_331),
.A2(n_207),
.B1(n_79),
.B2(n_81),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_315),
.B(n_316),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_336),
.B(n_207),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_327),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_347),
.A2(n_207),
.B1(n_9),
.B2(n_12),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_339),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_21),
.Y(n_394)
);

BUFx4f_ASAP7_75t_SL g395 ( 
.A(n_321),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_299),
.B(n_7),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_316),
.B(n_22),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_299),
.A2(n_86),
.B1(n_143),
.B2(n_142),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_301),
.B(n_23),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_301),
.B(n_25),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_301),
.B(n_27),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_301),
.B(n_29),
.Y(n_403)
);

OR2x2_ASAP7_75t_SL g404 ( 
.A(n_341),
.B(n_12),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_313),
.Y(n_405)
);

OAI21xp33_ASAP7_75t_L g406 ( 
.A1(n_321),
.A2(n_13),
.B(n_14),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_301),
.B(n_32),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_343),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_335),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_311),
.B(n_15),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

NOR2x2_ASAP7_75t_L g416 ( 
.A(n_340),
.B(n_16),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_340),
.A2(n_17),
.B1(n_33),
.B2(n_37),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_354),
.B(n_320),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_310),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_318),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_SL g423 ( 
.A(n_357),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_363),
.A2(n_415),
.B(n_355),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_371),
.B(n_393),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_295),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_356),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_292),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_352),
.B(n_301),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_314),
.B(n_333),
.C(n_317),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_330),
.B(n_334),
.C(n_329),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

BUFx4f_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_414),
.A2(n_309),
.B(n_306),
.C(n_350),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_355),
.A2(n_350),
.B(n_344),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_371),
.A2(n_350),
.B(n_344),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_353),
.B(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_344),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_350),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_38),
.Y(n_442)
);

BUFx8_ASAP7_75t_L g443 ( 
.A(n_396),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_42),
.B(n_43),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_397),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_361),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_351),
.A2(n_47),
.B(n_49),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_359),
.A2(n_50),
.B(n_52),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_377),
.B(n_53),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_366),
.A2(n_57),
.B(n_58),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_395),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_366),
.A2(n_59),
.B(n_60),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_362),
.B(n_62),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_387),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_358),
.B(n_63),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_392),
.B(n_64),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_368),
.B(n_66),
.Y(n_469)
);

OAI22x1_ASAP7_75t_L g470 ( 
.A1(n_412),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_368),
.B(n_72),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_417),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_472)
);

NAND2x1_ASAP7_75t_L g473 ( 
.A(n_373),
.B(n_77),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_398),
.A2(n_82),
.B1(n_87),
.B2(n_89),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_420),
.A2(n_384),
.B(n_378),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_438),
.A2(n_407),
.B(n_403),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_432),
.A2(n_407),
.B(n_403),
.Y(n_479)
);

BUFx12f_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

BUFx2_ASAP7_75t_R g481 ( 
.A(n_446),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_443),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_428),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_450),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_449),
.A2(n_431),
.B(n_426),
.Y(n_487)
);

BUFx2_ASAP7_75t_R g488 ( 
.A(n_457),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_425),
.A2(n_402),
.B(n_401),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_367),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_437),
.A2(n_402),
.B(n_401),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_441),
.A2(n_400),
.B(n_399),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_453),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_464),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_400),
.B(n_382),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_379),
.B(n_381),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_375),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_427),
.Y(n_502)
);

BUFx4f_ASAP7_75t_SL g503 ( 
.A(n_459),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_SL g504 ( 
.A(n_465),
.B(n_373),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_444),
.A2(n_391),
.B(n_375),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_422),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_418),
.B(n_375),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_448),
.A2(n_90),
.B(n_91),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_434),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_466),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_93),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_442),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_469),
.A2(n_96),
.B(n_97),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_424),
.B(n_98),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_451),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_454),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_454),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_481),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g522 ( 
.A1(n_491),
.A2(n_472),
.B(n_471),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_489),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_463),
.B1(n_507),
.B2(n_460),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_495),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_495),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_517),
.A2(n_470),
.B1(n_452),
.B2(n_461),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_423),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_515),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_462),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_477),
.A2(n_473),
.B(n_440),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_490),
.A2(n_430),
.B(n_468),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_506),
.A2(n_429),
.B1(n_455),
.B2(n_474),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_496),
.Y(n_537)
);

BUFx4f_ASAP7_75t_SL g538 ( 
.A(n_480),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_515),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_429),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_445),
.B(n_458),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_483),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_475),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

AO21x1_ASAP7_75t_SL g548 ( 
.A1(n_500),
.A2(n_456),
.B(n_102),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_513),
.A2(n_501),
.B1(n_517),
.B2(n_476),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_498),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_486),
.B(n_101),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_494),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_498),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_492),
.A2(n_108),
.B(n_109),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_R g560 ( 
.A1(n_510),
.A2(n_110),
.B1(n_112),
.B2(n_114),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_494),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_561)
);

BUFx2_ASAP7_75t_R g562 ( 
.A(n_502),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_525),
.Y(n_563)
);

AND4x1_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_488),
.C(n_503),
.D(n_480),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_521),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_509),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_521),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_527),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_538),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_542),
.B(n_494),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_484),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_537),
.B(n_484),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_533),
.B(n_503),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_520),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_562),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_R g577 ( 
.A(n_554),
.B(n_505),
.Y(n_577)
);

BUFx4f_ASAP7_75t_SL g578 ( 
.A(n_552),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_524),
.B(n_529),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_R g580 ( 
.A(n_554),
.B(n_482),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_532),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_553),
.Y(n_583)
);

O2A1O1Ixp33_ASAP7_75t_SL g584 ( 
.A1(n_522),
.A2(n_512),
.B(n_516),
.C(n_505),
.Y(n_584)
);

AND2x4_ASAP7_75t_SL g585 ( 
.A(n_554),
.B(n_519),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_528),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_540),
.B(n_482),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

NOR3xp33_ASAP7_75t_SL g589 ( 
.A(n_549),
.B(n_478),
.C(n_520),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_R g591 ( 
.A(n_540),
.B(n_478),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_539),
.B(n_520),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_SL g593 ( 
.A(n_536),
.B(n_545),
.C(n_547),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_560),
.A2(n_548),
.B1(n_530),
.B2(n_543),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_540),
.B(n_511),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_556),
.A2(n_512),
.B1(n_519),
.B2(n_511),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_540),
.B(n_511),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_523),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_516),
.B1(n_511),
.B2(n_498),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_531),
.B(n_493),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_532),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_SL g605 ( 
.A(n_531),
.B(n_497),
.C(n_493),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_SL g607 ( 
.A1(n_551),
.A2(n_497),
.B(n_479),
.C(n_120),
.Y(n_607)
);

NOR2x1_ASAP7_75t_SL g608 ( 
.A(n_548),
.B(n_479),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_568),
.B(n_557),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_541),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_546),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_586),
.Y(n_613)
);

AOI21xp33_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_550),
.B(n_534),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_604),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_535),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_575),
.B(n_551),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_602),
.Y(n_619)
);

NAND2x1p5_ASAP7_75t_L g620 ( 
.A(n_601),
.B(n_559),
.Y(n_620)
);

OAI211xp5_ASAP7_75t_L g621 ( 
.A1(n_593),
.A2(n_535),
.B(n_559),
.C(n_523),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_579),
.B(n_534),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_594),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_590),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_608),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_583),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_605),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_589),
.B(n_492),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_145),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_592),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_594),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_607),
.A2(n_118),
.B(n_119),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_599),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_594),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_600),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_600),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_124),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_584),
.Y(n_641)
);

OAI211xp5_ASAP7_75t_SL g642 ( 
.A1(n_566),
.A2(n_125),
.B(n_127),
.C(n_128),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_627),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_581),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_612),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_612),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_615),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_628),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_611),
.B(n_578),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_625),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_634),
.B(n_564),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_638),
.B(n_565),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_610),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_629),
.B(n_574),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_625),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_623),
.B(n_603),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_619),
.B(n_597),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_642),
.A2(n_621),
.B(n_614),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_631),
.B(n_587),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_635),
.B(n_567),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_616),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_635),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_616),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_623),
.B(n_565),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_632),
.B(n_576),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_609),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_651),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_648),
.B(n_619),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_650),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_650),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_647),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_664),
.B(n_641),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_658),
.B(n_617),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_654),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_655),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_662),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_643),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_645),
.B(n_646),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_645),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_646),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_669),
.B(n_641),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_669),
.B(n_617),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_676),
.A2(n_652),
.B1(n_656),
.B2(n_667),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_672),
.Y(n_687)
);

OAI211xp5_ASAP7_75t_SL g688 ( 
.A1(n_675),
.A2(n_649),
.B(n_657),
.C(n_665),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_673),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_680),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_674),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_683),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_682),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_677),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_678),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_684),
.B(n_656),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_692),
.Y(n_697)
);

AOI21xp33_ASAP7_75t_L g698 ( 
.A1(n_688),
.A2(n_652),
.B(n_675),
.Y(n_698)
);

XOR2x2_ASAP7_75t_L g699 ( 
.A(n_686),
.B(n_661),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_644),
.B(n_660),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_696),
.A2(n_630),
.B(n_684),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_697),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_690),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_700),
.A2(n_653),
.B(n_668),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_699),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_698),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_706),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.C(n_702),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_705),
.B(n_690),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_705),
.B(n_569),
.Y(n_709)
);

AOI221xp5_ASAP7_75t_L g710 ( 
.A1(n_706),
.A2(n_644),
.B1(n_691),
.B2(n_694),
.C(n_687),
.Y(n_710)
);

NOR2x1_ASAP7_75t_L g711 ( 
.A(n_708),
.B(n_671),
.Y(n_711)
);

OAI21xp33_ASAP7_75t_SL g712 ( 
.A1(n_707),
.A2(n_710),
.B(n_709),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_667),
.B(n_670),
.Y(n_713)
);

NOR2x1_ASAP7_75t_L g714 ( 
.A(n_713),
.B(n_631),
.Y(n_714)
);

XNOR2xp5_ASAP7_75t_L g715 ( 
.A(n_711),
.B(n_653),
.Y(n_715)
);

AOI221x1_ASAP7_75t_L g716 ( 
.A1(n_712),
.A2(n_689),
.B1(n_633),
.B2(n_639),
.C(n_679),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_SL g717 ( 
.A(n_712),
.B(n_618),
.C(n_663),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_714),
.B(n_658),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_716),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_659),
.B1(n_685),
.B2(n_695),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_659),
.B1(n_685),
.B2(n_630),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_715),
.Y(n_723)
);

NOR2x1_ASAP7_75t_L g724 ( 
.A(n_715),
.B(n_591),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_693),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_719),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_720),
.B(n_681),
.Y(n_728)
);

NAND5xp2_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_721),
.C(n_640),
.D(n_620),
.E(n_580),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_723),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_720),
.B(n_681),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_720),
.B(n_636),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_727),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_726),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_725),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_732),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_730),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_728),
.A2(n_640),
.B(n_634),
.Y(n_738)
);

NOR2x1p5_ASAP7_75t_L g739 ( 
.A(n_731),
.B(n_637),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_729),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_SL g741 ( 
.A1(n_735),
.A2(n_630),
.B(n_585),
.Y(n_741)
);

OAI22x1_ASAP7_75t_SL g742 ( 
.A1(n_736),
.A2(n_636),
.B1(n_637),
.B2(n_598),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_733),
.B(n_637),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_734),
.Y(n_745)
);

XNOR2x1_ASAP7_75t_L g746 ( 
.A(n_737),
.B(n_129),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_739),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_740),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_743),
.B(n_738),
.Y(n_749)
);

OAI31xp33_ASAP7_75t_L g750 ( 
.A1(n_744),
.A2(n_620),
.A3(n_596),
.B(n_626),
.Y(n_750)
);

OAI22x1_ASAP7_75t_L g751 ( 
.A1(n_747),
.A2(n_746),
.B1(n_742),
.B2(n_741),
.Y(n_751)
);

XOR2xp5_ASAP7_75t_L g752 ( 
.A(n_751),
.B(n_132),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_749),
.B(n_626),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_753),
.Y(n_755)
);

AO22x2_ASAP7_75t_L g756 ( 
.A1(n_752),
.A2(n_750),
.B1(n_622),
.B2(n_613),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_755),
.B(n_754),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_756),
.B1(n_624),
.B2(n_634),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_758),
.B(n_624),
.Y(n_759)
);

AOI211xp5_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_133),
.B(n_134),
.C(n_135),
.Y(n_760)
);


endmodule