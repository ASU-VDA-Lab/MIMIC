module real_jpeg_1624_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_59),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_59),
.B1(n_65),
.B2(n_67),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_2),
.A2(n_56),
.B1(n_65),
.B2(n_67),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_27),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_44),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_36),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_62),
.C(n_65),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_3),
.B(n_80),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_71),
.Y(n_173)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_65),
.B1(n_67),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_8),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_8),
.A2(n_40),
.B1(n_65),
.B2(n_67),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_11),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_12),
.A2(n_65),
.B1(n_67),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_15),
.A2(n_65),
.B1(n_67),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_117),
.B1(n_191),
.B2(n_192),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_19),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_96),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_87),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_22),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_23),
.B(n_42),
.C(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_24),
.A2(n_33),
.B1(n_39),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_28),
.A2(n_31),
.A3(n_36),
.B1(n_38),
.B2(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_30),
.B(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_34),
.B(n_128),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_36),
.A2(n_46),
.A3(n_48),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_41)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_52),
.B1(n_54),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_43),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_43),
.A2(n_54),
.B1(n_89),
.B2(n_150),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

AO22x2_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_45),
.B(n_50),
.Y(n_129)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_46),
.B(n_159),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_68),
.B2(n_71),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_60),
.B1(n_71),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_60),
.A2(n_71),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_60),
.A2(n_71),
.B1(n_141),
.B2(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_69),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_64),
.A2(n_113),
.B1(n_124),
.B2(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_65),
.B(n_169),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_87),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_80),
.B1(n_132),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_78),
.A2(n_80),
.B1(n_128),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_78),
.A2(n_80),
.B1(n_171),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_85),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_109),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_79),
.A2(n_109),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.C(n_93),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_136),
.B(n_190),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_134),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_134),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_120),
.B(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_125),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_185),
.B(n_189),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_154),
.B(n_184),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_146),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_143),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.C(n_152),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_165),
.B(n_183),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_177),
.B(n_182),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_172),
.B(n_176),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_188),
.Y(n_189)
);


endmodule