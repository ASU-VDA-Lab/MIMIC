module fake_jpeg_3571_n_689 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_689);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_689;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_61),
.Y(n_169)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_71),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_9),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_77),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_0),
.CON(n_73),
.SN(n_73)
);

HAxp5_ASAP7_75t_SL g199 ( 
.A(n_73),
.B(n_15),
.CON(n_199),
.SN(n_199)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_9),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_80),
.Y(n_219)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_40),
.B(n_8),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_82),
.B(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_20),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g172 ( 
.A(n_84),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_30),
.A2(n_10),
.B(n_18),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_89),
.B(n_99),
.Y(n_166)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_90),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_42),
.A2(n_7),
.B1(n_18),
.B2(n_17),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_101),
.Y(n_211)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_105),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g183 ( 
.A(n_110),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_31),
.Y(n_111)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_7),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_129),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_45),
.B(n_19),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_132),
.Y(n_148)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_31),
.Y(n_125)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_27),
.Y(n_128)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_57),
.B(n_7),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_27),
.Y(n_130)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_45),
.B(n_11),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_75),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_155),
.B(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_158),
.A2(n_198),
.B(n_201),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_73),
.B(n_32),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_108),
.A2(n_31),
.B1(n_58),
.B2(n_27),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_177),
.A2(n_198),
.B1(n_217),
.B2(n_37),
.Y(n_248)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_84),
.B(n_42),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_180),
.B(n_197),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_91),
.B(n_25),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_128),
.A2(n_58),
.B1(n_39),
.B2(n_48),
.Y(n_198)
);

NAND2x1_ASAP7_75t_L g284 ( 
.A(n_199),
.B(n_11),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_91),
.B(n_25),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_218),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_87),
.A2(n_58),
.B1(n_39),
.B2(n_49),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_201),
.A2(n_206),
.B1(n_208),
.B2(n_212),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_88),
.A2(n_39),
.B1(n_53),
.B2(n_43),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_130),
.A2(n_37),
.B1(n_43),
.B2(n_53),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_117),
.A2(n_37),
.B1(n_52),
.B2(n_32),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_118),
.A2(n_52),
.B1(n_33),
.B2(n_23),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_127),
.B(n_23),
.Y(n_218)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_67),
.Y(n_224)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_68),
.B(n_37),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_0),
.Y(n_301)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_90),
.Y(n_226)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_80),
.B(n_33),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_148),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_133),
.B(n_37),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_229),
.B(n_257),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_233),
.Y(n_338)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_235),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_241),
.Y(n_357)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_150),
.Y(n_242)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_243),
.B(n_255),
.Y(n_356)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_245),
.A2(n_259),
.B1(n_296),
.B2(n_304),
.Y(n_345)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_248),
.B(n_295),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_142),
.A2(n_92),
.B1(n_106),
.B2(n_104),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_165),
.A2(n_96),
.B1(n_103),
.B2(n_100),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_163),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_137),
.B(n_95),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_166),
.A2(n_28),
.B1(n_26),
.B2(n_98),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_173),
.B(n_14),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_261),
.B(n_263),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_262),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_173),
.B(n_14),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_271),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_155),
.B(n_112),
.C(n_28),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_225),
.C(n_216),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_135),
.B(n_28),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_267),
.Y(n_336)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_157),
.Y(n_269)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_168),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_272),
.B(n_274),
.Y(n_337)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_170),
.Y(n_273)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_273),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_141),
.B(n_166),
.Y(n_274)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_160),
.A2(n_56),
.A3(n_11),
.B1(n_15),
.B2(n_19),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_280),
.A2(n_154),
.B(n_219),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_141),
.B(n_11),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_282),
.B(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_283),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_292),
.Y(n_348)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

INVx4_ASAP7_75t_SL g286 ( 
.A(n_172),
.Y(n_286)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_286),
.Y(n_364)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_288),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_289),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_191),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_160),
.B(n_6),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_293),
.Y(n_320)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_149),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_138),
.A2(n_56),
.B1(n_6),
.B2(n_15),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_145),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_297),
.B(n_298),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_161),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_139),
.B(n_19),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_185),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_300),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_305),
.Y(n_319)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_302),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_212),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_307),
.B1(n_216),
.B2(n_162),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_140),
.A2(n_56),
.B1(n_18),
.B2(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_136),
.B(n_17),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g307 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_162),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_190),
.B(n_0),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_1),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_194),
.B(n_214),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_208),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_241),
.A2(n_275),
.B(n_271),
.C(n_288),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_315),
.A2(n_307),
.B(n_284),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_328),
.B(n_329),
.C(n_346),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_246),
.B(n_236),
.C(n_266),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_SL g407 ( 
.A1(n_331),
.A2(n_293),
.B(n_297),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_248),
.A2(n_205),
.B1(n_209),
.B2(n_204),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_353),
.B1(n_369),
.B2(n_252),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_339),
.B(n_372),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_246),
.B(n_202),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_352),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_259),
.A2(n_188),
.B1(n_187),
.B2(n_189),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_370),
.B1(n_289),
.B2(n_262),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_254),
.B(n_199),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_231),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_192),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_275),
.A2(n_196),
.B1(n_184),
.B2(n_171),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_280),
.B(n_167),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_291),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_267),
.B(n_240),
.C(n_237),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_328),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_303),
.A2(n_176),
.B1(n_196),
.B2(n_184),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_275),
.A2(n_221),
.B1(n_154),
.B2(n_219),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_373),
.B(n_394),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_286),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_384),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_376),
.A2(n_386),
.B1(n_407),
.B2(n_343),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_267),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_377),
.B(n_322),
.C(n_317),
.Y(n_442)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_315),
.A2(n_250),
.B(n_230),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_381),
.B(n_400),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_380),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_341),
.A2(n_357),
.B(n_336),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_382),
.A2(n_412),
.B1(n_421),
.B2(n_314),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_383),
.B(n_406),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_230),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_370),
.A2(n_268),
.B1(n_281),
.B2(n_251),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_385),
.A2(n_391),
.B1(n_420),
.B2(n_376),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_350),
.A2(n_363),
.B1(n_344),
.B2(n_345),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_387),
.B(n_389),
.Y(n_437)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_388),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_330),
.B(n_235),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_393),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_232),
.B1(n_234),
.B2(n_221),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_233),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_285),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_372),
.B(n_294),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_401),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_313),
.A2(n_276),
.B(n_253),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_398),
.A2(n_369),
.B(n_366),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_359),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_405),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_348),
.A2(n_304),
.B(n_296),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_321),
.B(n_308),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_356),
.B(n_249),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_408),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_427)
);

INVx13_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_410),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_359),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_311),
.B(n_365),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_319),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_339),
.B(n_249),
.Y(n_414)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_320),
.B(n_273),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_239),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_418),
.A2(n_419),
.B1(n_231),
.B2(n_334),
.Y(n_449)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_342),
.A2(n_302),
.B1(n_269),
.B2(n_222),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_359),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_422),
.A2(n_431),
.B(n_434),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_442),
.C(n_403),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_313),
.B1(n_343),
.B2(n_331),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_428),
.A2(n_440),
.B1(n_450),
.B2(n_399),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_401),
.A2(n_408),
.B1(n_373),
.B2(n_374),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_430),
.A2(n_432),
.B1(n_433),
.B2(n_435),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_408),
.A2(n_333),
.B1(n_348),
.B2(n_358),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_374),
.A2(n_319),
.B1(n_352),
.B2(n_366),
.Y(n_433)
);

O2A1O1Ixp33_ASAP7_75t_SL g434 ( 
.A1(n_379),
.A2(n_362),
.B(n_347),
.C(n_312),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_397),
.A2(n_258),
.B1(n_371),
.B2(n_354),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_397),
.A2(n_371),
.B1(n_354),
.B2(n_318),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_436),
.A2(n_441),
.B1(n_444),
.B2(n_451),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_382),
.A2(n_346),
.B1(n_318),
.B2(n_355),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_381),
.A2(n_322),
.B1(n_317),
.B2(n_355),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_385),
.A2(n_314),
.B1(n_323),
.B2(n_312),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_446),
.A2(n_449),
.B(n_398),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_349),
.B1(n_323),
.B2(n_361),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_414),
.A2(n_335),
.B1(n_327),
.B2(n_361),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_414),
.A2(n_335),
.B1(n_327),
.B2(n_153),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_457),
.A2(n_340),
.B1(n_388),
.B2(n_338),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_383),
.B(n_368),
.C(n_298),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_403),
.C(n_394),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_437),
.B(n_384),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_463),
.B(n_471),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_483),
.B1(n_485),
.B2(n_441),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_396),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_467),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_454),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_377),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_480),
.C(n_492),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_406),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_473),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_454),
.B(n_413),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_430),
.A2(n_375),
.B1(n_412),
.B2(n_421),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_472),
.A2(n_479),
.B1(n_481),
.B2(n_486),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_416),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_455),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g531 ( 
.A(n_475),
.Y(n_531)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_476),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_433),
.B(n_393),
.Y(n_477)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_435),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_422),
.A2(n_446),
.B1(n_428),
.B2(n_456),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_432),
.A2(n_400),
.B1(n_394),
.B2(n_390),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_482),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_456),
.A2(n_394),
.B1(n_420),
.B2(n_391),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_456),
.A2(n_415),
.B1(n_417),
.B2(n_419),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_431),
.A2(n_460),
.B1(n_440),
.B2(n_427),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_426),
.A2(n_404),
.B(n_395),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_487),
.A2(n_493),
.B(n_452),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_444),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_488),
.B(n_494),
.Y(n_522)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_489),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_392),
.Y(n_490)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_442),
.C(n_424),
.Y(n_492)
);

OAI32xp33_ASAP7_75t_L g493 ( 
.A1(n_460),
.A2(n_378),
.A3(n_380),
.B1(n_368),
.B2(n_340),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_458),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_439),
.Y(n_495)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_495),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_450),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_496),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_388),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_497),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_462),
.A2(n_411),
.B1(n_402),
.B2(n_409),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_427),
.A2(n_411),
.B1(n_402),
.B2(n_316),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_484),
.A2(n_426),
.B1(n_462),
.B2(n_434),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_502),
.A2(n_494),
.B1(n_485),
.B2(n_483),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_473),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_514),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_461),
.C(n_424),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_513),
.C(n_515),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_511),
.A2(n_521),
.B1(n_523),
.B2(n_529),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_497),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_480),
.B(n_438),
.C(n_425),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_445),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_524),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_425),
.C(n_445),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_517),
.B(n_518),
.C(n_520),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_451),
.C(n_457),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_490),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_519),
.B(n_465),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_469),
.B(n_434),
.C(n_449),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_466),
.A2(n_429),
.B1(n_443),
.B2(n_447),
.Y(n_521)
);

AOI22x1_ASAP7_75t_L g523 ( 
.A1(n_479),
.A2(n_453),
.B1(n_447),
.B2(n_452),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_492),
.B(n_452),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_471),
.B(n_453),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_532),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_466),
.A2(n_443),
.B1(n_452),
.B2(n_316),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_530),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_472),
.B(n_410),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_410),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_537),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_481),
.B(n_409),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_484),
.B(n_423),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_468),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_475),
.Y(n_539)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_526),
.A2(n_486),
.B1(n_464),
.B2(n_467),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_540),
.A2(n_549),
.B1(n_553),
.B2(n_556),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_517),
.B(n_463),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_557),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_487),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_544),
.B(n_567),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_528),
.Y(n_545)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_537),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_512),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_522),
.Y(n_550)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_550),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_560),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_511),
.A2(n_496),
.B1(n_488),
.B2(n_491),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_554),
.A2(n_570),
.B1(n_532),
.B2(n_520),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_527),
.B(n_493),
.Y(n_555)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_555),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_504),
.Y(n_556)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_501),
.Y(n_559)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_559),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_515),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g561 ( 
.A(n_504),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_561),
.A2(n_562),
.B1(n_525),
.B2(n_498),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_534),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g564 ( 
.A(n_506),
.B(n_468),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g584 ( 
.A(n_564),
.B(n_565),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_506),
.B(n_470),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_566),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_524),
.B(n_491),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_510),
.B(n_476),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_513),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_505),
.A2(n_482),
.B1(n_499),
.B2(n_474),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_534),
.B(n_495),
.Y(n_571)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_571),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_553),
.A2(n_526),
.B1(n_530),
.B2(n_521),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_574),
.A2(n_554),
.B1(n_555),
.B2(n_568),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_578),
.B(n_590),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_535),
.Y(n_581)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_502),
.B(n_509),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_582),
.A2(n_588),
.B(n_423),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_593),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_539),
.B(n_489),
.Y(n_585)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_585),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_586),
.A2(n_589),
.B1(n_598),
.B2(n_541),
.Y(n_616)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_542),
.Y(n_587)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_540),
.A2(n_533),
.B(n_529),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_548),
.A2(n_518),
.B1(n_523),
.B2(n_500),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_523),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_536),
.Y(n_593)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_545),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_596),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_551),
.B(n_546),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_597),
.B(n_423),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_599),
.A2(n_601),
.B1(n_586),
.B2(n_589),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_577),
.A2(n_570),
.B1(n_552),
.B2(n_563),
.Y(n_601)
);

NOR2x1_ASAP7_75t_SL g602 ( 
.A(n_572),
.B(n_547),
.Y(n_602)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_602),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_546),
.C(n_560),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_604),
.B(n_605),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_567),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_565),
.Y(n_607)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_607),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_573),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_608),
.B(n_609),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_558),
.C(n_564),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_573),
.Y(n_610)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_610),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_613),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_558),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_544),
.C(n_563),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_584),
.C(n_579),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_591),
.B(n_541),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_615),
.B(n_618),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_616),
.A2(n_574),
.B1(n_576),
.B2(n_578),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_619),
.B(n_620),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g620 ( 
.A1(n_588),
.A2(n_338),
.B(n_270),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_622),
.B(n_629),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_576),
.C(n_579),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_623),
.B(n_628),
.Y(n_652)
);

NOR2x1_ASAP7_75t_SL g625 ( 
.A(n_603),
.B(n_575),
.Y(n_625)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_625),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_610),
.A2(n_582),
.B1(n_585),
.B2(n_581),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_630),
.B(n_638),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_584),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_634),
.B(n_606),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_612),
.B(n_594),
.Y(n_635)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_635),
.Y(n_649)
);

BUFx24_ASAP7_75t_SL g637 ( 
.A(n_611),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_600),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_611),
.B(n_592),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_SL g639 ( 
.A1(n_602),
.A2(n_618),
.B(n_599),
.C(n_614),
.Y(n_639)
);

BUFx4f_ASAP7_75t_SL g643 ( 
.A(n_639),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_642),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_626),
.B(n_617),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_623),
.B(n_609),
.C(n_606),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_644),
.B(n_654),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_639),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_601),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_647),
.B(n_640),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_627),
.A2(n_621),
.B(n_620),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_653),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_632),
.A2(n_621),
.B(n_239),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_265),
.C(n_270),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_628),
.B(n_265),
.C(n_238),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_656),
.C(n_639),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_630),
.B(n_2),
.C(n_3),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_649),
.B(n_636),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_657),
.B(n_662),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g669 ( 
.A1(n_658),
.A2(n_648),
.B(n_663),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_643),
.A2(n_625),
.B1(n_633),
.B2(n_639),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_659),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_646),
.A2(n_622),
.B(n_629),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_660),
.A2(n_667),
.B(n_653),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_634),
.Y(n_662)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_650),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_644),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_668),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_652),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_669),
.B(n_670),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_SL g678 ( 
.A1(n_671),
.A2(n_664),
.B(n_668),
.C(n_654),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_659),
.A2(n_645),
.B(n_656),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_673),
.A2(n_664),
.B(n_666),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_661),
.B(n_655),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_674),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_677),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_678),
.B(n_672),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_676),
.A2(n_672),
.B(n_675),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_680),
.A2(n_3),
.B(n_4),
.Y(n_684)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_683),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_684),
.A2(n_679),
.B(n_4),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_685),
.A2(n_682),
.B(n_686),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g688 ( 
.A(n_687),
.B(n_681),
.C(n_3),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_688),
.A2(n_3),
.B(n_635),
.Y(n_689)
);


endmodule