module fake_jpeg_24907_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_59),
.B1(n_26),
.B2(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_25),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_18),
.B1(n_26),
.B2(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_33),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_20),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_57),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_39),
.B1(n_40),
.B2(n_33),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_78),
.B(n_17),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_40),
.B(n_1),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_83),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_40),
.B1(n_35),
.B2(n_23),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_34),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_38),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_34),
.B1(n_63),
.B2(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_34),
.B1(n_23),
.B2(n_29),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_41),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_93),
.B1(n_96),
.B2(n_102),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_94),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_51),
.B1(n_60),
.B2(n_66),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_108),
.B(n_85),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_63),
.C(n_49),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_105),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_104),
.B1(n_87),
.B2(n_47),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_42),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_63),
.C(n_47),
.Y(n_107)
);

NAND2x1_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_42),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_67),
.B1(n_43),
.B2(n_42),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_132),
.B(n_107),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_69),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_99),
.C(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_88),
.B1(n_57),
.B2(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_87),
.B1(n_82),
.B2(n_66),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_50),
.B1(n_85),
.B2(n_43),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_42),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_84),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_43),
.B1(n_23),
.B2(n_31),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_102),
.B1(n_97),
.B2(n_94),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_108),
.C(n_99),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_28),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_31),
.C(n_29),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_146),
.B1(n_117),
.B2(n_119),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_89),
.B1(n_92),
.B2(n_108),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_155),
.B(n_158),
.Y(n_170)
);

NOR4xp25_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_107),
.C(n_103),
.D(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_95),
.B(n_90),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_24),
.B(n_1),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_104),
.B(n_84),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_116),
.B1(n_131),
.B2(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_77),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_114),
.B1(n_120),
.B2(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_178),
.C(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_183),
.Y(n_191)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_144),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_77),
.C(n_24),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_197),
.B(n_198),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_147),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_202),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_208),
.B(n_186),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_162),
.C(n_138),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_176),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_151),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_205),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_146),
.B1(n_141),
.B2(n_15),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_184),
.B1(n_195),
.B2(n_201),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_170),
.B1(n_187),
.B2(n_182),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_225),
.B(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_202),
.C(n_196),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_200),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_203),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_165),
.B(n_196),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_173),
.B(n_172),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_141),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_193),
.B1(n_191),
.B2(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_234),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_179),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_238),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_165),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_174),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_226),
.C(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_249),
.C(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_0),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_212),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_228),
.B1(n_231),
.B2(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_220),
.B1(n_211),
.B2(n_239),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_214),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_213),
.C(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_254),
.B(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_224),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_256),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_2),
.B(n_5),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_248),
.B(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_6),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_246),
.B(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_263),
.B(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_8),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_249),
.B(n_7),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_266),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.C(n_12),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_10),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_268),
.B(n_13),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_272),
.B(n_269),
.Y(n_275)
);

OAI31xp33_ASAP7_75t_SL g276 ( 
.A1(n_275),
.A2(n_14),
.A3(n_12),
.B(n_13),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_14),
.Y(n_277)
);


endmodule