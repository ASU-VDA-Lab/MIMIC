module real_aes_9806_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_1994, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_1994;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1284;
wire n_1987;
wire n_859;
wire n_1465;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1812;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_730;
wire n_1023;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_1457;
wire n_465;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_1969;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_1584;
wire n_466;
wire n_1277;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_0), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_1), .A2(n_189), .B1(n_949), .B2(n_1333), .C(n_1334), .Y(n_1332) );
AOI221xp5_ASAP7_75t_L g1365 ( .A1(n_1), .A2(n_371), .B1(n_622), .B2(n_851), .C(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_2), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_2), .A2(n_361), .B1(n_798), .B2(n_928), .Y(n_1311) );
OA22x2_ASAP7_75t_L g741 ( .A1(n_3), .A2(n_742), .B1(n_816), .B2(n_817), .Y(n_741) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_3), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g1908 ( .A1(n_4), .A2(n_74), .B1(n_1909), .B2(n_1911), .Y(n_1908) );
INVx1_ASAP7_75t_L g1920 ( .A(n_4), .Y(n_1920) );
INVx1_ASAP7_75t_L g1011 ( .A(n_5), .Y(n_1011) );
INVx1_ASAP7_75t_L g1953 ( .A(n_6), .Y(n_1953) );
INVx1_ASAP7_75t_L g1481 ( .A(n_7), .Y(n_1481) );
INVxp33_ASAP7_75t_L g1305 ( .A(n_8), .Y(n_1305) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_8), .A2(n_614), .B(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1716 ( .A(n_9), .Y(n_1716) );
INVx1_ASAP7_75t_L g1916 ( .A(n_10), .Y(n_1916) );
OAI22xp5_ASAP7_75t_L g1931 ( .A1(n_10), .A2(n_93), .B1(n_1013), .B2(n_1017), .Y(n_1931) );
INVx1_ASAP7_75t_L g1293 ( .A(n_11), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_12), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_12), .A2(n_333), .B1(n_999), .B2(n_1000), .Y(n_998) );
INVx1_ASAP7_75t_L g1905 ( .A(n_13), .Y(n_1905) );
OAI221xp5_ASAP7_75t_L g1922 ( .A1(n_13), .A2(n_1088), .B1(n_1108), .B2(n_1923), .C(n_1924), .Y(n_1922) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_14), .A2(n_288), .B1(n_628), .B2(n_833), .C(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g880 ( .A(n_14), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_15), .A2(n_311), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_15), .A2(n_346), .B1(n_798), .B2(n_1222), .Y(n_1221) );
INVxp33_ASAP7_75t_L g1303 ( .A(n_16), .Y(n_1303) );
NAND2xp33_ASAP7_75t_SL g1316 ( .A(n_16), .B(n_1317), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_17), .Y(n_1444) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_18), .A2(n_256), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_18), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_19), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_20), .A2(n_136), .B1(n_1654), .B2(n_1662), .Y(n_1705) );
INVxp67_ASAP7_75t_L g1393 ( .A(n_21), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1414 ( .A1(n_21), .A2(n_66), .B1(n_623), .B2(n_624), .C(n_933), .Y(n_1414) );
INVxp33_ASAP7_75t_L g1956 ( .A(n_22), .Y(n_1956) );
AOI221xp5_ASAP7_75t_L g1976 ( .A1(n_22), .A2(n_89), .B1(n_874), .B2(n_1080), .C(n_1977), .Y(n_1976) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_23), .A2(n_78), .B1(n_599), .B2(n_601), .C(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g655 ( .A(n_23), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g1298 ( .A1(n_24), .A2(n_338), .B1(n_752), .B2(n_895), .C(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1320 ( .A(n_24), .Y(n_1320) );
OAI22xp5_ASAP7_75t_L g1562 ( .A1(n_25), .A2(n_364), .B1(n_441), .B2(n_992), .Y(n_1562) );
INVxp67_ASAP7_75t_SL g1592 ( .A(n_25), .Y(n_1592) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_26), .A2(n_373), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g861 ( .A(n_26), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g1390 ( .A1(n_27), .A2(n_141), .B1(n_895), .B2(n_896), .C(n_1299), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_27), .A2(n_141), .B1(n_829), .B2(n_1211), .Y(n_1412) );
INVx1_ASAP7_75t_L g1520 ( .A(n_28), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_28), .A2(n_60), .B1(n_1044), .B2(n_1548), .Y(n_1547) );
INVxp67_ASAP7_75t_SL g903 ( .A(n_29), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_29), .A2(n_355), .B1(n_472), .B2(n_622), .C(n_624), .Y(n_926) );
INVx1_ASAP7_75t_L g1228 ( .A(n_30), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_31), .A2(n_180), .B1(n_1078), .B2(n_1200), .Y(n_1204) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_31), .Y(n_1218) );
INVxp33_ASAP7_75t_L g1512 ( .A(n_32), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1539 ( .A1(n_32), .A2(n_91), .B1(n_602), .B2(n_995), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1965 ( .A1(n_33), .A2(n_360), .B1(n_1047), .B2(n_1314), .Y(n_1965) );
INVxp67_ASAP7_75t_SL g1983 ( .A(n_33), .Y(n_1983) );
CKINVDCx5p33_ASAP7_75t_R g1424 ( .A(n_34), .Y(n_1424) );
INVx1_ASAP7_75t_L g631 ( .A(n_35), .Y(n_631) );
INVxp33_ASAP7_75t_SL g1019 ( .A(n_36), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_36), .A2(n_149), .B1(n_874), .B2(n_1078), .C(n_1080), .Y(n_1077) );
INVx1_ASAP7_75t_L g380 ( .A(n_37), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_38), .A2(n_129), .B1(n_1654), .B2(n_1662), .Y(n_1726) );
INVx1_ASAP7_75t_L g1688 ( .A(n_39), .Y(n_1688) );
INVx1_ASAP7_75t_L g844 ( .A(n_40), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_40), .A2(n_335), .B1(n_872), .B2(n_874), .Y(n_871) );
INVxp33_ASAP7_75t_SL g952 ( .A(n_41), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_41), .A2(n_297), .B1(n_628), .B2(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1900 ( .A1(n_42), .A2(n_197), .B1(n_702), .B2(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1926 ( .A(n_42), .Y(n_1926) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_43), .A2(n_327), .B1(n_1148), .B2(n_1150), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_43), .A2(n_169), .B1(n_479), .B2(n_702), .C(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1427 ( .A(n_44), .Y(n_1427) );
AOI221xp5_ASAP7_75t_L g1450 ( .A1(n_44), .A2(n_201), .B1(n_618), .B2(n_1451), .C(n_1453), .Y(n_1450) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_45), .A2(n_215), .B1(n_534), .B2(n_545), .C(n_751), .Y(n_1517) );
OAI33xp33_ASAP7_75t_L g1543 ( .A1(n_45), .A2(n_215), .A3(n_487), .B1(n_691), .B2(n_792), .B3(n_1994), .Y(n_1543) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_46), .A2(n_79), .B1(n_534), .B2(n_751), .C(n_752), .Y(n_750) );
OAI222xp33_ASAP7_75t_L g789 ( .A1(n_46), .A2(n_79), .B1(n_246), .B2(n_630), .C1(n_790), .C2(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g1296 ( .A(n_47), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_48), .A2(n_70), .B1(n_441), .B2(n_829), .Y(n_1475) );
OAI221xp5_ASAP7_75t_L g1494 ( .A1(n_48), .A2(n_70), .B1(n_752), .B2(n_895), .C(n_1299), .Y(n_1494) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_49), .A2(n_702), .B(n_704), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_49), .A2(n_100), .B1(n_528), .B2(n_567), .C(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1565 ( .A(n_50), .Y(n_1565) );
OAI221xp5_ASAP7_75t_L g1575 ( .A1(n_50), .A2(n_317), .B1(n_947), .B2(n_949), .C(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1960 ( .A(n_51), .Y(n_1960) );
INVxp33_ASAP7_75t_SL g1195 ( .A(n_52), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_52), .A2(n_170), .B1(n_455), .B2(n_804), .Y(n_1213) );
INVx1_ASAP7_75t_L g856 ( .A(n_53), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_53), .A2(n_344), .B1(n_866), .B2(n_869), .Y(n_868) );
CKINVDCx16_ASAP7_75t_R g1555 ( .A(n_54), .Y(n_1555) );
INVx1_ASAP7_75t_L g1156 ( .A(n_55), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_56), .A2(n_346), .B1(n_566), .B2(n_866), .Y(n_1201) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_56), .A2(n_311), .B1(n_612), .B2(n_624), .C(n_1220), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_57), .A2(n_186), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_1251) );
INVxp33_ASAP7_75t_SL g1266 ( .A(n_57), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1706 ( .A1(n_58), .A2(n_86), .B1(n_1670), .B2(n_1684), .Y(n_1706) );
INVx1_ASAP7_75t_L g1237 ( .A(n_59), .Y(n_1237) );
INVx1_ASAP7_75t_L g1523 ( .A(n_60), .Y(n_1523) );
INVxp67_ASAP7_75t_SL g902 ( .A(n_61), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_61), .A2(n_233), .B1(n_798), .B2(n_928), .Y(n_927) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_62), .A2(n_127), .B1(n_534), .B2(n_545), .C(n_1339), .Y(n_1338) );
OAI221xp5_ASAP7_75t_SL g1362 ( .A1(n_62), .A2(n_127), .B1(n_790), .B2(n_791), .C(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1527 ( .A(n_63), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_64), .Y(n_764) );
XOR2xp5_ASAP7_75t_L g1231 ( .A(n_65), .B(n_1232), .Y(n_1231) );
INVxp33_ASAP7_75t_L g1397 ( .A(n_66), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1967 ( .A1(n_67), .A2(n_222), .B1(n_1968), .B2(n_1969), .Y(n_1967) );
OAI22xp5_ASAP7_75t_L g1989 ( .A1(n_67), .A2(n_222), .B1(n_1111), .B2(n_1113), .Y(n_1989) );
INVx1_ASAP7_75t_L g972 ( .A(n_68), .Y(n_972) );
INVxp67_ASAP7_75t_L g1595 ( .A(n_69), .Y(n_1595) );
XOR2xp5_ASAP7_75t_L g1947 ( .A(n_71), .B(n_1948), .Y(n_1947) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_72), .A2(n_226), .B1(n_999), .B2(n_1000), .Y(n_1570) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_72), .A2(n_226), .B1(n_872), .B2(n_1584), .Y(n_1583) );
AOI22xp33_ASAP7_75t_L g1678 ( .A1(n_73), .A2(n_228), .B1(n_1654), .B2(n_1662), .Y(n_1678) );
INVx1_ASAP7_75t_L g1921 ( .A(n_74), .Y(n_1921) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_75), .A2(n_155), .B1(n_685), .B2(n_691), .C(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g740 ( .A(n_75), .Y(n_740) );
INVxp67_ASAP7_75t_L g1617 ( .A(n_76), .Y(n_1617) );
AOI22xp33_ASAP7_75t_L g1640 ( .A1(n_76), .A2(n_118), .B1(n_714), .B2(n_1162), .Y(n_1640) );
AO22x1_ASAP7_75t_SL g1697 ( .A1(n_77), .A2(n_137), .B1(n_1654), .B2(n_1662), .Y(n_1697) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_78), .A2(n_227), .B1(n_650), .B2(n_652), .C(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g1507 ( .A(n_80), .Y(n_1507) );
INVx1_ASAP7_75t_L g1024 ( .A(n_81), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1441 ( .A(n_82), .Y(n_1441) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_83), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_84), .A2(n_108), .B1(n_1049), .B2(n_1051), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_84), .A2(n_108), .B1(n_1111), .B2(n_1113), .Y(n_1110) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_85), .A2(n_458), .B(n_460), .Y(n_457) );
INVxp33_ASAP7_75t_L g521 ( .A(n_85), .Y(n_521) );
INVx1_ASAP7_75t_L g1035 ( .A(n_87), .Y(n_1035) );
INVxp33_ASAP7_75t_L g1515 ( .A(n_88), .Y(n_1515) );
AOI21xp33_ASAP7_75t_L g1540 ( .A1(n_88), .A2(n_714), .B(n_715), .Y(n_1540) );
INVxp33_ASAP7_75t_L g1957 ( .A(n_89), .Y(n_1957) );
INVx1_ASAP7_75t_L g1623 ( .A(n_90), .Y(n_1623) );
INVxp33_ASAP7_75t_L g1516 ( .A(n_91), .Y(n_1516) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_92), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1917 ( .A1(n_93), .A2(n_367), .B1(n_642), .B2(n_1200), .C(n_1918), .Y(n_1917) );
AOI22xp5_ASAP7_75t_L g1679 ( .A1(n_94), .A2(n_245), .B1(n_1666), .B2(n_1670), .Y(n_1679) );
INVx1_ASAP7_75t_L g1906 ( .A(n_95), .Y(n_1906) );
OAI211xp5_ASAP7_75t_L g1913 ( .A1(n_95), .A2(n_1068), .B(n_1914), .C(n_1919), .Y(n_1913) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_96), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g1907 ( .A1(n_97), .A2(n_249), .B1(n_781), .B2(n_1042), .Y(n_1907) );
OAI22xp5_ASAP7_75t_L g1927 ( .A1(n_97), .A2(n_249), .B1(n_1928), .B2(n_1929), .Y(n_1927) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_98), .A2(n_366), .B1(n_460), .B2(n_779), .C(n_1409), .Y(n_1472) );
INVxp33_ASAP7_75t_L g1490 ( .A(n_98), .Y(n_1490) );
INVxp33_ASAP7_75t_L g1389 ( .A(n_99), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_99), .A2(n_374), .B1(n_798), .B2(n_1411), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_100), .A2(n_254), .B1(n_602), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_101), .A2(n_194), .B1(n_627), .B2(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g665 ( .A(n_101), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_102), .A2(n_115), .B1(n_566), .B2(n_1148), .Y(n_1152) );
INVx1_ASAP7_75t_L g1182 ( .A(n_102), .Y(n_1182) );
OAI221xp5_ASAP7_75t_SL g946 ( .A1(n_103), .A2(n_297), .B1(n_947), .B2(n_949), .C(n_951), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_103), .A2(n_316), .B1(n_460), .B2(n_981), .C(n_985), .Y(n_980) );
INVxp33_ASAP7_75t_SL g1573 ( .A(n_104), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_104), .A2(n_362), .B1(n_1584), .B2(n_1586), .Y(n_1588) );
OAI221xp5_ASAP7_75t_L g1429 ( .A1(n_105), .A2(n_176), .B1(n_534), .B2(n_544), .C(n_1299), .Y(n_1429) );
OAI22xp33_ASAP7_75t_L g1449 ( .A1(n_105), .A2(n_176), .B1(n_830), .B2(n_992), .Y(n_1449) );
AOI22xp5_ASAP7_75t_L g1665 ( .A1(n_106), .A2(n_124), .B1(n_1666), .B2(n_1670), .Y(n_1665) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_107), .A2(n_318), .B1(n_618), .B2(n_1480), .Y(n_1479) );
INVxp67_ASAP7_75t_SL g1502 ( .A(n_107), .Y(n_1502) );
INVx1_ASAP7_75t_L g939 ( .A(n_109), .Y(n_939) );
AOI22xp33_ASAP7_75t_SL g1473 ( .A1(n_110), .A2(n_242), .B1(n_617), .B2(n_798), .Y(n_1473) );
INVxp33_ASAP7_75t_SL g1493 ( .A(n_110), .Y(n_1493) );
OR2x2_ASAP7_75t_L g409 ( .A(n_111), .B(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g413 ( .A(n_111), .Y(n_413) );
BUFx2_ASAP7_75t_L g501 ( .A(n_111), .Y(n_501) );
INVx1_ASAP7_75t_L g513 ( .A(n_111), .Y(n_513) );
INVx1_ASAP7_75t_L g1692 ( .A(n_112), .Y(n_1692) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_113), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_114), .A2(n_248), .B1(n_470), .B2(n_473), .C(n_477), .Y(n_469) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_114), .Y(n_564) );
INVx1_ASAP7_75t_L g1159 ( .A(n_115), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_116), .A2(n_313), .B1(n_1654), .B2(n_1662), .Y(n_1674) );
AOI221xp5_ASAP7_75t_SL g611 ( .A1(n_117), .A2(n_123), .B1(n_460), .B2(n_612), .C(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g644 ( .A(n_117), .Y(n_644) );
INVxp33_ASAP7_75t_L g1608 ( .A(n_118), .Y(n_1608) );
INVx1_ASAP7_75t_L g606 ( .A(n_119), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g1417 ( .A1(n_120), .A2(n_1418), .B1(n_1461), .B2(n_1462), .Y(n_1417) );
INVx1_ASAP7_75t_L g1461 ( .A(n_120), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1727 ( .A1(n_120), .A2(n_273), .B1(n_1670), .B2(n_1684), .Y(n_1727) );
INVx1_ASAP7_75t_L g1350 ( .A(n_121), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_122), .A2(n_203), .B1(n_534), .B2(n_896), .C(n_956), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_122), .A2(n_203), .B1(n_441), .B2(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g641 ( .A(n_123), .Y(n_641) );
XOR2x2_ASAP7_75t_L g676 ( .A(n_124), .B(n_677), .Y(n_676) );
INVxp67_ASAP7_75t_SL g1524 ( .A(n_125), .Y(n_1524) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_125), .A2(n_324), .B1(n_704), .B2(n_1049), .C(n_1546), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_126), .A2(n_246), .B1(n_408), .B2(n_748), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_126), .Y(n_808) );
INVx1_ASAP7_75t_L g1629 ( .A(n_128), .Y(n_1629) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_130), .Y(n_1358) );
INVxp67_ASAP7_75t_L g1604 ( .A(n_131), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g1634 ( .A1(n_131), .A2(n_161), .B1(n_628), .B2(n_995), .Y(n_1634) );
INVx1_ASAP7_75t_L g1700 ( .A(n_132), .Y(n_1700) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_133), .A2(n_278), .B1(n_455), .B2(n_712), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g716 ( .A1(n_133), .A2(n_717), .B(n_719), .C(n_721), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_134), .A2(n_200), .B1(n_441), .B2(n_1239), .Y(n_1238) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_134), .A2(n_200), .B1(n_751), .B2(n_752), .C(n_895), .Y(n_1273) );
INVx1_ASAP7_75t_L g1643 ( .A(n_135), .Y(n_1643) );
INVx1_ASAP7_75t_L g1885 ( .A(n_136), .Y(n_1885) );
AOI22xp33_ASAP7_75t_L g1941 ( .A1(n_136), .A2(n_1942), .B1(n_1946), .B2(n_1990), .Y(n_1941) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_138), .A2(n_206), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_138), .A2(n_194), .B1(n_660), .B2(n_662), .C(n_664), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_139), .A2(n_345), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_139), .Y(n_1105) );
XNOR2x1_ASAP7_75t_L g1380 ( .A(n_140), .B(n_1381), .Y(n_1380) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_142), .A2(n_358), .B1(n_866), .B2(n_1203), .Y(n_1202) );
INVxp33_ASAP7_75t_L g1227 ( .A(n_142), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_143), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_144), .A2(n_329), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_144), .A2(n_205), .B1(n_642), .B2(n_732), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_145), .A2(n_328), .B1(n_479), .B2(n_846), .C(n_848), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_145), .A2(n_240), .B1(n_866), .B2(n_867), .Y(n_865) );
INVxp67_ASAP7_75t_L g1603 ( .A(n_146), .Y(n_1603) );
AOI221xp5_ASAP7_75t_L g1633 ( .A1(n_146), .A2(n_210), .B1(n_458), .B2(n_460), .C(n_1409), .Y(n_1633) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_147), .A2(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g722 ( .A(n_147), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_148), .A2(n_205), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_148), .A2(n_329), .B1(n_508), .B2(n_730), .Y(n_729) );
INVxp33_ASAP7_75t_SL g1015 ( .A(n_149), .Y(n_1015) );
XNOR2xp5_ASAP7_75t_L g1006 ( .A(n_150), .B(n_1007), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g894 ( .A1(n_151), .A2(n_191), .B1(n_541), .B2(n_895), .C(n_896), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_151), .A2(n_191), .B1(n_436), .B2(n_937), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g1569 ( .A1(n_152), .A2(n_325), .B1(n_623), .B2(n_996), .C(n_997), .Y(n_1569) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_152), .A2(n_325), .B1(n_1586), .B2(n_1587), .Y(n_1585) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_153), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g1605 ( .A1(n_154), .A2(n_198), .B1(n_534), .B2(n_751), .C(n_752), .Y(n_1605) );
OAI22xp5_ASAP7_75t_L g1635 ( .A1(n_154), .A2(n_198), .B1(n_1211), .B2(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g720 ( .A(n_155), .Y(n_720) );
INVx1_ASAP7_75t_L g609 ( .A(n_156), .Y(n_609) );
INVx1_ASAP7_75t_L g1246 ( .A(n_157), .Y(n_1246) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_158), .Y(n_771) );
INVx1_ASAP7_75t_L g1329 ( .A(n_159), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_160), .Y(n_1446) );
INVxp67_ASAP7_75t_L g1600 ( .A(n_161), .Y(n_1600) );
INVx1_ASAP7_75t_L g1400 ( .A(n_162), .Y(n_1400) );
INVxp33_ASAP7_75t_SL g1572 ( .A(n_163), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_163), .A2(n_305), .B1(n_872), .B2(n_1587), .Y(n_1589) );
INVx1_ASAP7_75t_L g1658 ( .A(n_164), .Y(n_1658) );
INVx1_ASAP7_75t_L g1131 ( .A(n_165), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_165), .A2(n_275), .B1(n_830), .B2(n_992), .Y(n_1160) );
XNOR2x1_ASAP7_75t_L g1183 ( .A(n_166), .B(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1255 ( .A(n_167), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_168), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_169), .A2(n_326), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
INVxp33_ASAP7_75t_SL g1190 ( .A(n_170), .Y(n_1190) );
XOR2x1_ASAP7_75t_L g1124 ( .A(n_171), .B(n_1125), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1682 ( .A1(n_171), .A2(n_260), .B1(n_1683), .B2(n_1685), .C(n_1687), .Y(n_1682) );
INVx1_ASAP7_75t_L g1513 ( .A(n_172), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_172), .B(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1353 ( .A(n_173), .Y(n_1353) );
INVx1_ASAP7_75t_L g1961 ( .A(n_174), .Y(n_1961) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_175), .A2(n_218), .B1(n_618), .B2(n_1241), .C(n_1243), .Y(n_1240) );
INVxp33_ASAP7_75t_L g1276 ( .A(n_175), .Y(n_1276) );
INVx1_ASAP7_75t_L g1402 ( .A(n_177), .Y(n_1402) );
INVx1_ASAP7_75t_L g1659 ( .A(n_178), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_178), .B(n_1657), .Y(n_1664) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_179), .A2(n_261), .B1(n_617), .B2(n_618), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_179), .A2(n_261), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_637) );
INVxp33_ASAP7_75t_L g1226 ( .A(n_180), .Y(n_1226) );
AOI22xp33_ASAP7_75t_SL g1964 ( .A1(n_181), .A2(n_213), .B1(n_1042), .B2(n_1045), .Y(n_1964) );
INVxp67_ASAP7_75t_SL g1982 ( .A(n_181), .Y(n_1982) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_182), .A2(n_240), .B1(n_851), .B2(n_853), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_182), .A2(n_328), .B1(n_642), .B2(n_864), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_183), .A2(n_458), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g879 ( .A(n_183), .Y(n_879) );
INVx1_ASAP7_75t_L g1297 ( .A(n_184), .Y(n_1297) );
INVx2_ASAP7_75t_L g392 ( .A(n_185), .Y(n_392) );
INVxp67_ASAP7_75t_L g1259 ( .A(n_186), .Y(n_1259) );
AO221x2_ASAP7_75t_L g1712 ( .A1(n_187), .A2(n_236), .B1(n_1684), .B2(n_1713), .C(n_1714), .Y(n_1712) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_188), .A2(n_347), .B1(n_429), .B2(n_624), .C(n_1478), .Y(n_1477) );
INVxp33_ASAP7_75t_SL g1498 ( .A(n_188), .Y(n_1498) );
INVx1_ASAP7_75t_L g1364 ( .A(n_189), .Y(n_1364) );
BUFx3_ASAP7_75t_L g422 ( .A(n_190), .Y(n_422) );
INVx1_ASAP7_75t_L g451 ( .A(n_190), .Y(n_451) );
INVx1_ASAP7_75t_L g1432 ( .A(n_192), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_192), .A2(n_307), .B1(n_1044), .B2(n_1314), .Y(n_1458) );
INVx1_ASAP7_75t_L g1954 ( .A(n_193), .Y(n_1954) );
INVx1_ASAP7_75t_L g1529 ( .A(n_195), .Y(n_1529) );
INVxp33_ASAP7_75t_L g892 ( .A(n_196), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_196), .A2(n_244), .B1(n_714), .B2(n_715), .C(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1925 ( .A(n_197), .Y(n_1925) );
INVxp33_ASAP7_75t_L g1306 ( .A(n_199), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_199), .A2(n_314), .B1(n_1026), .B2(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1422 ( .A(n_201), .Y(n_1422) );
INVx1_ASAP7_75t_L g1192 ( .A(n_202), .Y(n_1192) );
INVx1_ASAP7_75t_L g1254 ( .A(n_204), .Y(n_1254) );
INVx1_ASAP7_75t_L g666 ( .A(n_206), .Y(n_666) );
INVxp67_ASAP7_75t_L g1343 ( .A(n_207), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_207), .A2(n_343), .B1(n_999), .B2(n_1314), .Y(n_1375) );
OAI221xp5_ASAP7_75t_SL g435 ( .A1(n_208), .A2(n_365), .B1(n_436), .B2(n_441), .C(n_445), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_208), .A2(n_365), .B1(n_534), .B2(n_541), .C(n_544), .Y(n_533) );
INVx1_ASAP7_75t_L g1336 ( .A(n_209), .Y(n_1336) );
INVxp67_ASAP7_75t_L g1601 ( .A(n_210), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_211), .A2(n_351), .B1(n_851), .B2(n_853), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1262 ( .A(n_211), .Y(n_1262) );
INVx1_ASAP7_75t_L g608 ( .A(n_212), .Y(n_608) );
INVxp67_ASAP7_75t_SL g1987 ( .A(n_213), .Y(n_1987) );
INVx1_ASAP7_75t_L g1250 ( .A(n_214), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_216), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g1972 ( .A(n_217), .Y(n_1972) );
INVxp33_ASAP7_75t_L g1279 ( .A(n_218), .Y(n_1279) );
INVx1_ASAP7_75t_L g1234 ( .A(n_219), .Y(n_1234) );
INVx1_ASAP7_75t_L g1324 ( .A(n_220), .Y(n_1324) );
INVx1_ASAP7_75t_L g1139 ( .A(n_221), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_221), .A2(n_315), .B1(n_617), .B2(n_1162), .C(n_1163), .Y(n_1161) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_223), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_223), .A2(n_276), .B1(n_779), .B2(n_798), .Y(n_1415) );
INVx1_ASAP7_75t_L g494 ( .A(n_224), .Y(n_494) );
INVx1_ASAP7_75t_L g417 ( .A(n_225), .Y(n_417) );
INVx1_ASAP7_75t_L g462 ( .A(n_225), .Y(n_462) );
INVx1_ASAP7_75t_L g605 ( .A(n_227), .Y(n_605) );
INVxp33_ASAP7_75t_SL g889 ( .A(n_229), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_229), .A2(n_234), .B1(n_623), .B2(n_935), .Y(n_934) );
INVxp33_ASAP7_75t_SL g1194 ( .A(n_230), .Y(n_1194) );
AOI21xp33_ASAP7_75t_L g1214 ( .A1(n_230), .A2(n_840), .B(n_930), .Y(n_1214) );
INVx1_ASAP7_75t_L g1526 ( .A(n_231), .Y(n_1526) );
INVx1_ASAP7_75t_L g1474 ( .A(n_232), .Y(n_1474) );
INVx1_ASAP7_75t_L g907 ( .A(n_233), .Y(n_907) );
INVxp33_ASAP7_75t_SL g893 ( .A(n_234), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_235), .Y(n_708) );
INVx1_ASAP7_75t_L g1399 ( .A(n_237), .Y(n_1399) );
AOI22xp33_ASAP7_75t_SL g1966 ( .A1(n_238), .A2(n_300), .B1(n_985), .B2(n_1045), .Y(n_1966) );
OAI211xp5_ASAP7_75t_SL g1974 ( .A1(n_238), .A2(n_1068), .B(n_1975), .C(n_1979), .Y(n_1974) );
AOI22xp5_ASAP7_75t_L g1653 ( .A1(n_239), .A2(n_287), .B1(n_1654), .B2(n_1662), .Y(n_1653) );
INVx1_ASAP7_75t_L g882 ( .A(n_241), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g1675 ( .A1(n_241), .A2(n_312), .B1(n_1666), .B2(n_1670), .Y(n_1675) );
INVxp33_ASAP7_75t_L g1489 ( .A(n_242), .Y(n_1489) );
INVx1_ASAP7_75t_L g1915 ( .A(n_243), .Y(n_1915) );
OAI22xp5_ASAP7_75t_L g1932 ( .A1(n_243), .A2(n_367), .B1(n_1933), .B2(n_1935), .Y(n_1932) );
INVxp33_ASAP7_75t_L g890 ( .A(n_244), .Y(n_890) );
INVx1_ASAP7_75t_L g1403 ( .A(n_247), .Y(n_1403) );
INVx1_ASAP7_75t_L g559 ( .A(n_248), .Y(n_559) );
INVxp67_ASAP7_75t_L g1614 ( .A(n_250), .Y(n_1614) );
AOI221xp5_ASAP7_75t_L g1638 ( .A1(n_250), .A2(n_264), .B1(n_454), .B2(n_1457), .C(n_1639), .Y(n_1638) );
INVxp33_ASAP7_75t_L g1290 ( .A(n_251), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_251), .A2(n_283), .B1(n_472), .B2(n_624), .C(n_933), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_252), .A2(n_319), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g553 ( .A(n_252), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_253), .A2(n_330), .B1(n_1045), .B2(n_1047), .Y(n_1046) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_253), .A2(n_1088), .B1(n_1090), .B2(n_1100), .C(n_1108), .Y(n_1087) );
INVx1_ASAP7_75t_L g735 ( .A(n_254), .Y(n_735) );
INVx1_ASAP7_75t_L g943 ( .A(n_255), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_256), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_257), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g1715 ( .A(n_258), .Y(n_1715) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_259), .A2(n_301), .B1(n_874), .B2(n_1144), .Y(n_1153) );
INVx1_ASAP7_75t_L g1181 ( .A(n_259), .Y(n_1181) );
INVxp67_ASAP7_75t_SL g964 ( .A(n_262), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_262), .A2(n_299), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_994) );
INVx1_ASAP7_75t_L g973 ( .A(n_263), .Y(n_973) );
INVxp33_ASAP7_75t_L g1612 ( .A(n_264), .Y(n_1612) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_265), .A2(n_271), .B1(n_454), .B2(n_455), .Y(n_453) );
INVxp33_ASAP7_75t_L g526 ( .A(n_265), .Y(n_526) );
INVx1_ASAP7_75t_L g1436 ( .A(n_266), .Y(n_1436) );
AOI221xp5_ASAP7_75t_L g1456 ( .A1(n_266), .A2(n_284), .B1(n_702), .B2(n_1173), .C(n_1457), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_267), .Y(n_1405) );
INVx1_ASAP7_75t_L g1351 ( .A(n_268), .Y(n_1351) );
BUFx3_ASAP7_75t_L g424 ( .A(n_269), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_269), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_270), .Y(n_759) );
INVxp33_ASAP7_75t_L g505 ( .A(n_271), .Y(n_505) );
INVx1_ASAP7_75t_L g589 ( .A(n_272), .Y(n_589) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_274), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_274), .B(n_354), .Y(n_410) );
AND2x2_ASAP7_75t_L g514 ( .A(n_274), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g588 ( .A(n_274), .Y(n_588) );
INVx1_ASAP7_75t_L g1130 ( .A(n_275), .Y(n_1130) );
INVxp67_ASAP7_75t_L g1394 ( .A(n_276), .Y(n_1394) );
INVx1_ASAP7_75t_L g970 ( .A(n_277), .Y(n_970) );
INVx1_ASAP7_75t_L g725 ( .A(n_278), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g1566 ( .A1(n_279), .A2(n_1319), .B(n_1542), .Y(n_1566) );
INVx1_ASAP7_75t_L g1578 ( .A(n_279), .Y(n_1578) );
OAI332xp33_ASAP7_75t_L g753 ( .A1(n_280), .A2(n_547), .A3(n_584), .B1(n_754), .B2(n_758), .B3(n_763), .C1(n_770), .C2(n_775), .Y(n_753) );
INVx1_ASAP7_75t_L g812 ( .A(n_280), .Y(n_812) );
INVx1_ASAP7_75t_L g968 ( .A(n_281), .Y(n_968) );
INVx1_ASAP7_75t_L g1245 ( .A(n_282), .Y(n_1245) );
INVxp67_ASAP7_75t_L g1286 ( .A(n_283), .Y(n_1286) );
INVx1_ASAP7_75t_L g1434 ( .A(n_284), .Y(n_1434) );
INVx1_ASAP7_75t_L g1483 ( .A(n_285), .Y(n_1483) );
INVx2_ASAP7_75t_L g419 ( .A(n_286), .Y(n_419) );
OR2x2_ASAP7_75t_L g433 ( .A(n_286), .B(n_417), .Y(n_433) );
INVx1_ASAP7_75t_L g876 ( .A(n_288), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_289), .Y(n_756) );
INVx1_ASAP7_75t_L g1621 ( .A(n_290), .Y(n_1621) );
INVxp67_ASAP7_75t_L g1347 ( .A(n_291), .Y(n_1347) );
AOI221xp5_ASAP7_75t_L g1371 ( .A1(n_291), .A2(n_341), .B1(n_1372), .B2(n_1373), .C(n_1374), .Y(n_1371) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_292), .Y(n_594) );
INVx1_ASAP7_75t_L g911 ( .A(n_293), .Y(n_911) );
INVx1_ASAP7_75t_L g857 ( .A(n_294), .Y(n_857) );
INVx1_ASAP7_75t_L g1484 ( .A(n_295), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_296), .A2(n_302), .B1(n_781), .B2(n_1042), .Y(n_1041) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_296), .Y(n_1094) );
INVx1_ASAP7_75t_L g468 ( .A(n_298), .Y(n_468) );
INVxp33_ASAP7_75t_SL g962 ( .A(n_299), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g1980 ( .A1(n_300), .A2(n_1088), .B1(n_1108), .B2(n_1981), .C(n_1984), .Y(n_1980) );
INVx1_ASAP7_75t_L g1171 ( .A(n_301), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1091 ( .A(n_302), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_303), .Y(n_1138) );
INVx1_ASAP7_75t_L g1354 ( .A(n_304), .Y(n_1354) );
INVxp67_ASAP7_75t_SL g1568 ( .A(n_305), .Y(n_1568) );
AOI221xp5_ASAP7_75t_L g1563 ( .A1(n_306), .A2(n_317), .B1(n_623), .B2(n_1000), .C(n_1564), .Y(n_1563) );
INVxp33_ASAP7_75t_L g1577 ( .A(n_306), .Y(n_1577) );
INVx1_ASAP7_75t_L g1438 ( .A(n_307), .Y(n_1438) );
INVx1_ASAP7_75t_L g1505 ( .A(n_308), .Y(n_1505) );
INVx1_ASAP7_75t_L g1029 ( .A(n_309), .Y(n_1029) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_310), .Y(n_1426) );
INVxp33_ASAP7_75t_L g1302 ( .A(n_314), .Y(n_1302) );
INVx1_ASAP7_75t_L g1134 ( .A(n_315), .Y(n_1134) );
INVxp33_ASAP7_75t_SL g953 ( .A(n_316), .Y(n_953) );
INVxp33_ASAP7_75t_L g1497 ( .A(n_318), .Y(n_1497) );
INVx1_ASAP7_75t_L g568 ( .A(n_319), .Y(n_568) );
INVx1_ASAP7_75t_L g1294 ( .A(n_320), .Y(n_1294) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_321), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_321), .A2(n_348), .B1(n_436), .B2(n_1211), .C(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1531 ( .A(n_322), .Y(n_1531) );
CKINVDCx5p33_ASAP7_75t_R g1440 ( .A(n_323), .Y(n_1440) );
INVxp33_ASAP7_75t_L g1521 ( .A(n_324), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_326), .A2(n_327), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
OAI211xp5_ASAP7_75t_SL g1067 ( .A1(n_330), .A2(n_1068), .B(n_1073), .C(n_1082), .Y(n_1067) );
INVx1_ASAP7_75t_L g1628 ( .A(n_331), .Y(n_1628) );
INVx1_ASAP7_75t_L g1485 ( .A(n_332), .Y(n_1485) );
INVxp67_ASAP7_75t_SL g965 ( .A(n_333), .Y(n_965) );
INVx1_ASAP7_75t_L g446 ( .A(n_334), .Y(n_446) );
INVx1_ASAP7_75t_L g855 ( .A(n_335), .Y(n_855) );
INVx1_ASAP7_75t_L g884 ( .A(n_336), .Y(n_884) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_337), .B(n_380), .Y(n_1661) );
AND3x2_ASAP7_75t_L g1667 ( .A(n_337), .B(n_380), .C(n_1658), .Y(n_1667) );
INVx1_ASAP7_75t_L g1321 ( .A(n_338), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g1888 ( .A(n_339), .Y(n_1888) );
INVx2_ASAP7_75t_L g393 ( .A(n_340), .Y(n_393) );
INVxp67_ASAP7_75t_SL g1348 ( .A(n_341), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_342), .Y(n_1136) );
INVxp33_ASAP7_75t_SL g1345 ( .A(n_343), .Y(n_1345) );
INVx1_ASAP7_75t_L g827 ( .A(n_344), .Y(n_827) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_345), .Y(n_1102) );
INVxp67_ASAP7_75t_SL g1501 ( .A(n_347), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g1188 ( .A(n_348), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g1899 ( .A(n_349), .Y(n_1899) );
AOI22x1_ASAP7_75t_L g1280 ( .A1(n_350), .A2(n_1281), .B1(n_1282), .B2(n_1325), .Y(n_1280) );
INVx1_ASAP7_75t_L g1325 ( .A(n_350), .Y(n_1325) );
INVxp33_ASAP7_75t_L g1264 ( .A(n_351), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_352), .Y(n_755) );
INVx1_ASAP7_75t_L g914 ( .A(n_353), .Y(n_914) );
INVx1_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
INVx2_ASAP7_75t_L g515 ( .A(n_354), .Y(n_515) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_355), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g1896 ( .A(n_356), .Y(n_1896) );
INVxp33_ASAP7_75t_L g1388 ( .A(n_357), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_357), .A2(n_359), .B1(n_460), .B2(n_614), .C(n_1409), .Y(n_1408) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_358), .Y(n_1209) );
INVxp33_ASAP7_75t_L g1386 ( .A(n_359), .Y(n_1386) );
INVxp67_ASAP7_75t_SL g1988 ( .A(n_360), .Y(n_1988) );
INVxp33_ASAP7_75t_L g1289 ( .A(n_361), .Y(n_1289) );
INVxp67_ASAP7_75t_SL g1561 ( .A(n_362), .Y(n_1561) );
INVx1_ASAP7_75t_L g912 ( .A(n_363), .Y(n_912) );
INVxp67_ASAP7_75t_SL g1591 ( .A(n_364), .Y(n_1591) );
INVxp33_ASAP7_75t_L g1492 ( .A(n_366), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g1558 ( .A(n_368), .Y(n_1558) );
INVx1_ASAP7_75t_L g490 ( .A(n_369), .Y(n_490) );
INVx1_ASAP7_75t_L g915 ( .A(n_370), .Y(n_915) );
INVxp33_ASAP7_75t_SL g1335 ( .A(n_371), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_372), .Y(n_838) );
INVx1_ASAP7_75t_L g860 ( .A(n_373), .Y(n_860) );
INVxp33_ASAP7_75t_L g1385 ( .A(n_374), .Y(n_1385) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_396), .B(n_1646), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_383), .Y(n_377) );
AND2x4_ASAP7_75t_L g1940 ( .A(n_378), .B(n_384), .Y(n_1940) );
NOR2xp33_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_SL g1945 ( .A(n_379), .Y(n_1945) );
NAND2xp5_ASAP7_75t_L g1992 ( .A(n_379), .B(n_381), .Y(n_1992) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g1944 ( .A(n_381), .B(n_1945), .Y(n_1944) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g658 ( .A(n_387), .B(n_395), .Y(n_658) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g548 ( .A(n_388), .B(n_549), .Y(n_548) );
OR2x6_ASAP7_75t_L g389 ( .A(n_390), .B(n_394), .Y(n_389) );
OR2x2_ASAP7_75t_L g408 ( .A(n_390), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g552 ( .A(n_390), .Y(n_552) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_390), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_390), .A2(n_696), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx2_ASAP7_75t_SL g960 ( .A(n_390), .Y(n_960) );
INVx2_ASAP7_75t_SL g1104 ( .A(n_390), .Y(n_1104) );
BUFx2_ASAP7_75t_L g1611 ( .A(n_390), .Y(n_1611) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x4_ASAP7_75t_L g510 ( .A(n_392), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g519 ( .A(n_392), .Y(n_519) );
AND2x2_ASAP7_75t_L g525 ( .A(n_392), .B(n_393), .Y(n_525) );
INVx2_ASAP7_75t_L g530 ( .A(n_392), .Y(n_530) );
INVx1_ASAP7_75t_L g558 ( .A(n_392), .Y(n_558) );
INVx2_ASAP7_75t_L g511 ( .A(n_393), .Y(n_511) );
INVx1_ASAP7_75t_L g532 ( .A(n_393), .Y(n_532) );
INVx1_ASAP7_75t_L g539 ( .A(n_393), .Y(n_539) );
INVx1_ASAP7_75t_L g557 ( .A(n_393), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_393), .B(n_530), .Y(n_563) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_1117), .B2(n_1118), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AO22x1_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_819), .B2(n_820), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_590), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
XNOR2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_589), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_502), .Y(n_404) );
AOI21xp33_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_425), .B(n_426), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_406), .A2(n_499), .B1(n_825), .B2(n_857), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g1205 ( .A1(n_406), .A2(n_1206), .B1(n_1207), .B2(n_1228), .Y(n_1205) );
AOI21xp33_ASAP7_75t_L g1233 ( .A1(n_406), .A2(n_1234), .B(n_1235), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_406), .A2(n_1206), .B1(n_1308), .B2(n_1324), .Y(n_1307) );
INVx1_ASAP7_75t_L g1357 ( .A(n_406), .Y(n_1357) );
AOI21xp33_ASAP7_75t_SL g1404 ( .A1(n_406), .A2(n_1405), .B(n_1406), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_406), .A2(n_1206), .B1(n_1470), .B2(n_1485), .Y(n_1469) );
INVx5_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g940 ( .A(n_407), .Y(n_940) );
INVx1_ASAP7_75t_L g1155 ( .A(n_407), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1642 ( .A(n_407), .Y(n_1642) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
INVx2_ASAP7_75t_L g667 ( .A(n_408), .Y(n_667) );
INVx3_ASAP7_75t_L g540 ( .A(n_409), .Y(n_540) );
INVx1_ASAP7_75t_L g1065 ( .A(n_410), .Y(n_1065) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x6_ASAP7_75t_L g1060 ( .A(n_412), .B(n_1061), .Y(n_1060) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
AND2x4_ASAP7_75t_L g1053 ( .A(n_413), .B(n_461), .Y(n_1053) );
INVx2_ASAP7_75t_L g630 ( .A(n_414), .Y(n_630) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_420), .Y(n_414) );
AND2x4_ASAP7_75t_L g437 ( .A(n_415), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g442 ( .A(n_415), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g487 ( .A(n_415), .Y(n_487) );
AND2x4_ASAP7_75t_L g607 ( .A(n_415), .B(n_438), .Y(n_607) );
BUFx2_ASAP7_75t_L g694 ( .A(n_415), .Y(n_694) );
AND2x2_ASAP7_75t_L g831 ( .A(n_415), .B(n_443), .Y(n_831) );
AND2x4_ASAP7_75t_L g938 ( .A(n_415), .B(n_443), .Y(n_938) );
NAND2x1p5_ASAP7_75t_L g1034 ( .A(n_415), .B(n_585), .Y(n_1034) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g461 ( .A(n_418), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g480 ( .A(n_419), .B(n_462), .Y(n_480) );
INVx6_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
BUFx2_ASAP7_75t_L g714 ( .A(n_420), .Y(n_714) );
INVx2_ASAP7_75t_L g1022 ( .A(n_420), .Y(n_1022) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g444 ( .A(n_421), .Y(n_444) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g430 ( .A(n_422), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_424), .Y(n_467) );
INVx1_ASAP7_75t_L g440 ( .A(n_423), .Y(n_440) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g456 ( .A(n_424), .B(n_451), .Y(n_456) );
AOI31xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_463), .A3(n_489), .B(n_498), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_434), .B(n_435), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_428), .A2(n_491), .B1(n_855), .B2(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g990 ( .A(n_428), .Y(n_990) );
AOI211xp5_ASAP7_75t_L g1158 ( .A1(n_428), .A2(n_1159), .B(n_1160), .C(n_1161), .Y(n_1158) );
AOI21xp33_ASAP7_75t_L g1208 ( .A1(n_428), .A2(n_1209), .B(n_1210), .Y(n_1208) );
AOI211xp5_ASAP7_75t_L g1236 ( .A1(n_428), .A2(n_1237), .B(n_1238), .C(n_1240), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_428), .A2(n_491), .B1(n_1293), .B2(n_1296), .Y(n_1322) );
HB1xp67_ASAP7_75t_L g1361 ( .A(n_428), .Y(n_1361) );
AOI221xp5_ASAP7_75t_L g1407 ( .A1(n_428), .A2(n_1399), .B1(n_1408), .B2(n_1410), .C(n_1412), .Y(n_1407) );
AOI211xp5_ASAP7_75t_L g1448 ( .A1(n_428), .A2(n_1441), .B(n_1449), .C(n_1450), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_428), .A2(n_1472), .B1(n_1473), .B2(n_1474), .C(n_1475), .Y(n_1471) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .Y(n_428) );
BUFx3_ASAP7_75t_L g617 ( .A(n_429), .Y(n_617) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_429), .Y(n_1050) );
INVx1_ASAP7_75t_L g1452 ( .A(n_429), .Y(n_1452) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_430), .Y(n_454) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
BUFx2_ASAP7_75t_L g623 ( .A(n_430), .Y(n_623) );
INVx2_ASAP7_75t_SL g703 ( .A(n_430), .Y(n_703) );
BUFx3_ASAP7_75t_L g712 ( .A(n_430), .Y(n_712) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_430), .Y(n_804) );
BUFx2_ASAP7_75t_L g995 ( .A(n_430), .Y(n_995) );
INVx1_ASAP7_75t_L g452 ( .A(n_431), .Y(n_452) );
AND2x4_ASAP7_75t_L g465 ( .A(n_432), .B(n_466), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_432), .A2(n_442), .B1(n_598), .B2(n_607), .C1(n_608), .C2(n_609), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_432), .A2(n_680), .B(n_683), .Y(n_679) );
AND2x2_ASAP7_75t_L g924 ( .A(n_432), .B(n_472), .Y(n_924) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g492 ( .A(n_433), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g496 ( .A(n_433), .B(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_SL g777 ( .A1(n_433), .A2(n_778), .B(n_783), .C(n_788), .Y(n_777) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_433), .B(n_513), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_434), .A2(n_494), .B1(n_570), .B2(n_573), .Y(n_569) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx4_ASAP7_75t_L g1636 ( .A(n_437), .Y(n_1636) );
INVxp67_ASAP7_75t_L g691 ( .A(n_438), .Y(n_691) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g1032 ( .A(n_439), .Y(n_1032) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g692 ( .A(n_443), .Y(n_692) );
INVx2_ASAP7_75t_L g792 ( .A(n_443), .Y(n_792) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_453), .C(n_457), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_446), .A2(n_505), .B1(n_506), .B2(n_516), .Y(n_504) );
OAI211xp5_ASAP7_75t_L g1212 ( .A1(n_447), .A2(n_1192), .B(n_1213), .C(n_1214), .Y(n_1212) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g685 ( .A(n_448), .Y(n_685) );
INVx1_ASAP7_75t_L g1164 ( .A(n_448), .Y(n_1164) );
BUFx4f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g698 ( .A(n_449), .Y(n_698) );
INVx1_ASAP7_75t_L g801 ( .A(n_449), .Y(n_801) );
BUFx2_ASAP7_75t_L g837 ( .A(n_449), .Y(n_837) );
INVx1_ASAP7_75t_L g1244 ( .A(n_449), .Y(n_1244) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
OR2x2_ASAP7_75t_L g493 ( .A(n_450), .B(n_452), .Y(n_493) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g834 ( .A(n_454), .Y(n_834) );
BUFx2_ASAP7_75t_L g1372 ( .A(n_454), .Y(n_1372) );
BUFx3_ASAP7_75t_L g1968 ( .A(n_454), .Y(n_1968) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_455), .Y(n_798) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_455), .Y(n_1051) );
INVx1_ASAP7_75t_L g1970 ( .A(n_455), .Y(n_1970) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_456), .Y(n_484) );
INVx2_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
INVx1_ASAP7_75t_L g619 ( .A(n_456), .Y(n_619) );
INVx1_ASAP7_75t_L g782 ( .A(n_456), .Y(n_782) );
BUFx3_ASAP7_75t_L g482 ( .A(n_458), .Y(n_482) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g615 ( .A(n_459), .Y(n_615) );
INVx1_ASAP7_75t_L g627 ( .A(n_459), .Y(n_627) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_459), .Y(n_689) );
INVx1_ASAP7_75t_L g700 ( .A(n_459), .Y(n_700) );
INVx2_ASAP7_75t_SL g930 ( .A(n_459), .Y(n_930) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_459), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g715 ( .A(n_461), .Y(n_715) );
INVx2_ASAP7_75t_L g840 ( .A(n_461), .Y(n_840) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_461), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_468), .B1(n_469), .B2(n_481), .C(n_485), .Y(n_463) );
INVx1_ASAP7_75t_L g1370 ( .A(n_464), .Y(n_1370) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_464), .A2(n_485), .B1(n_1403), .B2(n_1414), .C(n_1415), .Y(n_1413) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g843 ( .A(n_465), .Y(n_843) );
INVx1_ASAP7_75t_L g1002 ( .A(n_465), .Y(n_1002) );
INVx1_ASAP7_75t_L g1170 ( .A(n_465), .Y(n_1170) );
INVx1_ASAP7_75t_L g1217 ( .A(n_465), .Y(n_1217) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_465), .A2(n_485), .B1(n_1477), .B2(n_1479), .C(n_1481), .Y(n_1476) );
AOI221xp5_ASAP7_75t_L g1637 ( .A1(n_465), .A2(n_1224), .B1(n_1629), .B2(n_1638), .C(n_1640), .Y(n_1637) );
INVx2_ASAP7_75t_SL g613 ( .A(n_466), .Y(n_613) );
BUFx3_ASAP7_75t_L g622 ( .A(n_466), .Y(n_622) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_466), .Y(n_787) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_466), .B(n_694), .Y(n_1224) );
BUFx4f_ASAP7_75t_L g1409 ( .A(n_466), .Y(n_1409) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_467), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_468), .A2(n_490), .B1(n_577), .B2(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g1935 ( .A(n_471), .B(n_1014), .Y(n_1935) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_472), .A2(n_488), .B1(n_605), .B2(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g682 ( .A(n_472), .Y(n_682) );
BUFx2_ASAP7_75t_L g988 ( .A(n_472), .Y(n_988) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g1891 ( .A(n_474), .B(n_1057), .Y(n_1891) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_476), .Y(n_488) );
INVx2_ASAP7_75t_L g984 ( .A(n_476), .Y(n_984) );
BUFx6f_ASAP7_75t_L g1639 ( .A(n_476), .Y(n_1639) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_479), .Y(n_1374) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g625 ( .A(n_480), .Y(n_625) );
INVx2_ASAP7_75t_L g706 ( .A(n_480), .Y(n_706) );
INVx1_ASAP7_75t_L g1457 ( .A(n_480), .Y(n_1457) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g684 ( .A(n_484), .Y(n_684) );
BUFx6f_ASAP7_75t_L g1162 ( .A(n_484), .Y(n_1162) );
INVx1_ASAP7_75t_L g1315 ( .A(n_484), .Y(n_1315) );
INVx1_ASAP7_75t_L g1549 ( .A(n_484), .Y(n_1549) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_485), .A2(n_611), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g788 ( .A(n_485), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_485), .A2(n_842), .B1(n_844), .B2(n_845), .C(n_850), .Y(n_841) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_485), .A2(n_842), .B1(n_915), .B2(n_926), .C(n_927), .Y(n_925) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_485), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_485), .A2(n_1169), .B1(n_1171), .B2(n_1172), .C(n_1176), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_485), .A2(n_1216), .B1(n_1250), .B2(n_1251), .C(n_1252), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_485), .A2(n_1216), .B1(n_1294), .B2(n_1310), .C(n_1311), .Y(n_1309) );
INVx1_ASAP7_75t_L g1377 ( .A(n_485), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1455 ( .A1(n_485), .A2(n_1169), .B1(n_1444), .B2(n_1456), .C(n_1458), .Y(n_1455) );
AOI221xp5_ASAP7_75t_L g1544 ( .A1(n_485), .A2(n_1169), .B1(n_1531), .B2(n_1545), .C(n_1547), .Y(n_1544) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g791 ( .A(n_487), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g849 ( .A(n_488), .Y(n_849) );
BUFx6f_ASAP7_75t_L g933 ( .A(n_488), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_494), .B2(n_495), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_491), .A2(n_911), .B1(n_914), .B2(n_922), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_491), .A2(n_495), .B1(n_970), .B2(n_972), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_491), .A2(n_495), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_491), .A2(n_495), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_491), .A2(n_495), .B1(n_1254), .B2(n_1255), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_491), .A2(n_495), .B1(n_1351), .B2(n_1353), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_491), .A2(n_495), .B1(n_1400), .B2(n_1402), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_491), .A2(n_495), .B1(n_1440), .B2(n_1443), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_491), .A2(n_495), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_491), .A2(n_495), .B1(n_1527), .B2(n_1529), .Y(n_1550) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_491), .A2(n_495), .B1(n_1572), .B2(n_1573), .Y(n_1571) );
AOI22xp5_ASAP7_75t_L g1641 ( .A1(n_491), .A2(n_495), .B1(n_1623), .B2(n_1628), .Y(n_1641) );
INVx6_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g600 ( .A(n_493), .Y(n_600) );
INVx1_ASAP7_75t_L g1166 ( .A(n_493), .Y(n_1166) );
BUFx2_ASAP7_75t_L g1904 ( .A(n_493), .Y(n_1904) );
AOI211xp5_ASAP7_75t_L g826 ( .A1(n_495), .A2(n_827), .B(n_828), .C(n_832), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_495), .A2(n_912), .B1(n_932), .B2(n_934), .C(n_936), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_495), .B(n_1297), .Y(n_1323) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g603 ( .A(n_497), .Y(n_603) );
INVx1_ASAP7_75t_L g935 ( .A(n_497), .Y(n_935) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g919 ( .A(n_500), .Y(n_919) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x6_ASAP7_75t_L g547 ( .A(n_501), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g634 ( .A(n_501), .Y(n_634) );
NOR3xp33_ASAP7_75t_SL g502 ( .A(n_503), .B(n_533), .C(n_546), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_520), .Y(n_503) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g877 ( .A(n_507), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_507), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_507), .Y(n_1135) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_507), .Y(n_1191) );
BUFx2_ASAP7_75t_L g1277 ( .A(n_507), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_507), .A2(n_516), .B1(n_1385), .B2(n_1386), .Y(n_1384) );
BUFx2_ASAP7_75t_L g1423 ( .A(n_507), .Y(n_1423) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
BUFx3_ASAP7_75t_L g867 ( .A(n_508), .Y(n_867) );
INVx1_ASAP7_75t_L g1271 ( .A(n_508), .Y(n_1271) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g575 ( .A(n_509), .Y(n_575) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_510), .Y(n_567) );
INVx1_ASAP7_75t_L g1099 ( .A(n_510), .Y(n_1099) );
AND2x4_ASAP7_75t_L g518 ( .A(n_511), .B(n_519), .Y(n_518) );
AND2x6_ASAP7_75t_L g516 ( .A(n_512), .B(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g522 ( .A(n_512), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g527 ( .A(n_512), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_512), .A2(n_637), .B1(n_648), .B2(n_649), .Y(n_636) );
AND2x2_ASAP7_75t_L g718 ( .A(n_512), .B(n_528), .Y(n_718) );
AND2x2_ASAP7_75t_L g723 ( .A(n_512), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g726 ( .A(n_512), .B(n_575), .Y(n_726) );
AND2x2_ASAP7_75t_L g738 ( .A(n_512), .B(n_732), .Y(n_738) );
AND2x2_ASAP7_75t_L g881 ( .A(n_512), .B(n_528), .Y(n_881) );
AND2x2_ASAP7_75t_L g950 ( .A(n_512), .B(n_528), .Y(n_950) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_512), .B(n_528), .Y(n_1428) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g585 ( .A(n_513), .Y(n_585) );
INVx2_ASAP7_75t_L g1071 ( .A(n_514), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_514), .B(n_643), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_514), .B(n_529), .Y(n_1112) );
INVx1_ASAP7_75t_L g549 ( .A(n_515), .Y(n_549) );
INVx1_ASAP7_75t_L g587 ( .A(n_515), .Y(n_587) );
INVx1_ASAP7_75t_SL g746 ( .A(n_516), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_516), .A2(n_838), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_516), .A2(n_877), .B1(n_889), .B2(n_890), .Y(n_888) );
BUFx2_ASAP7_75t_L g954 ( .A(n_516), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_516), .A2(n_1134), .B1(n_1135), .B2(n_1136), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_516), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_516), .A2(n_1245), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_516), .A2(n_1191), .B1(n_1302), .B2(n_1303), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_516), .A2(n_1422), .B1(n_1423), .B2(n_1424), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_516), .A2(n_877), .B1(n_1489), .B2(n_1490), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_516), .A2(n_1135), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_517), .B(n_540), .Y(n_545) );
BUFx2_ASAP7_75t_L g1200 ( .A(n_517), .Y(n_1200) );
BUFx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_518), .Y(n_647) );
BUFx2_ASAP7_75t_L g675 ( .A(n_518), .Y(n_675) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_518), .Y(n_732) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_518), .Y(n_1072) );
INVx1_ASAP7_75t_L g1146 ( .A(n_518), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_526), .B2(n_527), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_522), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_522), .A2(n_881), .B1(n_892), .B2(n_893), .Y(n_891) );
BUFx2_ASAP7_75t_L g948 ( .A(n_522), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_522), .A2(n_527), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_522), .A2(n_527), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_522), .A2(n_881), .B1(n_1246), .B2(n_1279), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_522), .A2(n_881), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_522), .A2(n_950), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_522), .A2(n_1426), .B1(n_1427), .B2(n_1428), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_522), .A2(n_527), .B1(n_1492), .B2(n_1493), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_522), .A2(n_1428), .B1(n_1515), .B2(n_1516), .Y(n_1514) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g724 ( .A(n_524), .Y(n_724) );
INVx2_ASAP7_75t_L g873 ( .A(n_524), .Y(n_873) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_525), .Y(n_643) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g651 ( .A(n_529), .Y(n_651) );
INVx1_ASAP7_75t_L g661 ( .A(n_529), .Y(n_661) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_529), .Y(n_730) );
BUFx2_ASAP7_75t_L g866 ( .A(n_529), .Y(n_866) );
BUFx6f_ASAP7_75t_L g1149 ( .A(n_529), .Y(n_1149) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g543 ( .A(n_530), .Y(n_543) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g895 ( .A(n_535), .Y(n_895) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2x1_ASAP7_75t_SL g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_539), .Y(n_670) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_540), .B(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g669 ( .A(n_540), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g671 ( .A(n_540), .B(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g674 ( .A(n_540), .B(n_675), .Y(n_674) );
BUFx4f_ASAP7_75t_L g751 ( .A(n_541), .Y(n_751) );
BUFx4f_ASAP7_75t_L g1299 ( .A(n_541), .Y(n_1299) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x6_ASAP7_75t_L g1086 ( .A(n_543), .B(n_1064), .Y(n_1086) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g752 ( .A(n_545), .Y(n_752) );
BUFx2_ASAP7_75t_L g896 ( .A(n_545), .Y(n_896) );
OAI33xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .A3(n_560), .B1(n_569), .B2(n_576), .B3(n_582), .Y(n_546) );
HB1xp67_ASAP7_75t_L g898 ( .A(n_547), .Y(n_898) );
OAI33xp33_ASAP7_75t_L g957 ( .A1(n_547), .A2(n_958), .A3(n_963), .B1(n_967), .B2(n_971), .B3(n_974), .Y(n_957) );
OAI33xp33_ASAP7_75t_L g1257 ( .A1(n_547), .A2(n_582), .A3(n_1258), .B1(n_1263), .B2(n_1269), .B3(n_1272), .Y(n_1257) );
OAI33xp33_ASAP7_75t_L g1284 ( .A1(n_547), .A2(n_582), .A3(n_1285), .B1(n_1288), .B2(n_1292), .B3(n_1295), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_547), .Y(n_1341) );
OAI33xp33_ASAP7_75t_L g1391 ( .A1(n_547), .A2(n_582), .A3(n_1392), .B1(n_1395), .B2(n_1398), .B3(n_1401), .Y(n_1391) );
OAI33xp33_ASAP7_75t_L g1430 ( .A1(n_547), .A2(n_582), .A3(n_1431), .B1(n_1435), .B2(n_1439), .B3(n_1442), .Y(n_1430) );
OAI33xp33_ASAP7_75t_L g1495 ( .A1(n_547), .A2(n_582), .A3(n_1496), .B1(n_1500), .B2(n_1503), .B3(n_1504), .Y(n_1495) );
OAI33xp33_ASAP7_75t_L g1606 ( .A1(n_547), .A2(n_1532), .A3(n_1607), .B1(n_1613), .B2(n_1620), .B3(n_1627), .Y(n_1606) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B1(n_554), .B2(n_559), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g760 ( .A(n_552), .Y(n_760) );
INVx1_ASAP7_75t_L g1344 ( .A(n_552), .Y(n_1344) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_554), .A2(n_900), .B1(n_1293), .B2(n_1294), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_554), .A2(n_1265), .B1(n_1481), .B2(n_1483), .Y(n_1504) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g581 ( .A(n_556), .Y(n_581) );
INVx2_ASAP7_75t_L g1109 ( .A(n_556), .Y(n_1109) );
INVx2_ASAP7_75t_L g1499 ( .A(n_556), .Y(n_1499) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_557), .B(n_558), .Y(n_737) );
INVx1_ASAP7_75t_L g673 ( .A(n_558), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B1(n_565), .B2(n_568), .Y(n_560) );
BUFx2_ASAP7_75t_L g905 ( .A(n_561), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g1914 ( .A1(n_561), .A2(n_757), .B1(n_1915), .B2(n_1916), .C(n_1917), .Y(n_1914) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1616 ( .A(n_562), .Y(n_1616) );
HB1xp67_ASAP7_75t_L g1986 ( .A(n_562), .Y(n_1986) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
BUFx2_ASAP7_75t_L g767 ( .A(n_563), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_565), .A2(n_570), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g969 ( .A(n_566), .Y(n_969) );
BUFx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_SL g639 ( .A(n_567), .Y(n_639) );
INVx2_ASAP7_75t_SL g663 ( .A(n_567), .Y(n_663) );
INVx4_ASAP7_75t_L g757 ( .A(n_567), .Y(n_757) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_567), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1151 ( .A(n_567), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_570), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g1075 ( .A(n_570), .Y(n_1075) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g638 ( .A(n_571), .Y(n_638) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_571), .Y(n_1093) );
INVx2_ASAP7_75t_L g1622 ( .A(n_571), .Y(n_1622) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g910 ( .A(n_572), .Y(n_910) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
INVx2_ASAP7_75t_L g768 ( .A(n_575), .Y(n_768) );
INVx2_ASAP7_75t_L g870 ( .A(n_575), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_577), .A2(n_1289), .B1(n_1290), .B2(n_1291), .Y(n_1288) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_579), .A2(n_581), .B1(n_606), .B2(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_579), .A2(n_581), .B1(n_665), .B2(n_666), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_579), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g901 ( .A(n_579), .Y(n_901) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_579), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1439 ( .A1(n_579), .A2(n_909), .B1(n_1440), .B2(n_1441), .Y(n_1439) );
OAI22xp33_ASAP7_75t_L g1528 ( .A1(n_579), .A2(n_1529), .B1(n_1530), .B2(n_1531), .Y(n_1528) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_580), .A2(n_900), .B1(n_902), .B2(n_903), .Y(n_899) );
OAI22xp33_ASAP7_75t_L g1272 ( .A1(n_580), .A2(n_959), .B1(n_1250), .B2(n_1254), .Y(n_1272) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_580), .A2(n_959), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
BUFx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g1268 ( .A(n_581), .Y(n_1268) );
OAI33xp33_ASAP7_75t_L g897 ( .A1(n_582), .A2(n_898), .A3(n_899), .B1(n_904), .B2(n_908), .B3(n_913), .Y(n_897) );
INVx1_ASAP7_75t_L g975 ( .A(n_582), .Y(n_975) );
CKINVDCx8_ASAP7_75t_R g582 ( .A(n_583), .Y(n_582) );
INVx5_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx6_ASAP7_75t_L g648 ( .A(n_584), .Y(n_648) );
OR2x6_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g1081 ( .A(n_586), .Y(n_1081) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OAI22x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_741), .B2(n_818), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
XNOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_676), .Y(n_592) );
XNOR2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_635), .Y(n_595) );
AOI31xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_610), .A3(n_620), .B(n_632), .Y(n_596) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g681 ( .A(n_600), .Y(n_681) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_600), .Y(n_796) );
INVx2_ASAP7_75t_L g811 ( .A(n_600), .Y(n_811) );
INVx1_ASAP7_75t_L g1934 ( .A(n_600), .Y(n_1934) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g1901 ( .A(n_602), .Y(n_1901) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g1179 ( .A(n_603), .Y(n_1179) );
INVx2_ASAP7_75t_SL g790 ( .A(n_607), .Y(n_790) );
INVx2_ASAP7_75t_SL g829 ( .A(n_607), .Y(n_829) );
INVx1_ASAP7_75t_L g992 ( .A(n_607), .Y(n_992) );
INVx1_ASAP7_75t_L g1239 ( .A(n_607), .Y(n_1239) );
AOI322xp5_ASAP7_75t_L g1312 ( .A1(n_607), .A2(n_831), .A3(n_1313), .B1(n_1316), .B2(n_1318), .C1(n_1320), .C2(n_1321), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_608), .A2(n_609), .B1(n_669), .B2(n_671), .C(n_674), .Y(n_668) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g1317 ( .A(n_613), .Y(n_1317) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_614), .Y(n_999) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g852 ( .A(n_615), .Y(n_852) );
INVxp67_ASAP7_75t_L g807 ( .A(n_617), .Y(n_807) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g628 ( .A(n_619), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_626), .B1(n_629), .B2(n_631), .Y(n_620) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_625), .A2(n_755), .B1(n_761), .B2(n_800), .C(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g997 ( .A(n_625), .Y(n_997) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_627), .Y(n_1047) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_631), .A2(n_657), .B1(n_659), .B2(n_667), .Y(n_656) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_633), .A2(n_678), .B(n_716), .C(n_727), .Y(n_677) );
NOR2xp67_ASAP7_75t_L g1061 ( .A(n_633), .B(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x4_ASAP7_75t_L g657 ( .A(n_634), .B(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g815 ( .A(n_634), .Y(n_815) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_634), .B(n_706), .Y(n_1040) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_634), .B(n_658), .Y(n_1142) );
AOI31xp33_ASAP7_75t_L g1535 ( .A1(n_634), .A2(n_1536), .A3(n_1544), .B(n_1550), .Y(n_1535) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_656), .C(n_668), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g1975 ( .A1(n_638), .A2(n_663), .B1(n_1953), .B2(n_1954), .C(n_1976), .Y(n_1975) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_639), .A2(n_1343), .B1(n_1344), .B2(n_1345), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_639), .A2(n_1074), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_644), .B2(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g1079 ( .A(n_642), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_642), .Y(n_1199) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_643), .Y(n_1144) );
INVx3_ASAP7_75t_L g1978 ( .A(n_643), .Y(n_1978) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g864 ( .A(n_646), .Y(n_864) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g728 ( .A1(n_648), .A2(n_657), .A3(n_708), .B1(n_729), .B2(n_731), .C1(n_733), .C2(n_738), .Y(n_728) );
AOI33xp33_ASAP7_75t_L g862 ( .A1(n_648), .A2(n_657), .A3(n_863), .B1(n_865), .B2(n_868), .B3(n_871), .Y(n_862) );
AOI33xp33_ASAP7_75t_L g1140 ( .A1(n_648), .A2(n_1141), .A3(n_1143), .B1(n_1147), .B2(n_1152), .B3(n_1153), .Y(n_1140) );
AOI33xp33_ASAP7_75t_L g1196 ( .A1(n_648), .A2(n_1197), .A3(n_1198), .B1(n_1201), .B2(n_1202), .B3(n_1204), .Y(n_1196) );
INVx1_ASAP7_75t_L g1532 ( .A(n_648), .Y(n_1532) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g1203 ( .A(n_653), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_657), .Y(n_1197) );
INVx1_ASAP7_75t_L g1107 ( .A(n_658), .Y(n_1107) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_663), .A2(n_773), .B1(n_1520), .B2(n_1521), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_667), .A2(n_671), .B1(n_687), .B2(n_720), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_669), .A2(n_674), .B(n_740), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_669), .A2(n_671), .B1(n_674), .B2(n_860), .C(n_861), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_669), .A2(n_1128), .B1(n_1130), .B2(n_1131), .C(n_1132), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g1186 ( .A1(n_669), .A2(n_671), .B1(n_674), .B2(n_1187), .C(n_1188), .Y(n_1186) );
AOI221xp5_ASAP7_75t_L g1590 ( .A1(n_669), .A2(n_671), .B1(n_674), .B2(n_1591), .C(n_1592), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_670), .B(n_1063), .Y(n_1084) );
INVx1_ASAP7_75t_L g1129 ( .A(n_671), .Y(n_1129) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_674), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1587 ( .A(n_675), .Y(n_1587) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_686), .C(n_695), .D(n_707), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_684), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
INVx1_ASAP7_75t_L g853 ( .A(n_684), .Y(n_853) );
INVx1_ASAP7_75t_L g1000 ( .A(n_684), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1363 ( .A1(n_684), .A2(n_1050), .B1(n_1336), .B2(n_1364), .C(n_1365), .Y(n_1363) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B(n_690), .C(n_693), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx4_ASAP7_75t_L g779 ( .A(n_689), .Y(n_779) );
INVx2_ASAP7_75t_L g986 ( .A(n_689), .Y(n_986) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .C(n_701), .Y(n_695) );
BUFx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g710 ( .A(n_698), .Y(n_710) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_698), .B(n_1014), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_700), .Y(n_1044) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g1026 ( .A(n_703), .Y(n_1026) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B(n_711), .C(n_713), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g1903 ( .A1(n_709), .A2(n_1904), .B1(n_1905), .B2(n_1906), .C(n_1907), .Y(n_1903) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g785 ( .A(n_712), .Y(n_785) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_712), .Y(n_1042) );
INVx1_ASAP7_75t_L g813 ( .A(n_715), .Y(n_813) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g745 ( .A(n_718), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g1602 ( .A1(n_718), .A2(n_723), .B1(n_1603), .B2(n_1604), .Y(n_1602) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_725), .B2(n_726), .Y(n_721) );
INVx1_ASAP7_75t_L g775 ( .A(n_723), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_724), .B(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g748 ( .A(n_726), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1599 ( .A1(n_726), .A2(n_738), .B1(n_1600), .B2(n_1601), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_739), .Y(n_727) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_732), .Y(n_874) );
BUFx3_ASAP7_75t_L g762 ( .A(n_736), .Y(n_762) );
INVx2_ASAP7_75t_L g774 ( .A(n_736), .Y(n_774) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g818 ( .A(n_741), .Y(n_818) );
INVx1_ASAP7_75t_L g816 ( .A(n_742), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_749), .C(n_776), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_751), .Y(n_956) );
HB1xp67_ASAP7_75t_L g1339 ( .A(n_751), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_756), .A2(n_759), .B1(n_795), .B2(n_797), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_757), .A2(n_905), .B1(n_906), .B2(n_907), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_757), .A2(n_909), .B1(n_911), .B2(n_912), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_757), .A2(n_1260), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
INVx2_ASAP7_75t_L g1584 ( .A(n_757), .Y(n_1584) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_762), .A2(n_959), .B1(n_961), .B2(n_962), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_762), .A2(n_959), .B1(n_972), .B2(n_973), .Y(n_971) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_762), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_768), .B2(n_769), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_764), .A2(n_772), .B1(n_784), .B2(n_786), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_765), .A2(n_1436), .B1(n_1437), .B2(n_1438), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1924 ( .A1(n_765), .A2(n_1437), .B1(n_1925), .B2(n_1926), .Y(n_1924) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1285 ( .A1(n_768), .A2(n_905), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_768), .A2(n_1260), .B1(n_1399), .B2(n_1400), .Y(n_1398) );
INVx2_ASAP7_75t_L g1619 ( .A(n_768), .Y(n_1619) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_769), .A2(n_771), .B1(n_779), .B2(n_780), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_773), .A2(n_900), .B1(n_914), .B2(n_915), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_773), .A2(n_1074), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
OAI22xp5_ASAP7_75t_SL g1627 ( .A1(n_773), .A2(n_1103), .B1(n_1628), .B2(n_1629), .Y(n_1627) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g1291 ( .A(n_774), .Y(n_1291) );
OAI31xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_789), .A3(n_793), .B(n_814), .Y(n_776) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OR2x6_ASAP7_75t_L g1013 ( .A(n_782), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_787), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_787), .B(n_1057), .Y(n_1056) );
OR2x6_ASAP7_75t_L g1037 ( .A(n_792), .B(n_1034), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1911 ( .A(n_792), .B(n_1034), .Y(n_1911) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_799), .B1(n_805), .B2(n_809), .Y(n_793) );
OAI21xp5_ASAP7_75t_SL g1564 ( .A1(n_795), .A2(n_1565), .B(n_1566), .Y(n_1564) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI221xp5_ASAP7_75t_L g809 ( .A1(n_800), .A2(n_810), .B1(n_811), .B2(n_812), .C(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g1542 ( .A(n_800), .Y(n_1542) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g1898 ( .A(n_801), .Y(n_1898) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_SL g847 ( .A(n_804), .Y(n_847) );
INVx2_ASAP7_75t_L g1242 ( .A(n_804), .Y(n_1242) );
OAI221xp5_ASAP7_75t_L g1895 ( .A1(n_811), .A2(n_1896), .B1(n_1897), .B2(n_1899), .C(n_1900), .Y(n_1895) );
INVx2_ASAP7_75t_L g1460 ( .A(n_814), .Y(n_1460) );
AOI22xp5_ASAP7_75t_L g1630 ( .A1(n_814), .A2(n_1631), .B1(n_1642), .B2(n_1643), .Y(n_1630) );
CKINVDCx8_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
AOI31xp33_ASAP7_75t_L g1157 ( .A1(n_815), .A2(n_1158), .A3(n_1168), .B(n_1180), .Y(n_1157) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_941), .B1(n_1115), .B2(n_1116), .Y(n_820) );
INVx1_ASAP7_75t_L g1115 ( .A(n_821), .Y(n_1115) );
XOR2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_883), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_882), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_858), .Y(n_823) );
NAND3xp33_ASAP7_75t_SL g825 ( .A(n_826), .B(n_841), .C(n_854), .Y(n_825) );
INVx2_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g1220 ( .A(n_834), .Y(n_1220) );
OAI21xp5_ASAP7_75t_SL g835 ( .A1(n_836), .A2(n_838), .B(n_839), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1454 ( .A(n_837), .Y(n_1454) );
INVx1_ASAP7_75t_L g1167 ( .A(n_840), .Y(n_1167) );
BUFx2_ASAP7_75t_L g1319 ( .A(n_840), .Y(n_1319) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1478 ( .A(n_849), .Y(n_1478) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
AND4x1_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .C(n_875), .D(n_878), .Y(n_858) );
HB1xp67_ASAP7_75t_L g1586 ( .A(n_866), .Y(n_1586) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_867), .Y(n_966) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
BUFx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
XNOR2x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_916), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_894), .C(n_897), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .Y(n_887) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_909), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_909), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_967) );
BUFx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g1261 ( .A(n_910), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_920), .B1(n_939), .B2(n_940), .Y(n_916) );
INVx1_ASAP7_75t_SL g1005 ( .A(n_917), .Y(n_1005) );
INVx5_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
AOI31xp33_ASAP7_75t_L g1235 ( .A1(n_918), .A2(n_1236), .A3(n_1249), .B(n_1253), .Y(n_1235) );
AOI31xp33_ASAP7_75t_L g1359 ( .A1(n_918), .A2(n_1360), .A3(n_1368), .B(n_1378), .Y(n_1359) );
AOI31xp33_ASAP7_75t_L g1406 ( .A1(n_918), .A2(n_1407), .A3(n_1413), .B(n_1416), .Y(n_1406) );
OAI31xp33_ASAP7_75t_L g1973 ( .A1(n_918), .A2(n_1974), .A3(n_1980), .B(n_1989), .Y(n_1973) );
BUFx8_ASAP7_75t_SL g918 ( .A(n_919), .Y(n_918) );
OAI31xp33_ASAP7_75t_L g1066 ( .A1(n_919), .A2(n_1067), .A3(n_1087), .B(n_1110), .Y(n_1066) );
INVx2_ASAP7_75t_L g1206 ( .A(n_919), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_925), .C(n_931), .Y(n_920) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g1632 ( .A1(n_924), .A2(n_1621), .B1(n_1633), .B2(n_1634), .C(n_1635), .Y(n_1632) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_933), .Y(n_996) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_938), .Y(n_1211) );
AOI21xp5_ASAP7_75t_L g976 ( .A1(n_940), .A2(n_977), .B(n_978), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g1557 ( .A1(n_940), .A2(n_1558), .B(n_1559), .Y(n_1557) );
INVx1_ASAP7_75t_L g1116 ( .A(n_941), .Y(n_1116) );
XOR2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_1006), .Y(n_941) );
XNOR2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
OAI22xp5_ASAP7_75t_SL g1698 ( .A1(n_943), .A2(n_1686), .B1(n_1699), .B2(n_1700), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_976), .Y(n_944) );
NOR3xp33_ASAP7_75t_SL g945 ( .A(n_946), .B(n_955), .C(n_957), .Y(n_945) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_948), .A2(n_1335), .B1(n_1336), .B2(n_1337), .Y(n_1334) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVxp67_ASAP7_75t_SL g1333 ( .A(n_954), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_954), .A2(n_1423), .B1(n_1577), .B2(n_1578), .Y(n_1576) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_959), .A2(n_1432), .B1(n_1433), .B2(n_1434), .Y(n_1431) );
OAI22xp33_ASAP7_75t_SL g1522 ( .A1(n_959), .A2(n_1074), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
OAI221xp5_ASAP7_75t_L g1923 ( .A1(n_959), .A2(n_1106), .B1(n_1291), .B2(n_1896), .C(n_1899), .Y(n_1923) );
INVx3_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_966), .A2(n_1259), .B1(n_1260), .B2(n_1262), .Y(n_1258) );
OAI22xp33_ASAP7_75t_L g1442 ( .A1(n_966), .A2(n_1433), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_966), .A2(n_1270), .B1(n_1474), .B2(n_1484), .Y(n_1503) );
AOI221xp5_ASAP7_75t_SL g979 ( .A1(n_968), .A2(n_980), .B1(n_987), .B2(n_989), .C(n_991), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_973), .A2(n_994), .B1(n_998), .B2(n_1001), .C(n_1003), .Y(n_993) );
OAI33xp33_ASAP7_75t_L g1340 ( .A1(n_974), .A2(n_1341), .A3(n_1342), .B1(n_1346), .B2(n_1349), .B3(n_1352), .Y(n_1340) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AOI33xp33_ASAP7_75t_L g1580 ( .A1(n_975), .A2(n_1581), .A3(n_1583), .B1(n_1585), .B2(n_1588), .B3(n_1589), .Y(n_1580) );
AOI31xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_993), .A3(n_1004), .B(n_1005), .Y(n_978) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx3_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx2_ASAP7_75t_L g1175 ( .A(n_984), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g1536 ( .A1(n_989), .A2(n_1526), .B(n_1537), .Y(n_1536) );
AOI211xp5_ASAP7_75t_SL g1560 ( .A1(n_989), .A2(n_1561), .B(n_1562), .C(n_1563), .Y(n_1560) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1567 ( .A1(n_1001), .A2(n_1003), .B1(n_1568), .B2(n_1569), .C(n_1570), .Y(n_1567) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_1002), .Y(n_1001) );
AOI31xp33_ASAP7_75t_L g1559 ( .A1(n_1005), .A2(n_1560), .A3(n_1567), .B(n_1571), .Y(n_1559) );
OAI31xp33_ASAP7_75t_L g1912 ( .A1(n_1005), .A2(n_1913), .A3(n_1922), .B(n_1927), .Y(n_1912) );
AND3x1_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1058), .C(n_1066), .Y(n_1007) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1027), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1018), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1012), .B1(n_1015), .B2(n_1016), .Y(n_1010) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_1011), .A2(n_1024), .B1(n_1074), .B2(n_1076), .C(n_1077), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1952 ( .A1(n_1012), .A2(n_1025), .B1(n_1953), .B2(n_1954), .Y(n_1952) );
CKINVDCx6p67_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1014), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1933 ( .A(n_1014), .B(n_1934), .Y(n_1933) );
AOI22xp33_ASAP7_75t_L g1955 ( .A1(n_1016), .A2(n_1020), .B1(n_1956), .B2(n_1957), .Y(n_1955) );
CKINVDCx6p67_ASAP7_75t_R g1016 ( .A(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1020), .B1(n_1024), .B2(n_1025), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1023), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_1021), .Y(n_1177) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1022), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1023), .B(n_1026), .Y(n_1025) );
NAND3xp33_ASAP7_75t_SL g1027 ( .A(n_1028), .B(n_1038), .C(n_1054), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1030), .B1(n_1035), .B2(n_1036), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_1029), .A2(n_1035), .B1(n_1083), .B2(n_1085), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1959 ( .A1(n_1030), .A2(n_1036), .B1(n_1960), .B2(n_1961), .Y(n_1959) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx2_ASAP7_75t_L g1910 ( .A(n_1031), .Y(n_1910) );
NAND2x1p5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1034), .Y(n_1057) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AOI33xp33_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1041), .A3(n_1043), .B1(n_1046), .B2(n_1048), .B3(n_1052), .Y(n_1038) );
CKINVDCx5p33_ASAP7_75t_R g1039 ( .A(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1894 ( .A(n_1040), .Y(n_1894) );
CKINVDCx5p33_ASAP7_75t_R g1963 ( .A(n_1040), .Y(n_1963) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1050), .Y(n_1411) );
BUFx4f_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx4_ASAP7_75t_L g1902 ( .A(n_1053), .Y(n_1902) );
AOI33xp33_ASAP7_75t_L g1962 ( .A1(n_1053), .A2(n_1963), .A3(n_1964), .B1(n_1965), .B2(n_1966), .B3(n_1967), .Y(n_1962) );
NAND3xp33_ASAP7_75t_SL g1958 ( .A(n_1054), .B(n_1959), .C(n_1962), .Y(n_1958) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1887 ( .A(n_1060), .B(n_1888), .Y(n_1887) );
NAND2xp5_ASAP7_75t_L g1971 ( .A(n_1060), .B(n_1972), .Y(n_1971) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1064), .B(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx8_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
AND2x4_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1072), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1114 ( .A(n_1070), .B(n_1098), .Y(n_1114) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
OAI22xp5_ASAP7_75t_SL g1500 ( .A1(n_1076), .A2(n_1270), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_1076), .A2(n_1092), .B1(n_1526), .B2(n_1527), .Y(n_1525) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1918 ( .A(n_1081), .Y(n_1918) );
AOI22xp33_ASAP7_75t_L g1919 ( .A1(n_1083), .A2(n_1085), .B1(n_1920), .B2(n_1921), .Y(n_1919) );
AOI22xp33_ASAP7_75t_L g1979 ( .A1(n_1083), .A2(n_1085), .B1(n_1960), .B2(n_1961), .Y(n_1979) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
CKINVDCx11_ASAP7_75t_R g1085 ( .A(n_1086), .Y(n_1085) );
CKINVDCx6p67_ASAP7_75t_R g1088 ( .A(n_1089), .Y(n_1088) );
OAI22xp5_ASAP7_75t_SL g1090 ( .A1(n_1091), .A2(n_1092), .B1(n_1094), .B2(n_1095), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1984 ( .A1(n_1095), .A2(n_1985), .B1(n_1987), .B2(n_1988), .Y(n_1984) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1099), .Y(n_1626) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1103), .B2(n_1105), .C(n_1106), .Y(n_1100) );
OAI22xp33_ASAP7_75t_L g1352 ( .A1(n_1101), .A2(n_1344), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
OAI221xp5_ASAP7_75t_L g1981 ( .A1(n_1101), .A2(n_1103), .B1(n_1106), .B2(n_1982), .C(n_1983), .Y(n_1981) );
OAI22xp33_ASAP7_75t_L g1395 ( .A1(n_1103), .A2(n_1291), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_1109), .Y(n_1530) );
INVx3_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx3_ASAP7_75t_L g1928 ( .A(n_1112), .Y(n_1928) );
INVx3_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx3_ASAP7_75t_L g1929 ( .A(n_1114), .Y(n_1929) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
XNOR2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1464), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1121), .B1(n_1326), .B2(n_1463), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
AO22x2_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1123), .B1(n_1229), .B2(n_1230), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
XNOR2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1183), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1154), .Y(n_1125) );
AND4x1_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1133), .C(n_1137), .D(n_1140), .Y(n_1126) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1337 ( .A(n_1135), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_1136), .A2(n_1138), .B1(n_1164), .B2(n_1165), .C(n_1167), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_L g1582 ( .A(n_1142), .Y(n_1582) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
AOI21xp33_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1156), .B(n_1157), .Y(n_1154) );
AOI21xp5_ASAP7_75t_L g1445 ( .A1(n_1155), .A2(n_1446), .B(n_1447), .Y(n_1445) );
AOI21xp5_ASAP7_75t_L g1533 ( .A1(n_1155), .A2(n_1534), .B(n_1535), .Y(n_1533) );
OAI221xp5_ASAP7_75t_L g1243 ( .A1(n_1165), .A2(n_1244), .B1(n_1245), .B2(n_1246), .C(n_1247), .Y(n_1243) );
OAI221xp5_ASAP7_75t_L g1453 ( .A1(n_1165), .A2(n_1167), .B1(n_1424), .B2(n_1426), .C(n_1454), .Y(n_1453) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1174), .Y(n_1373) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1205), .Y(n_1184) );
AND4x1_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1189), .C(n_1193), .D(n_1196), .Y(n_1185) );
INVx2_ASAP7_75t_SL g1437 ( .A(n_1203), .Y(n_1437) );
NAND3xp33_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1215), .C(n_1225), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1218), .B1(n_1219), .B2(n_1221), .C(n_1224), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
XOR2xp5_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1280), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1256), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_1237), .A2(n_1255), .B1(n_1270), .B2(n_1271), .Y(n_1269) );
INVx2_ASAP7_75t_SL g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1248), .Y(n_1367) );
NOR3xp33_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1273), .C(n_1274), .Y(n_1256) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1261), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B1(n_1266), .B2(n_1267), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1496 ( .A1(n_1265), .A2(n_1497), .B1(n_1498), .B2(n_1499), .Y(n_1496) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1268), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1307), .Y(n_1282) );
NOR3xp33_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1298), .C(n_1300), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1304), .Y(n_1300) );
NAND4xp25_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1312), .C(n_1322), .D(n_1323), .Y(n_1308) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1326), .Y(n_1463) );
XNOR2x1_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1379), .Y(n_1326) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
XNOR2x1_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1355), .Y(n_1330) );
NOR3xp33_ASAP7_75t_SL g1331 ( .A(n_1332), .B(n_1338), .C(n_1340), .Y(n_1331) );
OAI33xp33_ASAP7_75t_L g1518 ( .A1(n_1341), .A2(n_1519), .A3(n_1522), .B1(n_1525), .B2(n_1528), .B3(n_1532), .Y(n_1518) );
AOI21xp5_ASAP7_75t_L g1360 ( .A1(n_1350), .A2(n_1361), .B(n_1362), .Y(n_1360) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_1354), .A2(n_1369), .B1(n_1371), .B2(n_1375), .C(n_1376), .Y(n_1368) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1358), .B(n_1359), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
XOR2x2_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1417), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1404), .Y(n_1381) );
NOR3xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1390), .C(n_1391), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1387), .Y(n_1383) );
BUFx2_ASAP7_75t_L g1546 ( .A(n_1409), .Y(n_1546) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1418), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1445), .Y(n_1418) );
NOR3xp33_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1429), .C(n_1430), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1421), .B(n_1425), .Y(n_1420) );
AOI31xp33_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1455), .A3(n_1459), .B(n_1460), .Y(n_1447) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
AOI22xp33_ASAP7_75t_SL g1464 ( .A1(n_1465), .A2(n_1466), .B1(n_1553), .B2(n_1645), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
AO22x2_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1506), .B1(n_1551), .B2(n_1552), .Y(n_1466) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1467), .Y(n_1552) );
XOR2x2_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1505), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1486), .Y(n_1468) );
NAND3xp33_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1476), .C(n_1482), .Y(n_1470) );
NOR3xp33_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1494), .C(n_1495), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1491), .Y(n_1487) );
OAI22xp33_ASAP7_75t_L g1607 ( .A1(n_1499), .A2(n_1608), .B1(n_1609), .B2(n_1612), .Y(n_1607) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1506), .Y(n_1551) );
XNOR2xp5_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1508), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1533), .Y(n_1508) );
NOR3xp33_ASAP7_75t_SL g1509 ( .A(n_1510), .B(n_1517), .C(n_1518), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1514), .Y(n_1510) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
AOI31xp33_ASAP7_75t_L g1538 ( .A1(n_1539), .A2(n_1540), .A3(n_1541), .B(n_1543), .Y(n_1538) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1553), .Y(n_1645) );
AOI22xp5_ASAP7_75t_L g1553 ( .A1(n_1554), .A2(n_1593), .B1(n_1594), .B2(n_1644), .Y(n_1553) );
INVx2_ASAP7_75t_SL g1644 ( .A(n_1554), .Y(n_1644) );
XNOR2x1_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1556), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1574), .Y(n_1556) );
NOR2xp33_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1579), .Y(n_1574) );
NAND2xp5_ASAP7_75t_SL g1579 ( .A(n_1580), .B(n_1590), .Y(n_1579) );
INVx2_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
XNOR2x1_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1596), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1630), .Y(n_1596) );
NOR3xp33_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1605), .C(n_1606), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1602), .Y(n_1598) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1611), .Y(n_1610) );
OAI22xp5_ASAP7_75t_L g1613 ( .A1(n_1614), .A2(n_1615), .B1(n_1617), .B2(n_1618), .Y(n_1613) );
BUFx2_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
OAI22xp5_ASAP7_75t_SL g1620 ( .A1(n_1621), .A2(n_1622), .B1(n_1623), .B2(n_1624), .Y(n_1620) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
NAND3xp33_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1637), .C(n_1641), .Y(n_1631) );
OAI221xp5_ASAP7_75t_L g1646 ( .A1(n_1647), .A2(n_1879), .B1(n_1881), .B2(n_1936), .C(n_1941), .Y(n_1646) );
HB1xp67_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NOR4xp25_ASAP7_75t_L g1648 ( .A(n_1649), .B(n_1743), .C(n_1829), .D(n_1856), .Y(n_1648) );
O2A1O1Ixp33_ASAP7_75t_L g1649 ( .A1(n_1650), .A2(n_1680), .B(n_1701), .C(n_1735), .Y(n_1649) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
OAI211xp5_ASAP7_75t_L g1827 ( .A1(n_1651), .A2(n_1722), .B(n_1759), .C(n_1828), .Y(n_1827) );
AOI21xp5_ASAP7_75t_L g1854 ( .A1(n_1651), .A2(n_1707), .B(n_1774), .Y(n_1854) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_1651), .B(n_1860), .Y(n_1859) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1671), .Y(n_1651) );
CKINVDCx5p33_ASAP7_75t_R g1708 ( .A(n_1652), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1652), .B(n_1677), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1652), .B(n_1711), .Y(n_1788) );
NOR2xp33_ASAP7_75t_L g1798 ( .A(n_1652), .B(n_1799), .Y(n_1798) );
OR2x2_ASAP7_75t_L g1802 ( .A(n_1652), .B(n_1803), .Y(n_1802) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1652), .B(n_1799), .Y(n_1815) );
NOR2xp33_ASAP7_75t_L g1825 ( .A(n_1652), .B(n_1761), .Y(n_1825) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_1652), .B(n_1739), .Y(n_1831) );
AND2x2_ASAP7_75t_L g1837 ( .A(n_1652), .B(n_1771), .Y(n_1837) );
AND2x2_ASAP7_75t_L g1867 ( .A(n_1652), .B(n_1762), .Y(n_1867) );
AND2x4_ASAP7_75t_SL g1652 ( .A(n_1653), .B(n_1665), .Y(n_1652) );
AND2x4_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1660), .Y(n_1654) );
OAI21xp33_ASAP7_75t_SL g1991 ( .A1(n_1655), .A2(n_1945), .B(n_1992), .Y(n_1991) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1691 ( .A(n_1656), .B(n_1661), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1659), .Y(n_1656) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1659), .Y(n_1669) );
AND2x4_ASAP7_75t_L g1662 ( .A(n_1660), .B(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1661), .B(n_1664), .Y(n_1695) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1668), .Y(n_1666) );
AND2x4_ASAP7_75t_L g1670 ( .A(n_1667), .B(n_1669), .Y(n_1670) );
AND2x4_ASAP7_75t_L g1684 ( .A(n_1667), .B(n_1668), .Y(n_1684) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx2_ASAP7_75t_L g1686 ( .A(n_1670), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1671), .B(n_1708), .Y(n_1732) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1671), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1812 ( .A(n_1671), .B(n_1788), .Y(n_1812) );
AOI22xp33_ASAP7_75t_L g1877 ( .A1(n_1671), .A2(n_1736), .B1(n_1795), .B2(n_1878), .Y(n_1877) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1676), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1672), .B(n_1677), .Y(n_1739) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1672), .Y(n_1799) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1673), .B(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1673), .B(n_1677), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1675), .Y(n_1673) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
INVxp67_ASAP7_75t_SL g1720 ( .A(n_1677), .Y(n_1720) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1677), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1679), .Y(n_1677) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1680), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1696), .Y(n_1680) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1681), .Y(n_1746) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
BUFx3_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1684), .Y(n_1699) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx2_ASAP7_75t_L g1713 ( .A(n_1686), .Y(n_1713) );
OAI22xp33_ASAP7_75t_L g1687 ( .A1(n_1688), .A2(n_1689), .B1(n_1692), .B2(n_1693), .Y(n_1687) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1689), .Y(n_1880) );
BUFx3_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
OAI22xp33_ASAP7_75t_L g1714 ( .A1(n_1690), .A2(n_1715), .B1(n_1716), .B2(n_1717), .Y(n_1714) );
BUFx6f_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
HB1xp67_ASAP7_75t_L g1717 ( .A(n_1695), .Y(n_1717) );
CKINVDCx6p67_ASAP7_75t_R g1755 ( .A(n_1696), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1696), .B(n_1765), .Y(n_1769) );
OR2x2_ASAP7_75t_L g1796 ( .A(n_1696), .B(n_1765), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1696), .B(n_1725), .Y(n_1819) );
OR2x2_ASAP7_75t_L g1826 ( .A(n_1696), .B(n_1740), .Y(n_1826) );
OR2x6_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1698), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1759 ( .A(n_1697), .B(n_1698), .Y(n_1759) );
OAI22xp5_ASAP7_75t_L g1701 ( .A1(n_1702), .A2(n_1721), .B1(n_1728), .B2(n_1733), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1707), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_1703), .B(n_1711), .Y(n_1804) );
A2O1A1Ixp33_ASAP7_75t_L g1851 ( .A1(n_1703), .A2(n_1765), .B(n_1852), .C(n_1854), .Y(n_1851) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1704), .Y(n_1723) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1704), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1704), .B(n_1724), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1704), .B(n_1725), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1704), .B(n_1755), .Y(n_1754) );
OAI321xp33_ASAP7_75t_L g1790 ( .A1(n_1704), .A2(n_1744), .A3(n_1791), .B1(n_1793), .B2(n_1794), .C(n_1800), .Y(n_1790) );
NAND3xp33_ASAP7_75t_L g1811 ( .A(n_1704), .B(n_1795), .C(n_1812), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1706), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1709), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1737 ( .A(n_1708), .B(n_1738), .Y(n_1737) );
OR2x2_ASAP7_75t_L g1749 ( .A(n_1708), .B(n_1750), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1708), .B(n_1712), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1708), .B(n_1719), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1822 ( .A(n_1708), .B(n_1739), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1845 ( .A(n_1708), .B(n_1771), .Y(n_1845) );
AND2x2_ASAP7_75t_L g1853 ( .A(n_1708), .B(n_1752), .Y(n_1853) );
NOR2xp33_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1718), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1710), .B(n_1739), .Y(n_1738) );
NOR2x1p5_ASAP7_75t_L g1752 ( .A(n_1710), .B(n_1753), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1710), .B(n_1798), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1710), .B(n_1722), .Y(n_1816) );
HB1xp67_ASAP7_75t_L g1860 ( .A(n_1710), .Y(n_1860) );
INVx2_ASAP7_75t_SL g1710 ( .A(n_1711), .Y(n_1710) );
BUFx3_ASAP7_75t_L g1731 ( .A(n_1711), .Y(n_1731) );
BUFx2_ASAP7_75t_L g1751 ( .A(n_1711), .Y(n_1751) );
NOR2xp33_ASAP7_75t_L g1874 ( .A(n_1711), .B(n_1723), .Y(n_1874) );
INVx2_ASAP7_75t_SL g1711 ( .A(n_1712), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1712), .B(n_1723), .Y(n_1774) );
OR2x2_ASAP7_75t_L g1750 ( .A(n_1718), .B(n_1751), .Y(n_1750) );
NOR2xp33_ASAP7_75t_L g1861 ( .A(n_1718), .B(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1719), .B(n_1780), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_1719), .B(n_1788), .Y(n_1810) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
NAND2xp5_ASAP7_75t_SL g1870 ( .A(n_1722), .B(n_1755), .Y(n_1870) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1724), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1723), .B(n_1755), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1789 ( .A(n_1723), .B(n_1725), .Y(n_1789) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
BUFx6f_ASAP7_75t_L g1734 ( .A(n_1725), .Y(n_1734) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1725), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
INVxp67_ASAP7_75t_L g1833 ( .A(n_1728), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
INVx3_ASAP7_75t_L g1809 ( .A(n_1729), .Y(n_1809) );
AOI221xp5_ASAP7_75t_L g1842 ( .A1(n_1729), .A2(n_1744), .B1(n_1789), .B2(n_1843), .C(n_1846), .Y(n_1842) );
O2A1O1Ixp33_ASAP7_75t_L g1817 ( .A1(n_1730), .A2(n_1818), .B(n_1819), .C(n_1820), .Y(n_1817) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1732), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1847 ( .A(n_1731), .B(n_1845), .Y(n_1847) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1731), .Y(n_1869) );
A2O1A1Ixp33_ASAP7_75t_L g1848 ( .A1(n_1733), .A2(n_1797), .B(n_1849), .C(n_1851), .Y(n_1848) );
CKINVDCx14_ASAP7_75t_R g1733 ( .A(n_1734), .Y(n_1733) );
AOI32xp33_ASAP7_75t_L g1838 ( .A1(n_1734), .A2(n_1738), .A3(n_1744), .B1(n_1839), .B2(n_1840), .Y(n_1838) );
OAI21xp5_ASAP7_75t_L g1735 ( .A1(n_1736), .A2(n_1740), .B(n_1741), .Y(n_1735) );
INVx2_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
INVx2_ASAP7_75t_L g1753 ( .A(n_1739), .Y(n_1753) );
INVx2_ASAP7_75t_L g1832 ( .A(n_1740), .Y(n_1832) );
AOI21xp33_ASAP7_75t_L g1875 ( .A1(n_1741), .A2(n_1778), .B(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1742), .B(n_1751), .Y(n_1758) );
AOI21xp33_ASAP7_75t_L g1834 ( .A1(n_1742), .A2(n_1835), .B(n_1838), .Y(n_1834) );
OAI211xp5_ASAP7_75t_L g1743 ( .A1(n_1744), .A2(n_1747), .B(n_1776), .C(n_1817), .Y(n_1743) );
INVx3_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AOI31xp33_ASAP7_75t_L g1856 ( .A1(n_1745), .A2(n_1857), .A3(n_1863), .B(n_1877), .Y(n_1856) );
INVx2_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g1793 ( .A(n_1746), .B(n_1755), .Y(n_1793) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1746), .B(n_1765), .Y(n_1841) );
O2A1O1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1748), .A2(n_1752), .B(n_1754), .C(n_1756), .Y(n_1747) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
NAND2xp5_ASAP7_75t_L g1843 ( .A(n_1750), .B(n_1844), .Y(n_1843) );
OR2x2_ASAP7_75t_L g1766 ( .A(n_1751), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1751), .B(n_1771), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1824 ( .A(n_1751), .B(n_1825), .Y(n_1824) );
INVx2_ASAP7_75t_L g1828 ( .A(n_1751), .Y(n_1828) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1752), .Y(n_1871) );
AOI221xp5_ASAP7_75t_L g1777 ( .A1(n_1754), .A2(n_1778), .B1(n_1781), .B2(n_1782), .C(n_1784), .Y(n_1777) );
CKINVDCx5p33_ASAP7_75t_R g1868 ( .A(n_1754), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1764 ( .A(n_1755), .B(n_1765), .Y(n_1764) );
AOI31xp33_ASAP7_75t_L g1784 ( .A1(n_1755), .A2(n_1785), .A3(n_1788), .B(n_1789), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1864 ( .A(n_1755), .B(n_1789), .Y(n_1864) );
OAI321xp33_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1759), .A3(n_1760), .B1(n_1763), .B2(n_1766), .C(n_1768), .Y(n_1756) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
NOR3xp33_ASAP7_75t_L g1772 ( .A(n_1759), .B(n_1773), .C(n_1775), .Y(n_1772) );
OAI211xp5_ASAP7_75t_L g1813 ( .A1(n_1759), .A2(n_1814), .B(n_1815), .C(n_1816), .Y(n_1813) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
OAI221xp5_ASAP7_75t_SL g1820 ( .A1(n_1763), .A2(n_1782), .B1(n_1821), .B2(n_1826), .C(n_1827), .Y(n_1820) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1767), .Y(n_1873) );
AOI21xp5_ASAP7_75t_L g1768 ( .A1(n_1769), .A2(n_1770), .B(n_1772), .Y(n_1768) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1769), .Y(n_1807) );
AOI211xp5_ASAP7_75t_L g1863 ( .A1(n_1770), .A2(n_1864), .B(n_1865), .C(n_1875), .Y(n_1863) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1771), .Y(n_1775) );
OAI211xp5_ASAP7_75t_L g1800 ( .A1(n_1771), .A2(n_1801), .B(n_1804), .C(n_1805), .Y(n_1800) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
OR2x2_ASAP7_75t_L g1782 ( .A(n_1775), .B(n_1783), .Y(n_1782) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1775), .B(n_1787), .Y(n_1786) );
NOR3xp33_ASAP7_75t_SL g1776 ( .A(n_1777), .B(n_1790), .C(n_1806), .Y(n_1776) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1818 ( .A(n_1779), .B(n_1809), .Y(n_1818) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1780), .Y(n_1783) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
AOI21xp5_ASAP7_75t_L g1857 ( .A1(n_1789), .A2(n_1858), .B(n_1861), .Y(n_1857) );
NAND2xp5_ASAP7_75t_L g1835 ( .A(n_1791), .B(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1793), .Y(n_1855) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1795), .B(n_1797), .Y(n_1794) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
HB1xp67_ASAP7_75t_L g1814 ( .A(n_1798), .Y(n_1814) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1799), .Y(n_1803) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
OAI211xp5_ASAP7_75t_L g1806 ( .A1(n_1807), .A2(n_1808), .B(n_1811), .C(n_1813), .Y(n_1806) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1809), .B(n_1810), .Y(n_1808) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1809), .Y(n_1850) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1812), .Y(n_1876) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1816), .Y(n_1862) );
AOI21xp5_ASAP7_75t_L g1830 ( .A1(n_1818), .A2(n_1831), .B(n_1832), .Y(n_1830) );
NOR2xp33_ASAP7_75t_L g1821 ( .A(n_1822), .B(n_1823), .Y(n_1821) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1822), .Y(n_1839) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1826), .Y(n_1878) );
AOI321xp33_ASAP7_75t_L g1829 ( .A1(n_1830), .A2(n_1833), .A3(n_1834), .B1(n_1842), .B2(n_1848), .C(n_1855), .Y(n_1829) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1849 ( .A(n_1850), .Y(n_1849) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
OAI321xp33_ASAP7_75t_L g1865 ( .A1(n_1866), .A2(n_1868), .A3(n_1869), .B1(n_1870), .B2(n_1871), .C(n_1872), .Y(n_1865) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
NAND2xp5_ASAP7_75t_L g1872 ( .A(n_1873), .B(n_1874), .Y(n_1872) );
CKINVDCx16_ASAP7_75t_R g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1883), .Y(n_1882) );
INVx1_ASAP7_75t_L g1883 ( .A(n_1884), .Y(n_1883) );
XNOR2xp5_ASAP7_75t_L g1884 ( .A(n_1885), .B(n_1886), .Y(n_1884) );
AND4x1_ASAP7_75t_L g1886 ( .A(n_1887), .B(n_1889), .C(n_1912), .D(n_1930), .Y(n_1886) );
NOR3xp33_ASAP7_75t_SL g1889 ( .A(n_1890), .B(n_1892), .C(n_1908), .Y(n_1889) );
BUFx2_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
OAI22xp5_ASAP7_75t_L g1892 ( .A1(n_1893), .A2(n_1895), .B1(n_1902), .B2(n_1903), .Y(n_1892) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1894), .Y(n_1893) );
INVx2_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVx2_ASAP7_75t_L g1909 ( .A(n_1910), .Y(n_1909) );
NOR2xp33_ASAP7_75t_L g1930 ( .A(n_1931), .B(n_1932), .Y(n_1930) );
CKINVDCx5p33_ASAP7_75t_R g1936 ( .A(n_1937), .Y(n_1936) );
BUFx2_ASAP7_75t_L g1937 ( .A(n_1938), .Y(n_1937) );
INVx1_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
INVx1_ASAP7_75t_L g1939 ( .A(n_1940), .Y(n_1939) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
CKINVDCx5p33_ASAP7_75t_R g1943 ( .A(n_1944), .Y(n_1943) );
INVxp33_ASAP7_75t_L g1946 ( .A(n_1947), .Y(n_1946) );
HB1xp67_ASAP7_75t_L g1948 ( .A(n_1949), .Y(n_1948) );
NAND3xp33_ASAP7_75t_L g1949 ( .A(n_1950), .B(n_1971), .C(n_1973), .Y(n_1949) );
NOR2xp33_ASAP7_75t_L g1950 ( .A(n_1951), .B(n_1958), .Y(n_1950) );
NAND2xp5_ASAP7_75t_L g1951 ( .A(n_1952), .B(n_1955), .Y(n_1951) );
INVx1_ASAP7_75t_L g1969 ( .A(n_1970), .Y(n_1969) );
INVx2_ASAP7_75t_SL g1977 ( .A(n_1978), .Y(n_1977) );
INVx1_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
HB1xp67_ASAP7_75t_L g1990 ( .A(n_1991), .Y(n_1990) );
endmodule