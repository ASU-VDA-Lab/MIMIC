module real_aes_12158_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_351;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1802;
wire n_727;
wire n_397;
wire n_1083;
wire n_1056;
wire n_1605;
wire n_1855;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_0), .A2(n_425), .B1(n_1031), .B2(n_1371), .C(n_1377), .Y(n_1370) );
AOI21xp33_ASAP7_75t_L g1399 ( .A1(n_0), .A2(n_645), .B(n_1208), .Y(n_1399) );
INVxp67_ASAP7_75t_L g433 ( .A(n_1), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_1), .A2(n_196), .B1(n_495), .B2(n_524), .C(n_529), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g1516 ( .A1(n_2), .A2(n_68), .B1(n_1059), .B2(n_1321), .C(n_1517), .Y(n_1516) );
AOI22xp33_ASAP7_75t_SL g1537 ( .A1(n_2), .A2(n_183), .B1(n_377), .B2(n_610), .Y(n_1537) );
OAI221xp5_ASAP7_75t_L g949 ( .A1(n_3), .A2(n_950), .B1(n_952), .B2(n_958), .C(n_964), .Y(n_949) );
INVx1_ASAP7_75t_L g988 ( .A(n_3), .Y(n_988) );
INVx1_ASAP7_75t_L g1352 ( .A(n_4), .Y(n_1352) );
AOI22xp5_ASAP7_75t_L g1601 ( .A1(n_5), .A2(n_329), .B1(n_1576), .B2(n_1580), .Y(n_1601) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_6), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_7), .A2(n_249), .B1(n_375), .B2(n_386), .C(n_393), .Y(n_374) );
INVx1_ASAP7_75t_L g510 ( .A(n_7), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_8), .A2(n_111), .B1(n_389), .B2(n_941), .C(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g1003 ( .A(n_8), .Y(n_1003) );
OAI221xp5_ASAP7_75t_L g1380 ( .A1(n_9), .A2(n_188), .B1(n_410), .B2(n_419), .C(n_422), .Y(n_1380) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_9), .Y(n_1404) );
AO22x1_ASAP7_75t_L g924 ( .A1(n_10), .A2(n_925), .B1(n_1009), .B2(n_1010), .Y(n_924) );
INVx1_ASAP7_75t_L g1010 ( .A(n_10), .Y(n_1010) );
AOI221xp5_ASAP7_75t_L g1426 ( .A1(n_11), .A2(n_316), .B1(n_939), .B2(n_1427), .C(n_1429), .Y(n_1426) );
INVx1_ASAP7_75t_L g1436 ( .A(n_11), .Y(n_1436) );
INVx1_ASAP7_75t_L g1165 ( .A(n_12), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_13), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_14), .A2(n_307), .B1(n_1100), .B2(n_1102), .Y(n_1099) );
INVx1_ASAP7_75t_L g1131 ( .A(n_14), .Y(n_1131) );
INVx1_ASAP7_75t_L g1412 ( .A(n_15), .Y(n_1412) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_16), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_17), .A2(n_262), .B1(n_665), .B2(n_1512), .Y(n_1511) );
INVxp33_ASAP7_75t_SL g1529 ( .A(n_17), .Y(n_1529) );
AOI22xp33_ASAP7_75t_SL g1804 ( .A1(n_18), .A2(n_154), .B1(n_612), .B2(n_613), .Y(n_1804) );
AOI221xp5_ASAP7_75t_L g1823 ( .A1(n_18), .A2(n_245), .B1(n_1210), .B2(n_1824), .C(n_1826), .Y(n_1823) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_19), .A2(n_158), .B1(n_813), .B2(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g845 ( .A(n_19), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_20), .A2(n_117), .B1(n_408), .B2(n_417), .C(n_422), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_20), .A2(n_117), .B1(n_478), .B2(n_489), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g1060 ( .A1(n_21), .A2(n_83), .B1(n_489), .B2(n_1061), .C(n_1062), .Y(n_1060) );
INVx1_ASAP7_75t_L g1065 ( .A(n_21), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_22), .Y(n_1331) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_23), .A2(n_198), .B1(n_496), .B2(n_1097), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_23), .A2(n_198), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
AOI22xp5_ASAP7_75t_L g1788 ( .A1(n_24), .A2(n_1789), .B1(n_1790), .B2(n_1791), .Y(n_1788) );
CKINVDCx5p33_ASAP7_75t_R g1789 ( .A(n_24), .Y(n_1789) );
INVx1_ASAP7_75t_L g1863 ( .A(n_25), .Y(n_1863) );
OAI22xp5_ASAP7_75t_L g1874 ( .A1(n_25), .A2(n_315), .B1(n_1875), .B2(n_1879), .Y(n_1874) );
AOI22xp5_ASAP7_75t_L g1602 ( .A1(n_26), .A2(n_287), .B1(n_1547), .B2(n_1593), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_27), .A2(n_223), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_27), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1414 ( .A1(n_28), .A2(n_48), .B1(n_1349), .B2(n_1415), .C(n_1416), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_28), .A2(n_290), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
CKINVDCx16_ASAP7_75t_R g1616 ( .A(n_29), .Y(n_1616) );
CKINVDCx5p33_ASAP7_75t_R g1374 ( .A(n_30), .Y(n_1374) );
INVx1_ASAP7_75t_L g1418 ( .A(n_31), .Y(n_1418) );
AOI221xp5_ASAP7_75t_L g1438 ( .A1(n_31), .A2(n_48), .B1(n_1439), .B2(n_1440), .C(n_1441), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_32), .A2(n_324), .B1(n_607), .B2(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g651 ( .A(n_32), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_33), .A2(n_80), .B1(n_918), .B2(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1397 ( .A(n_33), .Y(n_1397) );
INVxp33_ASAP7_75t_L g1263 ( .A(n_34), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_34), .A2(n_101), .B1(n_1291), .B2(n_1292), .C(n_1294), .Y(n_1290) );
INVx1_ASAP7_75t_L g1431 ( .A(n_35), .Y(n_1431) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_36), .A2(n_237), .B1(n_530), .B2(n_662), .C(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g708 ( .A(n_36), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g1272 ( .A1(n_37), .A2(n_171), .B1(n_1273), .B2(n_1275), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_37), .A2(n_171), .B1(n_1305), .B2(n_1307), .Y(n_1304) );
OAI221xp5_ASAP7_75t_L g1466 ( .A1(n_38), .A2(n_103), .B1(n_408), .B2(n_418), .C(n_1467), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1490 ( .A1(n_38), .A2(n_103), .B1(n_671), .B2(n_1173), .Y(n_1490) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_39), .A2(n_131), .B1(n_613), .B2(n_1123), .C(n_1125), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_39), .A2(n_157), .B1(n_1135), .B2(n_1137), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_40), .A2(n_43), .B1(n_761), .B2(n_939), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_40), .A2(n_111), .B1(n_1005), .B2(n_1007), .Y(n_1004) );
INVx1_ASAP7_75t_L g350 ( .A(n_41), .Y(n_350) );
INVx1_ASAP7_75t_L g749 ( .A(n_42), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_42), .A2(n_276), .B1(n_792), .B2(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g1001 ( .A(n_43), .Y(n_1001) );
INVx1_ASAP7_75t_L g736 ( .A(n_44), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_45), .A2(n_115), .B1(n_597), .B2(n_600), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_45), .A2(n_214), .B1(n_643), .B2(n_647), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1597 ( .A1(n_46), .A2(n_165), .B1(n_1576), .B2(n_1580), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g1582 ( .A1(n_47), .A2(n_220), .B1(n_1545), .B2(n_1553), .Y(n_1582) );
AOI22xp33_ASAP7_75t_SL g1277 ( .A1(n_49), .A2(n_302), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_49), .A2(n_302), .B1(n_675), .B2(n_1300), .C(n_1302), .Y(n_1299) );
INVx1_ASAP7_75t_L g616 ( .A(n_50), .Y(n_616) );
INVx1_ASAP7_75t_L g1480 ( .A(n_51), .Y(n_1480) );
INVxp33_ASAP7_75t_L g739 ( .A(n_52), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_52), .A2(n_297), .B1(n_665), .B2(n_780), .C(n_783), .Y(n_779) );
INVx1_ASAP7_75t_L g1095 ( .A(n_53), .Y(n_1095) );
OAI211xp5_ASAP7_75t_SL g1118 ( .A1(n_53), .A2(n_928), .B(n_1119), .C(n_1126), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_54), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g1811 ( .A(n_55), .Y(n_1811) );
INVx1_ASAP7_75t_L g870 ( .A(n_56), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_56), .A2(n_288), .B1(n_897), .B2(n_898), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_57), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_58), .A2(n_108), .B1(n_944), .B2(n_948), .Y(n_943) );
OAI22xp5_ASAP7_75t_SL g973 ( .A1(n_58), .A2(n_108), .B1(n_974), .B2(n_978), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g1591 ( .A1(n_59), .A2(n_136), .B1(n_1576), .B2(n_1580), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_60), .A2(n_340), .B1(n_533), .B2(n_1324), .Y(n_1326) );
OAI22xp33_ASAP7_75t_L g1360 ( .A1(n_60), .A2(n_320), .B1(n_950), .B2(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1189 ( .A(n_61), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_61), .A2(n_284), .B1(n_1195), .B2(n_1196), .C(n_1198), .Y(n_1194) );
AOI22xp33_ASAP7_75t_SL g1280 ( .A1(n_62), .A2(n_134), .B1(n_1275), .B2(n_1278), .Y(n_1280) );
INVxp67_ASAP7_75t_SL g1288 ( .A(n_62), .Y(n_1288) );
AO221x2_ASAP7_75t_L g1603 ( .A1(n_63), .A2(n_247), .B1(n_1547), .B2(n_1593), .C(n_1604), .Y(n_1603) );
CKINVDCx16_ASAP7_75t_R g1617 ( .A(n_64), .Y(n_1617) );
INVx1_ASAP7_75t_L g1498 ( .A(n_65), .Y(n_1498) );
AOI22xp5_ASAP7_75t_SL g1586 ( .A1(n_66), .A2(n_233), .B1(n_1547), .B2(n_1553), .Y(n_1586) );
INVx1_ASAP7_75t_L g768 ( .A(n_67), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g1536 ( .A1(n_68), .A2(n_162), .B1(n_600), .B2(n_604), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g1801 ( .A(n_69), .Y(n_1801) );
INVx1_ASAP7_75t_L g1411 ( .A(n_70), .Y(n_1411) );
INVxp33_ASAP7_75t_SL g1802 ( .A(n_71), .Y(n_1802) );
AOI221xp5_ASAP7_75t_L g1817 ( .A1(n_71), .A2(n_239), .B1(n_628), .B2(n_1818), .C(n_1820), .Y(n_1817) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_72), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_73), .A2(n_179), .B1(n_971), .B2(n_1376), .Y(n_1379) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_73), .A2(n_179), .B1(n_548), .B2(n_807), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_74), .A2(n_318), .B1(n_489), .B2(n_1214), .Y(n_1213) );
OAI221xp5_ASAP7_75t_L g1237 ( .A1(n_74), .A2(n_318), .B1(n_742), .B2(n_743), .C(n_744), .Y(n_1237) );
INVx1_ASAP7_75t_L g766 ( .A(n_75), .Y(n_766) );
CKINVDCx14_ASAP7_75t_R g1563 ( .A(n_76), .Y(n_1563) );
INVx1_ASAP7_75t_L g966 ( .A(n_77), .Y(n_966) );
INVxp67_ASAP7_75t_SL g1513 ( .A(n_78), .Y(n_1513) );
AOI22xp33_ASAP7_75t_SL g1538 ( .A1(n_78), .A2(n_201), .B1(n_377), .B2(n_597), .Y(n_1538) );
AOI22xp33_ASAP7_75t_SL g1805 ( .A1(n_79), .A2(n_245), .B1(n_1278), .B2(n_1806), .Y(n_1805) );
AOI22xp33_ASAP7_75t_L g1828 ( .A1(n_79), .A2(n_154), .B1(n_648), .B2(n_1829), .Y(n_1828) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_80), .A2(n_124), .B1(n_471), .B2(n_1395), .Y(n_1398) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_81), .A2(n_306), .B1(n_560), .B2(n_917), .Y(n_1037) );
INVx1_ASAP7_75t_L g1063 ( .A(n_81), .Y(n_1063) );
INVxp67_ASAP7_75t_SL g1796 ( .A(n_82), .Y(n_1796) );
OAI22xp33_ASAP7_75t_L g1815 ( .A1(n_82), .A2(n_291), .B1(n_621), .B2(n_1816), .Y(n_1815) );
INVx1_ASAP7_75t_L g1066 ( .A(n_83), .Y(n_1066) );
INVx1_ASAP7_75t_L g1226 ( .A(n_84), .Y(n_1226) );
XOR2xp5_ASAP7_75t_L g1315 ( .A(n_85), .B(n_1316), .Y(n_1315) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_86), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g1281 ( .A1(n_87), .A2(n_121), .B1(n_1273), .B2(n_1279), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1298 ( .A(n_87), .Y(n_1298) );
INVx1_ASAP7_75t_L g1350 ( .A(n_88), .Y(n_1350) );
INVx1_ASAP7_75t_L g1799 ( .A(n_89), .Y(n_1799) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_90), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_91), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_92), .A2(n_212), .B1(n_1576), .B2(n_1579), .Y(n_1575) );
CKINVDCx5p33_ASAP7_75t_R g1890 ( .A(n_93), .Y(n_1890) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_94), .A2(n_303), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1339 ( .A(n_94), .Y(n_1339) );
INVx1_ASAP7_75t_L g575 ( .A(n_95), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_95), .A2(n_169), .B1(n_621), .B2(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g1462 ( .A(n_96), .Y(n_1462) );
OAI222xp33_ASAP7_75t_L g1148 ( .A1(n_97), .A2(n_146), .B1(n_300), .B2(n_560), .C1(n_743), .C2(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1175 ( .A(n_97), .Y(n_1175) );
OAI211xp5_ASAP7_75t_SL g880 ( .A1(n_98), .A2(n_881), .B(n_882), .C(n_885), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_98), .A2(n_192), .B1(n_901), .B2(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g771 ( .A(n_99), .Y(n_771) );
AO22x2_ASAP7_75t_L g1011 ( .A1(n_100), .A2(n_1012), .B1(n_1067), .B2(n_1068), .Y(n_1011) );
CKINVDCx14_ASAP7_75t_R g1067 ( .A(n_100), .Y(n_1067) );
INVxp33_ASAP7_75t_SL g1267 ( .A(n_101), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_102), .A2(n_333), .B1(n_671), .B2(n_825), .Y(n_824) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_102), .A2(n_333), .B1(n_408), .B2(n_418), .C(n_696), .Y(n_840) );
INVx1_ASAP7_75t_L g383 ( .A(n_104), .Y(n_383) );
OR2x2_ASAP7_75t_L g415 ( .A(n_104), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g428 ( .A(n_104), .Y(n_428) );
BUFx2_ASAP7_75t_L g563 ( .A(n_104), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_105), .A2(n_142), .B1(n_971), .B2(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1393 ( .A(n_105), .Y(n_1393) );
INVx1_ASAP7_75t_L g772 ( .A(n_106), .Y(n_772) );
INVx1_ASAP7_75t_L g957 ( .A(n_107), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_107), .A2(n_225), .B1(n_629), .B2(n_878), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1212 ( .A(n_109), .Y(n_1212) );
AOI22xp33_ASAP7_75t_SL g1808 ( .A1(n_110), .A2(n_204), .B1(n_1278), .B2(n_1806), .Y(n_1808) );
INVxp33_ASAP7_75t_SL g1832 ( .A(n_110), .Y(n_1832) );
INVx1_ASAP7_75t_L g935 ( .A(n_112), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_112), .A2(n_260), .B1(n_470), .B2(n_629), .Y(n_990) );
INVx1_ASAP7_75t_L g738 ( .A(n_113), .Y(n_738) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_114), .A2(n_325), .B1(n_742), .B2(n_743), .C(n_744), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_114), .A2(n_325), .B1(n_489), .B2(n_778), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_115), .A2(n_272), .B1(n_530), .B2(n_638), .C(n_640), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_116), .A2(n_193), .B1(n_662), .B2(n_782), .C(n_810), .Y(n_809) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_116), .Y(n_849) );
AOI22xp33_ASAP7_75t_SL g1809 ( .A1(n_118), .A2(n_258), .B1(n_612), .B2(n_613), .Y(n_1809) );
INVxp33_ASAP7_75t_L g1831 ( .A(n_118), .Y(n_1831) );
INVx1_ASAP7_75t_L g589 ( .A(n_119), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_119), .A2(n_127), .B1(n_625), .B2(n_628), .C(n_630), .Y(n_624) );
INVxp33_ASAP7_75t_L g1461 ( .A(n_120), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1491 ( .A1(n_120), .A2(n_343), .B1(n_665), .B2(n_1439), .C(n_1492), .Y(n_1491) );
INVxp33_ASAP7_75t_L g1309 ( .A(n_121), .Y(n_1309) );
INVx1_ASAP7_75t_L g1092 ( .A(n_122), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1107 ( .A1(n_122), .A2(n_950), .B1(n_1108), .B2(n_1111), .C(n_1117), .Y(n_1107) );
INVx1_ASAP7_75t_L g1430 ( .A(n_123), .Y(n_1430) );
OAI221xp5_ASAP7_75t_L g1434 ( .A1(n_123), .A2(n_316), .B1(n_823), .B2(n_1178), .C(n_1435), .Y(n_1434) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_124), .A2(n_140), .B1(n_560), .B2(n_917), .Y(n_1384) );
INVx1_ASAP7_75t_L g567 ( .A(n_125), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_126), .A2(n_173), .B1(n_622), .B2(n_778), .Y(n_1514) );
INVxp67_ASAP7_75t_SL g1526 ( .A(n_126), .Y(n_1526) );
INVx1_ASAP7_75t_L g584 ( .A(n_127), .Y(n_584) );
INVx1_ASAP7_75t_L g1266 ( .A(n_128), .Y(n_1266) );
INVx1_ASAP7_75t_L g394 ( .A(n_129), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_130), .A2(n_161), .B1(n_534), .B2(n_662), .C(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g837 ( .A(n_130), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_131), .A2(n_202), .B1(n_1005), .B2(n_1007), .Y(n_1133) );
INVxp67_ASAP7_75t_L g758 ( .A(n_132), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_132), .A2(n_206), .B1(n_530), .B2(n_787), .C(n_789), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_133), .Y(n_683) );
INVxp33_ASAP7_75t_L g1310 ( .A(n_134), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1505 ( .A(n_135), .Y(n_1505) );
AOI22xp5_ASAP7_75t_L g1838 ( .A1(n_136), .A2(n_1839), .B1(n_1844), .B2(n_1926), .Y(n_1838) );
XOR2xp5_ASAP7_75t_L g1847 ( .A(n_136), .B(n_1848), .Y(n_1847) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_137), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_138), .Y(n_884) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_139), .Y(n_1260) );
OAI22xp33_ASAP7_75t_L g1289 ( .A1(n_139), .A2(n_176), .B1(n_478), .B2(n_489), .Y(n_1289) );
INVx1_ASAP7_75t_L g1401 ( .A(n_140), .Y(n_1401) );
INVx1_ASAP7_75t_L g808 ( .A(n_141), .Y(n_808) );
INVx1_ASAP7_75t_L g1390 ( .A(n_142), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_143), .Y(n_1073) );
AOI21xp33_ASAP7_75t_L g877 ( .A1(n_144), .A2(n_530), .B(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_144), .A2(n_175), .B1(n_901), .B2(n_903), .Y(n_900) );
INVxp33_ASAP7_75t_L g1470 ( .A(n_145), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_145), .A2(n_156), .B1(n_1443), .B2(n_1444), .Y(n_1496) );
INVx1_ASAP7_75t_L g1186 ( .A(n_146), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_147), .Y(n_1024) );
INVx1_ASAP7_75t_L g1860 ( .A(n_148), .Y(n_1860) );
OAI22xp5_ASAP7_75t_L g1896 ( .A1(n_148), .A2(n_282), .B1(n_1897), .B2(n_1899), .Y(n_1896) );
AOI22xp5_ASAP7_75t_SL g1585 ( .A1(n_149), .A2(n_172), .B1(n_1576), .B2(n_1580), .Y(n_1585) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_150), .A2(n_192), .B1(n_548), .B2(n_550), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_150), .A2(n_264), .B1(n_898), .B2(n_909), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_151), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_152), .Y(n_883) );
INVx1_ASAP7_75t_L g1551 ( .A(n_153), .Y(n_1551) );
INVx1_ASAP7_75t_L g1020 ( .A(n_155), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g1056 ( .A1(n_155), .A2(n_305), .B1(n_629), .B2(n_1057), .Y(n_1056) );
INVxp67_ASAP7_75t_SL g1477 ( .A(n_156), .Y(n_1477) );
INVx1_ASAP7_75t_L g1120 ( .A(n_157), .Y(n_1120) );
INVx1_ASAP7_75t_L g851 ( .A(n_158), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_159), .A2(n_799), .B1(n_861), .B2(n_862), .Y(n_798) );
INVx1_ASAP7_75t_L g862 ( .A(n_159), .Y(n_862) );
INVx1_ASAP7_75t_L g1483 ( .A(n_160), .Y(n_1483) );
INVx1_ASAP7_75t_L g834 ( .A(n_161), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_162), .A2(n_183), .B1(n_643), .B2(n_1089), .Y(n_1519) );
CKINVDCx16_ASAP7_75t_R g1613 ( .A(n_163), .Y(n_1613) );
INVx1_ASAP7_75t_L g1870 ( .A(n_164), .Y(n_1870) );
OAI22xp33_ASAP7_75t_SL g1921 ( .A1(n_164), .A2(n_181), .B1(n_359), .B2(n_1922), .Y(n_1921) );
INVx1_ASAP7_75t_L g1456 ( .A(n_165), .Y(n_1456) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_166), .A2(n_215), .B1(n_821), .B2(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g832 ( .A(n_166), .Y(n_832) );
INVx1_ASAP7_75t_L g1549 ( .A(n_167), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_167), .B(n_1562), .Y(n_1568) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_168), .A2(n_197), .B1(n_627), .B2(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g688 ( .A(n_168), .Y(n_688) );
INVx1_ASAP7_75t_L g580 ( .A(n_169), .Y(n_580) );
INVx1_ASAP7_75t_L g1157 ( .A(n_170), .Y(n_1157) );
INVx1_ASAP7_75t_L g796 ( .A(n_172), .Y(n_796) );
INVxp67_ASAP7_75t_SL g1527 ( .A(n_173), .Y(n_1527) );
INVx2_ASAP7_75t_L g362 ( .A(n_174), .Y(n_362) );
INVx1_ASAP7_75t_L g872 ( .A(n_175), .Y(n_872) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_176), .Y(n_1261) );
INVxp67_ASAP7_75t_L g1159 ( .A(n_177), .Y(n_1159) );
OAI222xp33_ASAP7_75t_L g1177 ( .A1(n_177), .A2(n_185), .B1(n_271), .B2(n_626), .C1(n_1178), .C2(n_1180), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_178), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_180), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1872 ( .A1(n_181), .A2(n_273), .B1(n_629), .B2(n_782), .Y(n_1872) );
BUFx3_ASAP7_75t_L g473 ( .A(n_182), .Y(n_473) );
INVx1_ASAP7_75t_L g503 ( .A(n_182), .Y(n_503) );
XNOR2x2_ASAP7_75t_L g371 ( .A(n_184), .B(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g1164 ( .A(n_185), .Y(n_1164) );
INVxp67_ASAP7_75t_L g447 ( .A(n_186), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_186), .A2(n_254), .B1(n_533), .B2(n_537), .Y(n_532) );
INVx1_ASAP7_75t_L g1347 ( .A(n_187), .Y(n_1347) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_188), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_189), .A2(n_295), .B1(n_1206), .B2(n_1207), .C(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1233 ( .A(n_189), .Y(n_1233) );
INVx1_ASAP7_75t_L g1015 ( .A(n_190), .Y(n_1015) );
AOI21xp33_ASAP7_75t_L g1058 ( .A1(n_190), .A2(n_470), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1419 ( .A(n_191), .Y(n_1419) );
INVxp67_ASAP7_75t_SL g846 ( .A(n_193), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_194), .A2(n_320), .B1(n_1210), .B2(n_1211), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1335 ( .A1(n_194), .A2(n_340), .B1(n_928), .B2(n_1336), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g1333 ( .A(n_195), .Y(n_1333) );
INVxp67_ASAP7_75t_L g441 ( .A(n_196), .Y(n_441) );
INVx1_ASAP7_75t_L g692 ( .A(n_197), .Y(n_692) );
INVx1_ASAP7_75t_L g476 ( .A(n_199), .Y(n_476) );
INVx1_ASAP7_75t_L g515 ( .A(n_199), .Y(n_515) );
INVx1_ASAP7_75t_L g804 ( .A(n_200), .Y(n_804) );
INVxp33_ASAP7_75t_L g1523 ( .A(n_201), .Y(n_1523) );
INVx1_ASAP7_75t_L g1121 ( .A(n_202), .Y(n_1121) );
INVx1_ASAP7_75t_L g1264 ( .A(n_203), .Y(n_1264) );
INVxp67_ASAP7_75t_SL g1814 ( .A(n_204), .Y(n_1814) );
XNOR2xp5_ASAP7_75t_L g1145 ( .A(n_205), .B(n_1146), .Y(n_1145) );
INVxp67_ASAP7_75t_L g753 ( .A(n_206), .Y(n_753) );
INVxp67_ASAP7_75t_SL g1476 ( .A(n_207), .Y(n_1476) );
AOI221xp5_ASAP7_75t_L g1495 ( .A1(n_207), .A2(n_279), .B1(n_675), .B2(n_1440), .C(n_1441), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_208), .Y(n_681) );
INVxp67_ASAP7_75t_L g1152 ( .A(n_209), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_209), .A2(n_308), .B1(n_782), .B2(n_810), .C(n_1043), .Y(n_1182) );
CKINVDCx20_ASAP7_75t_R g1556 ( .A(n_210), .Y(n_1556) );
OAI21xp33_ASAP7_75t_L g1408 ( .A1(n_211), .A2(n_1409), .B(n_1432), .Y(n_1408) );
INVx1_ASAP7_75t_L g1451 ( .A(n_211), .Y(n_1451) );
INVxp67_ASAP7_75t_SL g1857 ( .A(n_213), .Y(n_1857) );
AOI22xp33_ASAP7_75t_L g1868 ( .A1(n_213), .A2(n_319), .B1(n_629), .B2(n_878), .Y(n_1868) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_214), .A2(n_272), .B1(n_604), .B2(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g838 ( .A(n_215), .Y(n_838) );
INVxp67_ASAP7_75t_SL g1520 ( .A(n_216), .Y(n_1520) );
AOI22xp33_ASAP7_75t_SL g1539 ( .A1(n_216), .A2(n_281), .B1(n_600), .B2(n_612), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_217), .Y(n_1023) );
OA22x2_ASAP7_75t_L g654 ( .A1(n_218), .A2(n_655), .B1(n_721), .B2(n_722), .Y(n_654) );
INVx1_ASAP7_75t_L g722 ( .A(n_218), .Y(n_722) );
XOR2xp5_ASAP7_75t_L g1367 ( .A(n_219), .B(n_1368), .Y(n_1367) );
CKINVDCx14_ASAP7_75t_R g1605 ( .A(n_221), .Y(n_1605) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_222), .A2(n_268), .B1(n_470), .B2(n_629), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_222), .A2(n_336), .B1(n_917), .B2(n_918), .Y(n_916) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_223), .Y(n_1116) );
INVx1_ASAP7_75t_L g1425 ( .A(n_224), .Y(n_1425) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_224), .A2(n_293), .B1(n_790), .B2(n_793), .C(n_1208), .Y(n_1446) );
INVx1_ASAP7_75t_L g955 ( .A(n_225), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g1353 ( .A(n_226), .Y(n_1353) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_227), .A2(n_267), .B1(n_810), .B2(n_1217), .C(n_1219), .Y(n_1216) );
INVx1_ASAP7_75t_L g1244 ( .A(n_227), .Y(n_1244) );
INVx1_ASAP7_75t_L g1853 ( .A(n_228), .Y(n_1853) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_229), .A2(n_234), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1047 ( .A(n_229), .Y(n_1047) );
OA332x1_ASAP7_75t_L g1013 ( .A1(n_230), .A2(n_425), .A3(n_1014), .B1(n_1019), .B2(n_1022), .B3(n_1025), .C1(n_1030), .C2(n_1031), .Y(n_1013) );
AOI21xp5_ASAP7_75t_L g1052 ( .A1(n_230), .A2(n_819), .B(n_1053), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1508 ( .A1(n_231), .A2(n_243), .B1(n_1207), .B2(n_1324), .C(n_1509), .Y(n_1508) );
INVxp33_ASAP7_75t_SL g1531 ( .A(n_231), .Y(n_1531) );
INVx1_ASAP7_75t_L g828 ( .A(n_232), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_234), .A2(n_306), .B1(n_470), .B2(n_629), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_235), .A2(n_242), .B1(n_533), .B2(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1345 ( .A(n_235), .Y(n_1345) );
CKINVDCx20_ASAP7_75t_R g1502 ( .A(n_236), .Y(n_1502) );
INVx1_ASAP7_75t_L g703 ( .A(n_237), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_238), .A2(n_241), .B1(n_669), .B2(n_671), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_238), .A2(n_241), .B1(n_418), .B2(n_695), .C(n_696), .Y(n_694) );
INVxp33_ASAP7_75t_SL g1798 ( .A(n_239), .Y(n_1798) );
INVx1_ASAP7_75t_L g1174 ( .A(n_240), .Y(n_1174) );
INVx1_ASAP7_75t_L g1343 ( .A(n_242), .Y(n_1343) );
INVxp33_ASAP7_75t_L g1533 ( .A(n_243), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_244), .Y(n_962) );
INVx1_ASAP7_75t_L g1254 ( .A(n_246), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_248), .A2(n_263), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g689 ( .A(n_248), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_249), .A2(n_338), .B1(n_495), .B2(n_498), .C(n_504), .Y(n_494) );
INVx1_ASAP7_75t_L g1086 ( .A(n_250), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g1311 ( .A(n_251), .Y(n_1311) );
INVx1_ASAP7_75t_L g472 ( .A(n_252), .Y(n_472) );
BUFx3_ASAP7_75t_L g488 ( .A(n_252), .Y(n_488) );
AO221x2_ASAP7_75t_L g1544 ( .A1(n_253), .A2(n_317), .B1(n_1545), .B2(n_1552), .C(n_1555), .Y(n_1544) );
INVxp67_ASAP7_75t_L g430 ( .A(n_254), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g889 ( .A1(n_255), .A2(n_534), .B(n_819), .Y(n_889) );
INVx1_ASAP7_75t_L g914 ( .A(n_255), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_256), .A2(n_257), .B1(n_1547), .B2(n_1593), .Y(n_1592) );
INVxp67_ASAP7_75t_SL g1822 ( .A(n_258), .Y(n_1822) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_259), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_259), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_259), .B(n_322), .Y(n_416) );
INVx1_ASAP7_75t_L g464 ( .A(n_259), .Y(n_464) );
INVx1_ASAP7_75t_L g933 ( .A(n_260), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g1892 ( .A(n_261), .Y(n_1892) );
INVxp33_ASAP7_75t_SL g1534 ( .A(n_262), .Y(n_1534) );
INVx1_ASAP7_75t_L g691 ( .A(n_263), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_264), .A2(n_807), .B1(n_868), .B2(n_873), .C(n_879), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_265), .Y(n_959) );
OR2x2_ASAP7_75t_L g475 ( .A(n_266), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g483 ( .A(n_266), .Y(n_483) );
INVx1_ASAP7_75t_L g1242 ( .A(n_267), .Y(n_1242) );
INVx1_ASAP7_75t_L g915 ( .A(n_268), .Y(n_915) );
INVx1_ASAP7_75t_L g1154 ( .A(n_269), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_270), .A2(n_289), .B1(n_378), .B2(n_856), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1386 ( .A1(n_270), .A2(n_289), .B1(n_550), .B2(n_881), .Y(n_1386) );
INVxp67_ASAP7_75t_L g1162 ( .A(n_271), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g1905 ( .A1(n_273), .A2(n_315), .B1(n_1906), .B2(n_1908), .Y(n_1905) );
INVx1_ASAP7_75t_L g1372 ( .A(n_274), .Y(n_1372) );
AOI21xp33_ASAP7_75t_L g1391 ( .A1(n_274), .A2(n_530), .B(n_782), .Y(n_1391) );
INVx1_ASAP7_75t_L g1485 ( .A(n_275), .Y(n_1485) );
INVxp67_ASAP7_75t_L g763 ( .A(n_276), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_277), .A2(n_314), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
INVx1_ASAP7_75t_L g1231 ( .A(n_277), .Y(n_1231) );
AOI22xp5_ASAP7_75t_SL g1598 ( .A1(n_278), .A2(n_283), .B1(n_1547), .B2(n_1553), .Y(n_1598) );
INVxp33_ASAP7_75t_SL g1472 ( .A(n_279), .Y(n_1472) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_280), .A2(n_286), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g636 ( .A(n_280), .Y(n_636) );
INVxp33_ASAP7_75t_SL g1522 ( .A(n_281), .Y(n_1522) );
INVx1_ASAP7_75t_L g1859 ( .A(n_282), .Y(n_1859) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_284), .A2(n_304), .B1(n_661), .B2(n_663), .C(n_1191), .Y(n_1190) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_285), .Y(n_1222) );
INVx1_ASAP7_75t_L g650 ( .A(n_286), .Y(n_650) );
INVx1_ASAP7_75t_L g874 ( .A(n_288), .Y(n_874) );
INVxp67_ASAP7_75t_SL g1417 ( .A(n_290), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g1795 ( .A(n_291), .Y(n_1795) );
INVx1_ASAP7_75t_L g1871 ( .A(n_292), .Y(n_1871) );
OAI211xp5_ASAP7_75t_SL g1912 ( .A1(n_292), .A2(n_1473), .B(n_1913), .C(n_1917), .Y(n_1912) );
INVx1_ASAP7_75t_L g1424 ( .A(n_293), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_294), .A2(n_864), .B1(n_919), .B2(n_920), .Y(n_863) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_294), .Y(n_919) );
INVx1_ASAP7_75t_L g1235 ( .A(n_295), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_296), .Y(n_555) );
INVxp33_ASAP7_75t_L g734 ( .A(n_297), .Y(n_734) );
OAI221xp5_ASAP7_75t_SL g1422 ( .A1(n_298), .A2(n_332), .B1(n_757), .B2(n_850), .C(n_1423), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_298), .A2(n_332), .B1(n_648), .B2(n_878), .Y(n_1447) );
INVx1_ASAP7_75t_L g1486 ( .A(n_299), .Y(n_1486) );
INVx1_ASAP7_75t_L g1171 ( .A(n_300), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_301), .Y(n_1028) );
INVx1_ASAP7_75t_L g1340 ( .A(n_303), .Y(n_1340) );
OAI332xp33_ASAP7_75t_L g1150 ( .A1(n_304), .A2(n_425), .A3(n_860), .B1(n_1036), .B2(n_1151), .B3(n_1155), .C1(n_1158), .C2(n_1163), .Y(n_1150) );
INVx1_ASAP7_75t_L g1016 ( .A(n_305), .Y(n_1016) );
INVx1_ASAP7_75t_L g1129 ( .A(n_307), .Y(n_1129) );
INVx1_ASAP7_75t_L g1156 ( .A(n_308), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
AND3x2_ASAP7_75t_L g1550 ( .A(n_309), .B(n_350), .C(n_1551), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_309), .B(n_350), .Y(n_1560) );
INVx2_ASAP7_75t_L g363 ( .A(n_310), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_311), .A2(n_334), .B1(n_498), .B2(n_661), .Y(n_676) );
INVx1_ASAP7_75t_L g702 ( .A(n_311), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g927 ( .A1(n_312), .A2(n_928), .B(n_932), .C(n_937), .Y(n_927) );
INVx1_ASAP7_75t_L g989 ( .A(n_312), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_313), .A2(n_328), .B1(n_792), .B2(n_1041), .Y(n_1221) );
INVx1_ASAP7_75t_L g1240 ( .A(n_313), .Y(n_1240) );
INVx1_ASAP7_75t_L g1236 ( .A(n_314), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1855 ( .A(n_319), .Y(n_1855) );
INVx1_ASAP7_75t_L g1852 ( .A(n_321), .Y(n_1852) );
INVx1_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
INVx2_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
OR2x2_ASAP7_75t_L g865 ( .A(n_323), .B(n_559), .Y(n_865) );
INVx1_ASAP7_75t_L g619 ( .A(n_324), .Y(n_619) );
INVx1_ASAP7_75t_L g1464 ( .A(n_326), .Y(n_1464) );
INVx1_ASAP7_75t_L g1357 ( .A(n_327), .Y(n_1357) );
INVx1_ASAP7_75t_L g1245 ( .A(n_328), .Y(n_1245) );
INVx1_ASAP7_75t_L g817 ( .A(n_330), .Y(n_817) );
INVx1_ASAP7_75t_L g1070 ( .A(n_331), .Y(n_1070) );
INVx1_ASAP7_75t_L g711 ( .A(n_334), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_335), .Y(n_1225) );
INVx1_ASAP7_75t_L g886 ( .A(n_336), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_337), .Y(n_1021) );
INVxp33_ASAP7_75t_SL g400 ( .A(n_338), .Y(n_400) );
INVx1_ASAP7_75t_L g1082 ( .A(n_339), .Y(n_1082) );
INVx1_ASAP7_75t_L g803 ( .A(n_341), .Y(n_803) );
INVx1_ASAP7_75t_L g1864 ( .A(n_342), .Y(n_1864) );
INVxp33_ASAP7_75t_L g1465 ( .A(n_343), .Y(n_1465) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_366), .B(n_1541), .Y(n_344) );
INVx3_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
AND2x4_ASAP7_75t_L g1843 ( .A(n_348), .B(n_354), .Y(n_1843) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_SL g1837 ( .A(n_349), .Y(n_1837) );
NAND2xp5_ASAP7_75t_L g1929 ( .A(n_349), .B(n_351), .Y(n_1929) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_351), .B(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x6_ASAP7_75t_L g1925 ( .A(n_356), .B(n_563), .Y(n_1925) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g595 ( .A(n_357), .B(n_365), .Y(n_595) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g426 ( .A(n_358), .B(n_427), .Y(n_426) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g432 ( .A(n_360), .Y(n_432) );
OR2x2_ASAP7_75t_L g560 ( .A(n_360), .B(n_415), .Y(n_560) );
BUFx2_ASAP7_75t_L g701 ( .A(n_360), .Y(n_701) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_360), .Y(n_748) );
INVx2_ASAP7_75t_SL g844 ( .A(n_360), .Y(n_844) );
INVx2_ASAP7_75t_SL g961 ( .A(n_360), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g1416 ( .A1(n_360), .A2(n_436), .B1(n_1417), .B2(n_1418), .Y(n_1416) );
OAI22xp33_ASAP7_75t_L g1429 ( .A1(n_360), .A2(n_436), .B1(n_1430), .B2(n_1431), .Y(n_1429) );
HB1xp67_ASAP7_75t_L g1862 ( .A(n_360), .Y(n_1862) );
OR2x6_ASAP7_75t_L g1906 ( .A(n_360), .B(n_1907), .Y(n_1906) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
AND2x2_ASAP7_75t_L g399 ( .A(n_362), .B(n_363), .Y(n_399) );
AND2x4_ASAP7_75t_L g406 ( .A(n_362), .B(n_392), .Y(n_406) );
INVx1_ASAP7_75t_L g439 ( .A(n_362), .Y(n_439) );
INVx1_ASAP7_75t_L g381 ( .A(n_363), .Y(n_381) );
INVx2_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
INVx1_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
INVx1_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_363), .B(n_379), .Y(n_446) );
AND2x4_ASAP7_75t_L g1918 ( .A(n_364), .B(n_413), .Y(n_1918) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_1140), .B2(n_1540), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
XNOR2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_725), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
XNOR2x1_ASAP7_75t_L g370 ( .A(n_371), .B(n_565), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_465), .Y(n_372) );
NOR3xp33_ASAP7_75t_SL g373 ( .A(n_374), .B(n_407), .C(n_423), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_376), .A2(n_396), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_376), .A2(n_387), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_376), .A2(n_396), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_376), .A2(n_396), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g590 ( .A(n_377), .B(n_382), .Y(n_590) );
INVx2_ASAP7_75t_SL g608 ( .A(n_377), .Y(n_608) );
AND2x2_ASAP7_75t_L g693 ( .A(n_377), .B(n_382), .Y(n_693) );
AND2x2_ASAP7_75t_L g740 ( .A(n_377), .B(n_382), .Y(n_740) );
AND2x2_ASAP7_75t_L g839 ( .A(n_377), .B(n_382), .Y(n_839) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g902 ( .A(n_378), .Y(n_902) );
AND2x2_ASAP7_75t_L g934 ( .A(n_378), .B(n_384), .Y(n_934) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_378), .Y(n_939) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_378), .Y(n_1415) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x6_ASAP7_75t_L g388 ( .A(n_382), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g396 ( .A(n_382), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g403 ( .A(n_382), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g833 ( .A(n_382), .B(n_710), .Y(n_833) );
AND2x2_ASAP7_75t_L g835 ( .A(n_382), .B(n_602), .Y(n_835) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_382), .B(n_971), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_382), .A2(n_910), .B1(n_1422), .B2(n_1426), .Y(n_1421) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g461 ( .A(n_383), .Y(n_461) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_383), .B(n_475), .Y(n_1000) );
INVx2_ASAP7_75t_L g931 ( .A(n_384), .Y(n_931) );
AND2x4_ASAP7_75t_L g951 ( .A(n_384), .B(n_606), .Y(n_951) );
INVx1_ASAP7_75t_L g427 ( .A(n_385), .Y(n_427) );
INVx1_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_388), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_388), .A2(n_403), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_388), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_388), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_388), .A2(n_1268), .B1(n_1461), .B2(n_1462), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_388), .A2(n_1529), .B1(n_1530), .B2(n_1531), .Y(n_1528) );
AOI22xp33_ASAP7_75t_L g1797 ( .A1(n_388), .A2(n_585), .B1(n_1798), .B2(n_1799), .Y(n_1797) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_389), .B(n_414), .Y(n_422) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g582 ( .A(n_390), .Y(n_582) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_390), .Y(n_602) );
BUFx3_ASAP7_75t_L g899 ( .A(n_390), .Y(n_899) );
BUFx6f_ASAP7_75t_L g1376 ( .A(n_390), .Y(n_1376) );
AND2x4_ASAP7_75t_L g1914 ( .A(n_390), .B(n_1915), .Y(n_1914) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_400), .B2(n_401), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_394), .A2(n_505), .B1(n_510), .B2(n_511), .C(n_514), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_395), .A2(n_1266), .B1(n_1267), .B2(n_1268), .Y(n_1265) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_396), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_396), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_396), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_396), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_396), .A2(n_740), .B1(n_914), .B2(n_915), .C(n_916), .Y(n_913) );
INVx1_ASAP7_75t_L g1195 ( .A(n_396), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1800 ( .A1(n_396), .A2(n_693), .B1(n_1801), .B2(n_1802), .Y(n_1800) );
BUFx3_ASAP7_75t_L g612 ( .A(n_397), .Y(n_612) );
BUFx2_ASAP7_75t_L g897 ( .A(n_397), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_397), .A2(n_582), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g971 ( .A(n_398), .Y(n_971) );
INVx2_ASAP7_75t_L g1274 ( .A(n_398), .Y(n_1274) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_399), .Y(n_606) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g585 ( .A(n_403), .Y(n_585) );
BUFx2_ASAP7_75t_L g735 ( .A(n_403), .Y(n_735) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_403), .Y(n_1197) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_403), .Y(n_1232) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_403), .Y(n_1268) );
BUFx2_ASAP7_75t_L g1530 ( .A(n_403), .Y(n_1530) );
BUFx3_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
INVx2_ASAP7_75t_L g850 ( .A(n_404), .Y(n_850) );
INVx1_ASAP7_75t_L g956 ( .A(n_404), .Y(n_956) );
INVx1_ASAP7_75t_SL g1373 ( .A(n_404), .Y(n_1373) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g710 ( .A(n_405), .Y(n_710) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_405), .Y(n_762) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_406), .Y(n_599) );
INVx1_ASAP7_75t_L g857 ( .A(n_406), .Y(n_857) );
INVx1_ASAP7_75t_L g1911 ( .A(n_406), .Y(n_1911) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g742 ( .A(n_409), .Y(n_742) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_410), .Y(n_695) );
NAND2x1_ASAP7_75t_SL g410 ( .A(n_411), .B(n_414), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g944 ( .A(n_411), .B(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_411), .A2(n_420), .B1(n_1331), .B2(n_1333), .Y(n_1359) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_413), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_414), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g572 ( .A(n_414), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g578 ( .A(n_414), .B(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g581 ( .A(n_414), .B(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g947 ( .A(n_416), .Y(n_947) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx4f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx4f_ASAP7_75t_L g743 ( .A(n_419), .Y(n_743) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g948 ( .A(n_421), .B(n_946), .Y(n_948) );
BUFx3_ASAP7_75t_L g696 ( .A(n_422), .Y(n_696) );
BUFx2_ASAP7_75t_L g744 ( .A(n_422), .Y(n_744) );
BUFx2_ASAP7_75t_L g1467 ( .A(n_422), .Y(n_1467) );
OAI33xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_429), .A3(n_440), .B1(n_450), .B2(n_453), .B3(n_458), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g697 ( .A1(n_425), .A2(n_458), .A3(n_698), .B1(n_704), .B2(n_712), .B3(n_716), .Y(n_697) );
OAI33xp33_ASAP7_75t_L g745 ( .A1(n_425), .A2(n_458), .A3(n_746), .B1(n_754), .B2(n_764), .B3(n_769), .Y(n_745) );
OAI33xp33_ASAP7_75t_L g841 ( .A1(n_425), .A2(n_842), .A3(n_847), .B1(n_852), .B2(n_858), .B3(n_860), .Y(n_841) );
OAI33xp33_ASAP7_75t_L g1238 ( .A1(n_425), .A2(n_860), .A3(n_1239), .B1(n_1243), .B2(n_1247), .B3(n_1253), .Y(n_1238) );
OAI33xp33_ASAP7_75t_L g1468 ( .A1(n_425), .A2(n_458), .A3(n_1469), .B1(n_1475), .B2(n_1478), .B3(n_1484), .Y(n_1468) );
OAI33xp33_ASAP7_75t_L g1850 ( .A1(n_425), .A2(n_1851), .A3(n_1854), .B1(n_1858), .B2(n_1861), .B3(n_1865), .Y(n_1850) );
OR2x6_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g1907 ( .A(n_427), .Y(n_1907) );
BUFx2_ASAP7_75t_L g554 ( .A(n_428), .Y(n_554) );
INVx2_ASAP7_75t_L g594 ( .A(n_428), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_431), .A2(n_442), .B1(n_451), .B2(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g770 ( .A(n_432), .Y(n_770) );
INVx1_ASAP7_75t_L g1241 ( .A(n_432), .Y(n_1241) );
OAI22xp5_ASAP7_75t_SL g1163 ( .A1(n_434), .A2(n_770), .B1(n_1164), .B2(n_1165), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_434), .A2(n_1471), .B1(n_1485), .B2(n_1486), .Y(n_1484) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g456 ( .A(n_436), .Y(n_456) );
BUFx3_ASAP7_75t_L g859 ( .A(n_436), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_436), .A2(n_748), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_436), .A2(n_770), .B1(n_1352), .B2(n_1353), .C(n_1354), .Y(n_1351) );
OAI22xp33_ASAP7_75t_L g1851 ( .A1(n_436), .A2(n_748), .B1(n_1852), .B2(n_1853), .Y(n_1851) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_L g720 ( .A(n_438), .B(n_439), .Y(n_720) );
INVx1_ASAP7_75t_L g574 ( .A(n_439), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_447), .B2(n_448), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_442), .A2(n_1112), .B1(n_1113), .B2(n_1116), .Y(n_1111) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_443), .A2(n_1347), .B1(n_1348), .B2(n_1350), .Y(n_1346) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g848 ( .A(n_444), .Y(n_848) );
INVx2_ASAP7_75t_L g1153 ( .A(n_444), .Y(n_1153) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g757 ( .A(n_445), .Y(n_757) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g707 ( .A(n_446), .Y(n_707) );
BUFx2_ASAP7_75t_L g954 ( .A(n_446), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_448), .A2(n_454), .B1(n_455), .B2(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_449), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_451), .A2(n_454), .B1(n_547), .B2(n_549), .Y(n_546) );
AOI211xp5_ASAP7_75t_L g467 ( .A1(n_452), .A2(n_468), .B(n_477), .C(n_494), .Y(n_467) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_456), .A2(n_699), .B1(n_702), .B2(n_703), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_456), .A2(n_960), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_457), .A2(n_517), .B1(n_523), .B2(n_532), .C(n_540), .Y(n_516) );
INVx1_ASAP7_75t_L g1282 ( .A(n_458), .Y(n_1282) );
CKINVDCx8_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_L g614 ( .A(n_460), .Y(n_614) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g977 ( .A(n_461), .B(n_480), .Y(n_977) );
INVx2_ASAP7_75t_L g911 ( .A(n_462), .Y(n_911) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g1916 ( .A(n_463), .Y(n_1916) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_551), .B1(n_555), .B2(n_556), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_516), .C(n_546), .Y(n_466) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI211xp5_ASAP7_75t_SL g618 ( .A1(n_469), .A2(n_619), .B(n_620), .C(n_624), .Y(n_618) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_469), .A2(n_766), .B(n_777), .C(n_779), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g1204 ( .A1(n_469), .A2(n_1205), .B1(n_1209), .B2(n_1212), .C(n_1213), .Y(n_1204) );
AOI211xp5_ASAP7_75t_L g1287 ( .A1(n_469), .A2(n_1288), .B(n_1289), .C(n_1290), .Y(n_1287) );
AOI211xp5_ASAP7_75t_SL g1489 ( .A1(n_469), .A2(n_1480), .B(n_1490), .C(n_1491), .Y(n_1489) );
AOI221xp5_ASAP7_75t_L g1507 ( .A1(n_469), .A2(n_1508), .B1(n_1511), .B2(n_1513), .C(n_1514), .Y(n_1507) );
AOI211xp5_ASAP7_75t_L g1813 ( .A1(n_469), .A2(n_1814), .B(n_1815), .C(n_1817), .Y(n_1813) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
INVx2_ASAP7_75t_SL g788 ( .A(n_470), .Y(n_788) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g497 ( .A(n_471), .Y(n_497) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_471), .Y(n_627) );
BUFx2_ASAP7_75t_L g675 ( .A(n_471), .Y(n_675) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_471), .Y(n_782) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_471), .Y(n_821) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_471), .Y(n_878) );
INVx2_ASAP7_75t_SL g998 ( .A(n_471), .Y(n_998) );
AND2x6_ASAP7_75t_L g1898 ( .A(n_471), .B(n_1877), .Y(n_1898) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g509 ( .A(n_472), .Y(n_509) );
INVx2_ASAP7_75t_L g493 ( .A(n_473), .Y(n_493) );
AND2x2_ASAP7_75t_L g522 ( .A(n_473), .B(n_488), .Y(n_522) );
AND2x4_ASAP7_75t_L g520 ( .A(n_474), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g666 ( .A(n_474), .B(n_627), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_474), .A2(n_520), .B1(n_678), .B2(n_1165), .C(n_1177), .Y(n_1176) );
AOI222xp33_ASAP7_75t_L g1433 ( .A1(n_474), .A2(n_670), .B1(n_672), .B2(n_1411), .C1(n_1412), .C2(n_1434), .Y(n_1433) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g548 ( .A(n_475), .B(n_513), .Y(n_548) );
OR2x2_ASAP7_75t_L g550 ( .A(n_475), .B(n_501), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g1039 ( .A1(n_475), .A2(n_1040), .B(n_1042), .C(n_1044), .Y(n_1039) );
INVx1_ASAP7_75t_L g481 ( .A(n_476), .Y(n_481) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g621 ( .A(n_479), .Y(n_621) );
INVx1_ASAP7_75t_L g778 ( .A(n_479), .Y(n_778) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_479), .Y(n_1061) );
INVx1_ASAP7_75t_L g1214 ( .A(n_479), .Y(n_1214) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_484), .Y(n_479) );
AND2x2_ASAP7_75t_L g490 ( .A(n_480), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g544 ( .A(n_480), .Y(n_544) );
AND2x2_ASAP7_75t_L g564 ( .A(n_480), .B(n_536), .Y(n_564) );
AND2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_491), .Y(n_623) );
AND2x4_ASAP7_75t_L g670 ( .A(n_480), .B(n_484), .Y(n_670) );
AND2x4_ASAP7_75t_L g672 ( .A(n_480), .B(n_491), .Y(n_672) );
BUFx2_ASAP7_75t_L g679 ( .A(n_480), .Y(n_679) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_L g514 ( .A(n_482), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g531 ( .A(n_483), .B(n_515), .Y(n_531) );
INVx1_ASAP7_75t_L g1878 ( .A(n_483), .Y(n_1878) );
HB1xp67_ASAP7_75t_L g1882 ( .A(n_483), .Y(n_1882) );
INVx1_ASAP7_75t_L g1887 ( .A(n_483), .Y(n_1887) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_484), .A2(n_491), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g975 ( .A(n_485), .Y(n_975) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1889 ( .A(n_486), .Y(n_1889) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g536 ( .A(n_487), .B(n_493), .Y(n_536) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g502 ( .A(n_488), .B(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g979 ( .A(n_491), .Y(n_979) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x6_ASAP7_75t_L g1891 ( .A(n_492), .B(n_1878), .Y(n_1891) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g1188 ( .A(n_499), .Y(n_1188) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g794 ( .A(n_500), .Y(n_794) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g1395 ( .A(n_501), .Y(n_1395) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_502), .Y(n_629) );
INVx1_ASAP7_75t_L g1006 ( .A(n_502), .Y(n_1006) );
INVx1_ASAP7_75t_L g1293 ( .A(n_502), .Y(n_1293) );
INVx1_ASAP7_75t_L g508 ( .A(n_503), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g1869 ( .A1(n_505), .A2(n_869), .B1(n_1870), .B2(n_1871), .C(n_1872), .Y(n_1869) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g631 ( .A(n_507), .Y(n_631) );
BUFx4f_ASAP7_75t_L g876 ( .A(n_507), .Y(n_876) );
INVx2_ASAP7_75t_L g1008 ( .A(n_507), .Y(n_1008) );
INVx1_ASAP7_75t_L g1050 ( .A(n_507), .Y(n_1050) );
INVx1_ASAP7_75t_L g1085 ( .A(n_507), .Y(n_1085) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
OR2x2_ASAP7_75t_L g513 ( .A(n_508), .B(n_509), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_511), .A2(n_1092), .B1(n_1093), .B2(n_1095), .C(n_1096), .Y(n_1091) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g784 ( .A(n_512), .Y(n_784) );
INVx2_ASAP7_75t_L g869 ( .A(n_512), .Y(n_869) );
INVx1_ASAP7_75t_L g1136 ( .A(n_512), .Y(n_1136) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g633 ( .A(n_513), .Y(n_633) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_513), .Y(n_1081) );
INVx1_ASAP7_75t_L g1179 ( .A(n_513), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1875 ( .A(n_513), .B(n_1876), .Y(n_1875) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_514), .Y(n_634) );
INVx1_ASAP7_75t_L g663 ( .A(n_514), .Y(n_663) );
INVx2_ASAP7_75t_SL g819 ( .A(n_514), .Y(n_819) );
AND2x4_ASAP7_75t_L g986 ( .A(n_514), .B(n_563), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_514), .Y(n_1208) );
OAI221xp5_ASAP7_75t_L g1492 ( .A1(n_514), .A2(n_1050), .B1(n_1136), .B2(n_1462), .C(n_1464), .Y(n_1492) );
INVx2_ASAP7_75t_L g1510 ( .A(n_514), .Y(n_1510) );
INVx1_ASAP7_75t_L g1903 ( .A(n_515), .Y(n_1903) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_519), .A2(n_542), .B1(n_636), .B2(n_637), .C(n_642), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_519), .A2(n_542), .B1(n_768), .B2(n_786), .C(n_791), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_519), .A2(n_678), .B1(n_1216), .B2(n_1221), .C(n_1222), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g1515 ( .A1(n_519), .A2(n_542), .B1(n_1516), .B2(n_1519), .C(n_1520), .Y(n_1515) );
AOI221xp5_ASAP7_75t_L g1821 ( .A1(n_519), .A2(n_542), .B1(n_1822), .B2(n_1823), .C(n_1828), .Y(n_1821) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_520), .A2(n_674), .B1(n_676), .B2(n_677), .C(n_678), .Y(n_673) );
INVx2_ASAP7_75t_SL g807 ( .A(n_520), .Y(n_807) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_520), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1494 ( .A(n_520), .Y(n_1494) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_521), .Y(n_641) );
AND2x4_ASAP7_75t_L g678 ( .A(n_521), .B(n_679), .Y(n_678) );
BUFx4f_ASAP7_75t_L g1043 ( .A(n_521), .Y(n_1043) );
INVx1_ASAP7_75t_L g1192 ( .A(n_521), .Y(n_1192) );
BUFx3_ASAP7_75t_L g1206 ( .A(n_521), .Y(n_1206) );
INVx2_ASAP7_75t_SL g1220 ( .A(n_521), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_521), .A2(n_627), .B1(n_1431), .B2(n_1436), .Y(n_1435) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_522), .Y(n_528) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g662 ( .A(n_527), .Y(n_662) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_528), .Y(n_545) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_528), .Y(n_790) );
INVx1_ASAP7_75t_L g993 ( .A(n_528), .Y(n_993) );
AND2x4_ASAP7_75t_L g1894 ( .A(n_528), .B(n_1895), .Y(n_1894) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g1827 ( .A(n_530), .Y(n_1827) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g811 ( .A(n_531), .Y(n_811) );
INVx1_ASAP7_75t_L g982 ( .A(n_531), .Y(n_982) );
INVx1_ASAP7_75t_L g1059 ( .A(n_531), .Y(n_1059) );
INVx2_ASAP7_75t_L g1079 ( .A(n_531), .Y(n_1079) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_534), .B(n_999), .Y(n_1002) );
A2O1A1Ixp33_ASAP7_75t_L g1400 ( .A1(n_534), .A2(n_1401), .B(n_1402), .C(n_1406), .Y(n_1400) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g1053 ( .A(n_535), .Y(n_1053) );
INVx1_ASAP7_75t_L g1829 ( .A(n_535), .Y(n_1829) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx6_ASAP7_75t_L g646 ( .A(n_536), .Y(n_646) );
BUFx2_ASAP7_75t_L g1306 ( .A(n_536), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1880 ( .A(n_536), .B(n_1881), .Y(n_1880) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI221xp5_ASAP7_75t_SL g1181 ( .A1(n_538), .A2(n_1154), .B1(n_1157), .B2(n_1178), .C(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_539), .Y(n_648) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_539), .Y(n_815) );
INVx1_ASAP7_75t_L g823 ( .A(n_539), .Y(n_823) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_539), .Y(n_1041) );
INVx2_ASAP7_75t_L g1180 ( .A(n_539), .Y(n_1180) );
AND2x6_ASAP7_75t_L g1900 ( .A(n_539), .B(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g1296 ( .A1(n_542), .A2(n_1297), .B1(n_1298), .B2(n_1299), .C(n_1304), .Y(n_1296) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g1816 ( .A(n_544), .B(n_979), .Y(n_1816) );
INVx1_ASAP7_75t_L g1325 ( .A(n_545), .Y(n_1325) );
INVx1_ASAP7_75t_L g1518 ( .A(n_545), .Y(n_1518) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_547), .A2(n_549), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_547), .A2(n_549), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_547), .A2(n_549), .B1(n_771), .B2(n_772), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_547), .A2(n_549), .B1(n_803), .B2(n_804), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_547), .A2(n_549), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_547), .A2(n_549), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_547), .A2(n_549), .B1(n_1483), .B2(n_1485), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_547), .A2(n_549), .B1(n_1522), .B2(n_1523), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g1830 ( .A1(n_547), .A2(n_549), .B1(n_1831), .B2(n_1832), .Y(n_1830) );
INVx6_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx5_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_552), .A2(n_927), .B(n_949), .Y(n_926) );
BUFx8_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g1202 ( .A(n_553), .Y(n_1202) );
AOI31xp33_ASAP7_75t_L g1286 ( .A1(n_553), .A2(n_1287), .A3(n_1296), .B(n_1308), .Y(n_1286) );
OAI31xp33_ASAP7_75t_L g1334 ( .A1(n_553), .A2(n_1335), .A3(n_1337), .B(n_1360), .Y(n_1334) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g653 ( .A(n_554), .Y(n_653) );
AND2x4_ASAP7_75t_L g1902 ( .A(n_554), .B(n_1903), .Y(n_1902) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_558), .A2(n_616), .B(n_617), .Y(n_615) );
AOI21xp33_ASAP7_75t_SL g773 ( .A1(n_558), .A2(n_774), .B(n_775), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g1504 ( .A1(n_558), .A2(n_1505), .B(n_1506), .Y(n_1504) );
AOI21xp5_ASAP7_75t_L g1810 ( .A1(n_558), .A2(n_1811), .B(n_1812), .Y(n_1810) );
INVx5_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g684 ( .A(n_559), .Y(n_684) );
INVx1_ASAP7_75t_L g1227 ( .A(n_559), .Y(n_1227) );
INVx2_ASAP7_75t_L g1284 ( .A(n_559), .Y(n_1284) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g1420 ( .A(n_560), .Y(n_1420) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x6_ASAP7_75t_L g967 ( .A(n_562), .B(n_968), .Y(n_967) );
AOI222xp33_ASAP7_75t_L g1362 ( .A1(n_562), .A2(n_1002), .B1(n_1350), .B2(n_1353), .C1(n_1357), .C2(n_1363), .Y(n_1362) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_564), .B(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1170 ( .A(n_564), .Y(n_1170) );
AO22x2_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_654), .B1(n_723), .B2(n_724), .Y(n_565) );
INVx1_ASAP7_75t_L g724 ( .A(n_566), .Y(n_724) );
XNOR2x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_615), .Y(n_568) );
AND4x1_ASAP7_75t_L g569 ( .A(n_570), .B(n_583), .C(n_587), .D(n_591), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B1(n_576), .B2(n_580), .C(n_581), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g1794 ( .A1(n_571), .A2(n_576), .B1(n_581), .B2(n_1795), .C(n_1796), .Y(n_1794) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_883), .C(n_884), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_1065), .C(n_1066), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1259 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_1260), .C(n_1261), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_1411), .C(n_1412), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_1526), .C(n_1527), .Y(n_1525) );
AND2x4_ASAP7_75t_L g1919 ( .A(n_573), .B(n_1920), .Y(n_1919) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g1198 ( .A1(n_578), .A2(n_581), .B(n_1174), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_579), .B(n_970), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_582), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_586), .A2(n_588), .B1(n_631), .B2(n_632), .C(n_634), .Y(n_630) );
AOI33xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .A3(n_603), .B1(n_609), .B2(n_611), .B3(n_614), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g1271 ( .A(n_593), .Y(n_1271) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
BUFx2_ASAP7_75t_L g827 ( .A(n_594), .Y(n_827) );
AND2x4_ASAP7_75t_L g895 ( .A(n_594), .B(n_595), .Y(n_895) );
AND2x2_ASAP7_75t_L g910 ( .A(n_594), .B(n_911), .Y(n_910) );
OR2x2_ASAP7_75t_L g981 ( .A(n_594), .B(n_982), .Y(n_981) );
OR2x6_ASAP7_75t_L g1078 ( .A(n_594), .B(n_1079), .Y(n_1078) );
BUFx2_ASAP7_75t_SL g963 ( .A(n_595), .Y(n_963) );
INVx1_ASAP7_75t_L g1110 ( .A(n_595), .Y(n_1110) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_598), .A2(n_770), .B1(n_771), .B2(n_772), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_598), .A2(n_1152), .B1(n_1153), .B2(n_1154), .Y(n_1151) );
INVx4_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g610 ( .A(n_599), .Y(n_610) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_599), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1807 ( .A(n_599), .Y(n_1807) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g613 ( .A(n_601), .Y(n_613) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g909 ( .A(n_605), .Y(n_909) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g941 ( .A(n_606), .Y(n_941) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g1246 ( .A(n_610), .Y(n_1246) );
INVx2_ASAP7_75t_L g860 ( .A(n_614), .Y(n_860) );
INVx1_ASAP7_75t_L g1030 ( .A(n_614), .Y(n_1030) );
AOI33xp33_ASAP7_75t_L g1535 ( .A1(n_614), .A2(n_1270), .A3(n_1536), .B1(n_1537), .B2(n_1538), .B3(n_1539), .Y(n_1535) );
AOI33xp33_ASAP7_75t_L g1803 ( .A1(n_614), .A2(n_1270), .A3(n_1804), .B1(n_1805), .B2(n_1808), .B3(n_1809), .Y(n_1803) );
AOI31xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_635), .A3(n_649), .B(n_652), .Y(n_617) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_626), .B(n_1000), .Y(n_1137) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g639 ( .A(n_627), .Y(n_639) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_629), .Y(n_665) );
INVx1_ASAP7_75t_L g871 ( .A(n_629), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_631), .A2(n_634), .B1(n_736), .B2(n_738), .C(n_784), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g1396 ( .A1(n_631), .A2(n_1397), .B(n_1398), .C(n_1399), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_632), .A2(n_875), .B1(n_988), .B2(n_989), .C(n_990), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_632), .A2(n_1374), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g1820 ( .A1(n_634), .A2(n_784), .B1(n_1008), .B2(n_1799), .C(n_1801), .Y(n_1820) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g1825 ( .A(n_641), .Y(n_1825) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g1443 ( .A(n_645), .Y(n_1443) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g661 ( .A(n_646), .Y(n_661) );
INVx2_ASAP7_75t_L g793 ( .A(n_646), .Y(n_793) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_646), .Y(n_814) );
INVx1_ASAP7_75t_L g1057 ( .A(n_646), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g1090 ( .A(n_648), .Y(n_1090) );
AOI31xp33_ASAP7_75t_L g775 ( .A1(n_652), .A2(n_776), .A3(n_785), .B(n_795), .Y(n_775) );
INVx1_ASAP7_75t_L g1193 ( .A(n_652), .Y(n_1193) );
AOI31xp33_ASAP7_75t_L g1812 ( .A1(n_652), .A2(n_1813), .A3(n_1821), .B(n_1830), .Y(n_1812) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI31xp33_ASAP7_75t_L g1038 ( .A1(n_653), .A2(n_1039), .A3(n_1045), .B(n_1060), .Y(n_1038) );
INVx3_ASAP7_75t_L g723 ( .A(n_654), .Y(n_723) );
INVx1_ASAP7_75t_L g721 ( .A(n_655), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_685), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_683), .B2(n_684), .Y(n_656) );
INVx2_ASAP7_75t_L g892 ( .A(n_657), .Y(n_892) );
NOR2xp67_ASAP7_75t_L g968 ( .A(n_657), .B(n_969), .Y(n_968) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_673), .C(n_680), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_664), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_659) );
INVx1_ASAP7_75t_L g1301 ( .A(n_662), .Y(n_1301) );
INVx1_ASAP7_75t_L g1295 ( .A(n_663), .Y(n_1295) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_666), .A2(n_817), .B1(n_818), .B2(n_820), .C(n_824), .Y(n_816) );
INVx1_ASAP7_75t_L g881 ( .A(n_666), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_667), .A2(n_682), .B1(n_705), .B2(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g825 ( .A(n_670), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_670), .A2(n_672), .B1(n_883), .B2(n_884), .Y(n_882) );
INVx4_ASAP7_75t_L g1173 ( .A(n_670), .Y(n_1173) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AOI222xp33_ASAP7_75t_SL g1168 ( .A1(n_672), .A2(n_1169), .B1(n_1171), .B2(n_1172), .C1(n_1174), .C2(n_1175), .Y(n_1168) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_677), .A2(n_681), .B1(n_699), .B2(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_678), .A2(n_806), .B1(n_808), .B2(n_809), .C(n_812), .Y(n_805) );
INVx1_ASAP7_75t_L g879 ( .A(n_678), .Y(n_879) );
INVx1_ASAP7_75t_L g1044 ( .A(n_678), .Y(n_1044) );
AOI21xp5_ASAP7_75t_L g1437 ( .A1(n_678), .A2(n_1438), .B(n_1442), .Y(n_1437) );
AOI221xp5_ASAP7_75t_L g1493 ( .A1(n_678), .A2(n_1486), .B1(n_1494), .B2(n_1495), .C(n_1496), .Y(n_1493) );
BUFx3_ASAP7_75t_L g1406 ( .A(n_679), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_684), .A2(n_801), .B1(n_826), .B2(n_828), .Y(n_800) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_694), .C(n_697), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_690), .Y(n_686) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g1344 ( .A(n_700), .Y(n_1344) );
INVx1_ASAP7_75t_L g1471 ( .A(n_700), .Y(n_1471) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_709), .B2(n_711), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_705), .A2(n_1348), .B1(n_1476), .B2(n_1477), .Y(n_1475) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_706), .Y(n_1027) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_707), .Y(n_854) );
INVx1_ASAP7_75t_L g1250 ( .A(n_707), .Y(n_1250) );
INVx2_ASAP7_75t_L g1856 ( .A(n_707), .Y(n_1856) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g715 ( .A(n_710), .Y(n_715) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_710), .Y(n_1018) );
INVx1_ASAP7_75t_L g1115 ( .A(n_710), .Y(n_1115) );
INVx2_ASAP7_75t_L g1428 ( .A(n_710), .Y(n_1428) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g903 ( .A(n_715), .Y(n_903) );
INVx2_ASAP7_75t_L g1482 ( .A(n_715), .Y(n_1482) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_717), .A2(n_843), .B1(n_845), .B2(n_846), .Y(n_842) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x6_ASAP7_75t_L g964 ( .A(n_719), .B(n_946), .Y(n_964) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_719), .B(n_946), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_719), .A2(n_960), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g752 ( .A(n_720), .Y(n_752) );
INVx2_ASAP7_75t_L g1342 ( .A(n_720), .Y(n_1342) );
BUFx2_ASAP7_75t_L g1474 ( .A(n_720), .Y(n_1474) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_922), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_797), .B2(n_921), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
XNOR2x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_796), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_773), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_741), .C(n_745), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B1(n_750), .B2(n_753), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_747), .A2(n_859), .B1(n_1222), .B2(n_1224), .Y(n_1253) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_748), .A2(n_803), .B1(n_808), .B2(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g767 ( .A(n_752), .Y(n_767) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_752), .A2(n_959), .B1(n_960), .B2(n_962), .C(n_963), .Y(n_958) );
AOI21xp33_ASAP7_75t_L g1358 ( .A1(n_752), .A2(n_946), .B(n_1359), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_758), .B1(n_759), .B2(n_763), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_755), .A2(n_1029), .B1(n_1120), .B2(n_1121), .C(n_1122), .Y(n_1119) );
OAI22xp5_ASAP7_75t_SL g1243 ( .A1(n_755), .A2(n_1244), .B1(n_1245), .B2(n_1246), .Y(n_1243) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g765 ( .A(n_756), .Y(n_765) );
INVx1_ASAP7_75t_L g1479 ( .A(n_756), .Y(n_1479) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx3_ASAP7_75t_L g1252 ( .A(n_762), .Y(n_1252) );
INVx2_ASAP7_75t_L g1349 ( .A(n_762), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_767), .A2(n_960), .B1(n_1082), .B2(n_1086), .C(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
BUFx3_ASAP7_75t_L g1185 ( .A(n_782), .Y(n_1185) );
OAI221xp5_ASAP7_75t_L g983 ( .A1(n_784), .A2(n_875), .B1(n_959), .B2(n_962), .C(n_984), .Y(n_983) );
OAI221xp5_ASAP7_75t_L g1867 ( .A1(n_784), .A2(n_1083), .B1(n_1852), .B2(n_1853), .C(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g1088 ( .A(n_788), .Y(n_1088) );
INVx1_ASAP7_75t_L g1512 ( .A(n_788), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_793), .A2(n_1023), .B1(n_1028), .B2(n_1041), .Y(n_1040) );
INVx2_ASAP7_75t_L g921 ( .A(n_797), .Y(n_921) );
XOR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_863), .Y(n_797) );
INVx1_ASAP7_75t_L g861 ( .A(n_799), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_829), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .C(n_816), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_804), .A2(n_817), .B1(n_853), .B2(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_L g1441 ( .A(n_811), .Y(n_1441) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx4_ASAP7_75t_L g1207 ( .A(n_814), .Y(n_1207) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1444 ( .A(n_823), .Y(n_1444) );
CKINVDCx8_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_840), .C(n_841), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_831), .B(n_836), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_831) );
INVx2_ASAP7_75t_L g917 ( .A(n_833), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_835), .Y(n_918) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_835), .Y(n_1036) );
INVx1_ASAP7_75t_L g1035 ( .A(n_839), .Y(n_1035) );
INVx1_ASAP7_75t_L g1149 ( .A(n_839), .Y(n_1149) );
INVx1_ASAP7_75t_L g1383 ( .A(n_839), .Y(n_1383) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_848), .A2(n_1029), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1858 ( .A1(n_850), .A2(n_1856), .B1(n_1859), .B2(n_1860), .Y(n_1858) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g907 ( .A(n_857), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_859), .A2(n_1240), .B1(n_1241), .B2(n_1242), .Y(n_1239) );
INVx1_ASAP7_75t_L g920 ( .A(n_864), .Y(n_920) );
NAND4xp75_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .C(n_893), .D(n_913), .Y(n_864) );
OAI31xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_880), .A3(n_890), .B(n_891), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_868) );
OAI21xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B(n_877), .Y(n_873) );
INVx2_ASAP7_75t_SL g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g887 ( .A(n_876), .Y(n_887) );
INVx1_ASAP7_75t_L g1055 ( .A(n_876), .Y(n_1055) );
BUFx3_ASAP7_75t_L g1210 ( .A(n_878), .Y(n_1210) );
INVx2_ASAP7_75t_L g1218 ( .A(n_878), .Y(n_1218) );
BUFx2_ASAP7_75t_L g1321 ( .A(n_878), .Y(n_1321) );
INVx1_ASAP7_75t_L g1819 ( .A(n_878), .Y(n_1819) );
OAI211xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B(n_888), .C(n_889), .Y(n_885) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
OAI31xp33_ASAP7_75t_SL g1103 ( .A1(n_892), .A2(n_1104), .A3(n_1107), .B(n_1118), .Y(n_1103) );
AOI31xp33_ASAP7_75t_SL g1432 ( .A1(n_892), .A2(n_1433), .A3(n_1437), .B(n_1445), .Y(n_1432) );
AOI31xp33_ASAP7_75t_L g1506 ( .A1(n_892), .A2(n_1507), .A3(n_1515), .B(n_1521), .Y(n_1506) );
AND2x2_ASAP7_75t_SL g893 ( .A(n_894), .B(n_912), .Y(n_893) );
AOI33xp33_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_896), .A3(n_900), .B1(n_904), .B2(n_908), .B3(n_910), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_895), .A2(n_1414), .B1(n_1419), .B2(n_1420), .Y(n_1413) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
AND2x4_ASAP7_75t_L g929 ( .A(n_899), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AND2x4_ASAP7_75t_L g936 ( .A(n_907), .B(n_930), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g1377 ( .A(n_910), .B(n_1378), .C(n_1379), .Y(n_1377) );
INVx1_ASAP7_75t_L g1865 ( .A(n_910), .Y(n_1865) );
INVx2_ASAP7_75t_SL g942 ( .A(n_911), .Y(n_942) );
INVx1_ASAP7_75t_L g1125 ( .A(n_911), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_1069), .B1(n_1138), .B2(n_1139), .Y(n_922) );
INVx1_ASAP7_75t_L g1138 ( .A(n_923), .Y(n_1138) );
XNOR2x1_ASAP7_75t_L g923 ( .A(n_924), .B(n_1011), .Y(n_923) );
INVx1_ASAP7_75t_L g1009 ( .A(n_925), .Y(n_1009) );
NAND4xp25_ASAP7_75t_L g925 ( .A(n_926), .B(n_965), .C(n_972), .D(n_995), .Y(n_925) );
INVx8_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_932) );
INVx3_ASAP7_75t_L g1105 ( .A(n_934), .Y(n_1105) );
INVx3_ASAP7_75t_L g1361 ( .A(n_934), .Y(n_1361) );
INVx3_ASAP7_75t_L g1106 ( .A(n_936), .Y(n_1106) );
INVx3_ASAP7_75t_L g1336 ( .A(n_936), .Y(n_1336) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_940), .B(n_943), .Y(n_937) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_939), .Y(n_1278) );
INVx1_ASAP7_75t_L g1124 ( .A(n_941), .Y(n_1124) );
INVx1_ASAP7_75t_L g1354 ( .A(n_942), .Y(n_1354) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g970 ( .A(n_946), .Y(n_970) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
CKINVDCx11_ASAP7_75t_R g1130 ( .A(n_948), .Y(n_1130) );
CKINVDCx6p67_ASAP7_75t_R g950 ( .A(n_951), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_953), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
BUFx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_L g1161 ( .A(n_954), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1922 ( .A(n_954), .B(n_1923), .Y(n_1922) );
INVx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_967), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_967), .B(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1356 ( .A(n_969), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
NOR3xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_980), .C(n_991), .Y(n_972) );
INVx2_ASAP7_75t_L g1101 ( .A(n_974), .Y(n_1101) );
INVx1_ASAP7_75t_L g1332 ( .A(n_974), .Y(n_1332) );
NAND2x1p5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
INVx2_ASAP7_75t_SL g976 ( .A(n_977), .Y(n_976) );
OR2x6_ASAP7_75t_L g978 ( .A(n_977), .B(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g994 ( .A(n_977), .Y(n_994) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_977), .B(n_979), .Y(n_1102) );
INVx2_ASAP7_75t_L g1330 ( .A(n_978), .Y(n_1330) );
OAI22xp5_ASAP7_75t_SL g980 ( .A1(n_981), .A2(n_983), .B1(n_985), .B2(n_987), .Y(n_980) );
OAI22xp5_ASAP7_75t_SL g1866 ( .A1(n_981), .A2(n_985), .B1(n_1867), .B2(n_1869), .Y(n_1866) );
OAI22xp33_ASAP7_75t_L g1075 ( .A1(n_985), .A2(n_1076), .B1(n_1080), .B2(n_1091), .Y(n_1075) );
INVx1_ASAP7_75t_L g1328 ( .A(n_985), .Y(n_1328) );
INVx4_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_991), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g1329 ( .A1(n_991), .A2(n_1330), .B1(n_1331), .B2(n_1332), .C(n_1333), .Y(n_1329) );
AND2x2_ASAP7_75t_L g991 ( .A(n_992), .B(n_994), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_1001), .B1(n_1002), .B2(n_1003), .C(n_1004), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g1364 ( .A1(n_996), .A2(n_1347), .B1(n_1352), .B2(n_1365), .Y(n_1364) );
AND2x2_ASAP7_75t_L g996 ( .A(n_997), .B(n_999), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_997), .A2(n_1024), .B1(n_1026), .B2(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_998), .Y(n_1291) );
INVx1_ASAP7_75t_L g1439 ( .A(n_998), .Y(n_1439) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_1000), .B(n_1006), .Y(n_1005) );
OR2x6_ASAP7_75t_L g1007 ( .A(n_1000), .B(n_1008), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1000), .B(n_1136), .Y(n_1135) );
CKINVDCx6p67_ASAP7_75t_R g1363 ( .A(n_1005), .Y(n_1363) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1006), .Y(n_1097) );
CKINVDCx6p67_ASAP7_75t_R g1365 ( .A(n_1007), .Y(n_1365) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1008), .Y(n_1094) );
OAI21xp33_ASAP7_75t_L g1389 ( .A1(n_1008), .A2(n_1390), .B(n_1391), .Y(n_1389) );
INVx1_ASAP7_75t_SL g1068 ( .A(n_1012), .Y(n_1068) );
NAND4xp75_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1033), .C(n_1038), .D(n_1064), .Y(n_1012) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI211xp5_ASAP7_75t_L g1054 ( .A1(n_1021), .A2(n_1055), .B(n_1056), .C(n_1058), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B1(n_1028), .B2(n_1029), .Y(n_1025) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
NOR2x1_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1037), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1054), .Y(n_1045) );
OAI211xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1048), .B(n_1051), .C(n_1052), .Y(n_1046) );
OAI221xp5_ASAP7_75t_L g1294 ( .A1(n_1048), .A2(n_1081), .B1(n_1264), .B2(n_1266), .C(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND2xp33_ASAP7_75t_L g1402 ( .A(n_1050), .B(n_1403), .Y(n_1402) );
OAI22xp5_ASAP7_75t_L g1604 ( .A1(n_1067), .A2(n_1559), .B1(n_1567), .B2(n_1605), .Y(n_1604) );
INVxp67_ASAP7_75t_SL g1139 ( .A(n_1069), .Y(n_1139) );
XNOR2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
AND4x1_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1074), .C(n_1103), .D(n_1132), .Y(n_1071) );
NOR3xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1098), .C(n_1099), .Y(n_1074) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_1078), .Y(n_1319) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1079), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B1(n_1083), .B2(n_1086), .C(n_1087), .Y(n_1080) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
BUFx2_ASAP7_75t_L g1322 ( .A(n_1097), .Y(n_1322) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1341 ( .A1(n_1109), .A2(n_1342), .B1(n_1343), .B2(n_1344), .C(n_1345), .Y(n_1341) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_SL g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_1115), .A2(n_1159), .B1(n_1160), .B2(n_1162), .Y(n_1158) );
OAI22xp33_ASAP7_75t_SL g1854 ( .A1(n_1115), .A2(n_1855), .B1(n_1856), .B2(n_1857), .Y(n_1854) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_1127), .A2(n_1129), .B1(n_1130), .B2(n_1131), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1134), .Y(n_1132) );
INVxp67_ASAP7_75t_SL g1540 ( .A(n_1140), .Y(n_1540) );
XNOR2xp5_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1312), .Y(n_1140) );
AO22x2_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1143), .B1(n_1255), .B2(n_1256), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
XNOR2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1199), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1166), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1150), .Y(n_1147) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
AOI21xp5_ASAP7_75t_SL g1166 ( .A1(n_1167), .A2(n_1193), .B(n_1194), .Y(n_1166) );
NAND4xp25_ASAP7_75t_SL g1167 ( .A(n_1168), .B(n_1176), .C(n_1181), .D(n_1183), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_1169), .A2(n_1419), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1180), .Y(n_1211) );
OAI221xp5_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1186), .B1(n_1187), .B2(n_1189), .C(n_1190), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
XNOR2x1_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1254), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1228), .Y(n_1200) );
AOI22xp5_ASAP7_75t_L g1201 ( .A1(n_1202), .A2(n_1203), .B1(n_1226), .B2(n_1227), .Y(n_1201) );
OAI31xp33_ASAP7_75t_SL g1385 ( .A1(n_1202), .A2(n_1386), .A3(n_1387), .B(n_1388), .Y(n_1385) );
AOI22xp5_ASAP7_75t_L g1487 ( .A1(n_1202), .A2(n_1284), .B1(n_1488), .B2(n_1498), .Y(n_1487) );
NAND3xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1215), .C(n_1223), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_1212), .A2(n_1225), .B1(n_1248), .B2(n_1251), .Y(n_1247) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1220), .Y(n_1440) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1220), .Y(n_1885) );
NOR3xp33_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1237), .C(n_1238), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1234), .Y(n_1229) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1371 ( .A1(n_1250), .A2(n_1372), .B1(n_1373), .B2(n_1374), .C(n_1375), .Y(n_1371) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
XOR2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1311), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1283), .Y(n_1257) );
AND4x1_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1262), .C(n_1265), .D(n_1269), .Y(n_1258) );
AOI33xp33_ASAP7_75t_L g1269 ( .A1(n_1270), .A2(n_1272), .A3(n_1277), .B1(n_1280), .B2(n_1281), .B3(n_1282), .Y(n_1269) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
BUFx3_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1285), .B(n_1286), .Y(n_1283) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1293), .Y(n_1307) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1612 ( .A1(n_1311), .A2(n_1558), .B1(n_1565), .B2(n_1613), .Y(n_1612) );
XNOR2xp5_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1452), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
XNOR2xp5_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1366), .Y(n_1314) );
NAND4xp75_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1334), .C(n_1362), .D(n_1364), .Y(n_1316) );
AND2x2_ASAP7_75t_SL g1317 ( .A(n_1318), .B(n_1329), .Y(n_1317) );
AOI33xp33_ASAP7_75t_L g1318 ( .A1(n_1319), .A2(n_1320), .A3(n_1323), .B1(n_1326), .B2(n_1327), .B3(n_1328), .Y(n_1318) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1341), .B1(n_1346), .B2(n_1351), .C(n_1355), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g1861 ( .A1(n_1342), .A2(n_1862), .B1(n_1863), .B2(n_1864), .Y(n_1861) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B(n_1358), .Y(n_1355) );
XNOR2xp5_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1407), .Y(n_1366) );
NAND3xp33_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1381), .C(n_1385), .Y(n_1368) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1380), .Y(n_1369) );
NOR2xp33_ASAP7_75t_SL g1381 ( .A(n_1382), .B(n_1384), .Y(n_1381) );
OAI211xp5_ASAP7_75t_SL g1388 ( .A1(n_1389), .A2(n_1392), .B(n_1396), .C(n_1400), .Y(n_1388) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NAND2xp5_ASAP7_75t_SL g1407 ( .A(n_1408), .B(n_1448), .Y(n_1407) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1409), .Y(n_1450) );
NAND3xp33_ASAP7_75t_SL g1409 ( .A(n_1410), .B(n_1413), .C(n_1421), .Y(n_1409) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1432), .Y(n_1449) );
NAND3xp33_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1450), .C(n_1451), .Y(n_1448) );
AOI22xp5_ASAP7_75t_L g1452 ( .A1(n_1453), .A2(n_1454), .B1(n_1499), .B2(n_1500), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
XNOR2xp5_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1487), .Y(n_1457) );
NOR3xp33_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1466), .C(n_1468), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1463), .Y(n_1459) );
OAI22xp33_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1471), .B1(n_1472), .B2(n_1473), .Y(n_1469) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1480), .B1(n_1481), .B2(n_1483), .Y(n_1478) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
NAND3xp33_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1493), .C(n_1497), .Y(n_1488) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
XNOR2x1_ASAP7_75t_SL g1501 ( .A(n_1502), .B(n_1503), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1504), .B(n_1524), .Y(n_1503) );
BUFx2_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
AND4x1_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1528), .C(n_1532), .D(n_1535), .Y(n_1524) );
OAI221xp5_ASAP7_75t_L g1541 ( .A1(n_1542), .A2(n_1785), .B1(n_1788), .B2(n_1833), .C(n_1838), .Y(n_1541) );
AOI211xp5_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1569), .B(n_1698), .C(n_1752), .Y(n_1542) );
OAI321xp33_ASAP7_75t_L g1698 ( .A1(n_1543), .A2(n_1630), .A3(n_1699), .B1(n_1705), .B2(n_1709), .C(n_1724), .Y(n_1698) );
INVx3_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
AOI211xp5_ASAP7_75t_L g1724 ( .A1(n_1544), .A2(n_1725), .B(n_1739), .C(n_1748), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1544), .B(n_1746), .Y(n_1745) );
INVx3_ASAP7_75t_L g1760 ( .A(n_1544), .Y(n_1760) );
NAND3xp33_ASAP7_75t_L g1766 ( .A(n_1544), .B(n_1603), .C(n_1660), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1778 ( .A(n_1544), .B(n_1779), .Y(n_1778) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_1546), .A2(n_1615), .B1(n_1616), .B2(n_1617), .Y(n_1614) );
INVx2_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
AND2x4_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1550), .Y(n_1547) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1548), .Y(n_1554) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1549), .B(n_1562), .Y(n_1561) );
AND2x4_ASAP7_75t_L g1553 ( .A(n_1550), .B(n_1554), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1550), .B(n_1554), .Y(n_1593) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1551), .Y(n_1562) );
BUFx3_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1553), .Y(n_1615) );
OAI22xp33_ASAP7_75t_L g1555 ( .A1(n_1556), .A2(n_1557), .B1(n_1563), .B2(n_1564), .Y(n_1555) );
BUFx3_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
BUFx6f_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1561), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1567 ( .A(n_1560), .B(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1560), .Y(n_1578) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1561), .Y(n_1577) );
BUFx2_ASAP7_75t_SL g1787 ( .A(n_1564), .Y(n_1787) );
HB1xp67_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1568), .Y(n_1581) );
NAND4xp25_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1648), .C(n_1661), .D(n_1683), .Y(n_1569) );
NOR3xp33_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1635), .C(n_1640), .Y(n_1570) );
OAI211xp5_ASAP7_75t_L g1571 ( .A1(n_1572), .A2(n_1587), .B(n_1606), .C(n_1627), .Y(n_1571) );
OAI221xp5_ASAP7_75t_L g1725 ( .A1(n_1572), .A2(n_1703), .B1(n_1726), .B2(n_1734), .C(n_1735), .Y(n_1725) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1573), .B(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1583), .Y(n_1573) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1574), .Y(n_1608) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1574), .Y(n_1626) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1574), .Y(n_1645) );
OR2x2_ASAP7_75t_L g1658 ( .A(n_1574), .B(n_1584), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1582), .Y(n_1574) );
AND2x4_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1578), .Y(n_1576) );
AND2x4_ASAP7_75t_L g1580 ( .A(n_1578), .B(n_1581), .Y(n_1580) );
BUFx2_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
HB1xp67_ASAP7_75t_L g1928 ( .A(n_1581), .Y(n_1928) );
OR2x2_ASAP7_75t_L g1625 ( .A(n_1583), .B(n_1626), .Y(n_1625) );
AND2x4_ASAP7_75t_L g1630 ( .A(n_1583), .B(n_1610), .Y(n_1630) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1583), .B(n_1611), .Y(n_1693) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1583), .Y(n_1712) );
NOR2xp33_ASAP7_75t_L g1719 ( .A(n_1583), .B(n_1720), .Y(n_1719) );
AOI221xp5_ASAP7_75t_L g1768 ( .A1(n_1583), .A2(n_1769), .B1(n_1771), .B2(n_1773), .C(n_1774), .Y(n_1768) );
INVx3_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1584), .B(n_1610), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1584), .B(n_1611), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1584), .B(n_1645), .Y(n_1674) );
AOI322xp5_ASAP7_75t_L g1683 ( .A1(n_1584), .A2(n_1589), .A3(n_1684), .B1(n_1686), .B2(n_1689), .C1(n_1692), .C2(n_1694), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1585), .B(n_1586), .Y(n_1584) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1594), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1589), .B(n_1633), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1669 ( .A(n_1589), .B(n_1596), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1589), .B(n_1603), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1589), .B(n_1711), .Y(n_1710) );
NOR2xp33_ASAP7_75t_L g1729 ( .A(n_1589), .B(n_1600), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1589), .B(n_1600), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1746 ( .A(n_1589), .B(n_1634), .Y(n_1746) );
BUFx3_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
BUFx2_ASAP7_75t_L g1622 ( .A(n_1590), .Y(n_1622) );
INVxp67_ASAP7_75t_L g1632 ( .A(n_1590), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1590), .B(n_1603), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1590), .B(n_1619), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1599), .Y(n_1594) );
NOR2xp33_ASAP7_75t_L g1639 ( .A(n_1595), .B(n_1620), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1595), .B(n_1630), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1595), .B(n_1619), .Y(n_1711) );
OAI21xp5_ASAP7_75t_SL g1739 ( .A1(n_1595), .A2(n_1740), .B(n_1747), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1595), .B(n_1678), .Y(n_1763) );
INVx2_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1596), .B(n_1608), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1596), .B(n_1622), .Y(n_1621) );
BUFx2_ASAP7_75t_L g1651 ( .A(n_1596), .Y(n_1651) );
INVx2_ASAP7_75t_L g1660 ( .A(n_1596), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1596), .B(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1596), .B(n_1599), .Y(n_1701) );
A2O1A1Ixp33_ASAP7_75t_L g1713 ( .A1(n_1596), .A2(n_1646), .B(n_1714), .C(n_1716), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1596), .B(n_1610), .Y(n_1720) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1596), .B(n_1693), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1770 ( .A(n_1596), .B(n_1715), .Y(n_1770) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1598), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1599), .B(n_1621), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1603), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1600), .B(n_1603), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1600), .B(n_1634), .Y(n_1633) );
INVx2_ASAP7_75t_L g1672 ( .A(n_1600), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1602), .Y(n_1600) );
AOI32xp33_ASAP7_75t_L g1606 ( .A1(n_1603), .A2(n_1607), .A3(n_1609), .B1(n_1618), .B2(n_1623), .Y(n_1606) );
INVx2_ASAP7_75t_SL g1634 ( .A(n_1603), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1603), .B(n_1672), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1608), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1608), .B(n_1693), .Y(n_1692) );
O2A1O1Ixp33_ASAP7_75t_L g1757 ( .A1(n_1608), .A2(n_1672), .B(n_1708), .C(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1609), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1609), .B(n_1723), .Y(n_1722) );
INVx2_ASAP7_75t_SL g1624 ( .A(n_1610), .Y(n_1624) );
HB1xp67_ASAP7_75t_L g1636 ( .A(n_1610), .Y(n_1636) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1610), .Y(n_1664) );
AOI21xp5_ASAP7_75t_L g1726 ( .A1(n_1610), .A2(n_1727), .B(n_1730), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1610), .B(n_1660), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1772 ( .A(n_1610), .B(n_1682), .Y(n_1772) );
OAI32xp33_ASAP7_75t_L g1776 ( .A1(n_1610), .A2(n_1624), .A3(n_1677), .B1(n_1711), .B2(n_1715), .Y(n_1776) );
CKINVDCx5p33_ASAP7_75t_R g1610 ( .A(n_1611), .Y(n_1610) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1612), .B(n_1614), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1618), .B(n_1624), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1621), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1619), .B(n_1632), .Y(n_1665) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_1620), .B(n_1669), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1621), .B(n_1678), .Y(n_1677) );
NOR2xp33_ASAP7_75t_L g1671 ( .A(n_1622), .B(n_1672), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1622), .B(n_1678), .Y(n_1697) );
NOR2x1_ASAP7_75t_L g1738 ( .A(n_1622), .B(n_1634), .Y(n_1738) );
NOR2xp33_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1625), .Y(n_1623) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1624), .Y(n_1654) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1624), .Y(n_1707) );
NOR2xp33_ASAP7_75t_L g1736 ( .A(n_1625), .B(n_1737), .Y(n_1736) );
OAI22xp5_ASAP7_75t_L g1767 ( .A1(n_1625), .A2(n_1653), .B1(n_1679), .B2(n_1731), .Y(n_1767) );
INVxp67_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
A2O1A1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1628), .A2(n_1684), .B(n_1703), .C(n_1717), .Y(n_1747) );
NOR2xp33_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1631), .Y(n_1628) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
AOI22xp5_ASAP7_75t_L g1740 ( .A1(n_1630), .A2(n_1741), .B1(n_1743), .B2(n_1744), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1630), .B(n_1682), .Y(n_1750) );
INVx2_ASAP7_75t_L g1723 ( .A(n_1631), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1633), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1632), .B(n_1639), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1632), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1632), .B(n_1678), .Y(n_1715) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1633), .Y(n_1641) );
NOR2xp33_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1637), .Y(n_1635) );
A2O1A1Ixp33_ASAP7_75t_L g1761 ( .A1(n_1637), .A2(n_1642), .B(n_1762), .C(n_1764), .Y(n_1761) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NOR2xp33_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1642), .Y(n_1640) );
OR2x2_ASAP7_75t_L g1679 ( .A(n_1641), .B(n_1669), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1641), .B(n_1688), .Y(n_1687) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1646), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1644), .Y(n_1779) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1645), .Y(n_1682) );
AOI21xp5_ASAP7_75t_L g1748 ( .A1(n_1646), .A2(n_1749), .B(n_1751), .Y(n_1748) );
CKINVDCx5p33_ASAP7_75t_R g1646 ( .A(n_1647), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1647), .B(n_1651), .Y(n_1650) );
O2A1O1Ixp33_ASAP7_75t_L g1648 ( .A1(n_1649), .A2(n_1652), .B(n_1655), .C(n_1656), .Y(n_1648) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1651), .Y(n_1696) );
NAND2xp5_ASAP7_75t_SL g1728 ( .A(n_1651), .B(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
OR2x2_ASAP7_75t_L g1782 ( .A(n_1654), .B(n_1770), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1655), .B(n_1660), .Y(n_1659) );
NOR2xp33_ASAP7_75t_L g1742 ( .A(n_1655), .B(n_1715), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1659), .Y(n_1656) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1660), .B(n_1671), .Y(n_1670) );
NAND2xp5_ASAP7_75t_L g1775 ( .A(n_1660), .B(n_1693), .Y(n_1775) );
AOI211xp5_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1665), .B(n_1666), .C(n_1675), .Y(n_1661) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1664), .B(n_1674), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1664), .B(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1664), .Y(n_1704) );
OAI22xp5_ASAP7_75t_L g1666 ( .A1(n_1667), .A2(n_1668), .B1(n_1670), .B2(n_1673), .Y(n_1666) );
OAI31xp33_ASAP7_75t_L g1780 ( .A1(n_1674), .A2(n_1710), .A3(n_1781), .B(n_1783), .Y(n_1780) );
AOI21xp33_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1679), .B(n_1680), .Y(n_1675) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1678), .Y(n_1688) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1680), .B(n_1755), .Y(n_1754) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx2_ASAP7_75t_L g1703 ( .A(n_1682), .Y(n_1703) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1697), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_1696), .B(n_1738), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1697), .B(n_1707), .Y(n_1784) );
AOI21xp33_ASAP7_75t_SL g1699 ( .A1(n_1700), .A2(n_1702), .B(n_1704), .Y(n_1699) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1701), .Y(n_1734) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
INVxp67_ASAP7_75t_SL g1705 ( .A(n_1706), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1708), .Y(n_1706) );
AOI211xp5_ASAP7_75t_L g1709 ( .A1(n_1710), .A2(n_1712), .B(n_1713), .C(n_1721), .Y(n_1709) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1710), .Y(n_1751) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1712), .Y(n_1743) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
O2A1O1Ixp33_ASAP7_75t_L g1764 ( .A1(n_1715), .A2(n_1750), .B(n_1765), .C(n_1767), .Y(n_1764) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1719), .Y(n_1716) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVxp67_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1733), .Y(n_1731) );
O2A1O1Ixp33_ASAP7_75t_SL g1774 ( .A1(n_1732), .A2(n_1775), .B(n_1776), .C(n_1777), .Y(n_1774) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
NAND3xp33_ASAP7_75t_L g1752 ( .A(n_1753), .B(n_1768), .C(n_1780), .Y(n_1752) );
O2A1O1Ixp33_ASAP7_75t_L g1753 ( .A1(n_1754), .A2(n_1757), .B(n_1759), .C(n_1761), .Y(n_1753) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
INVx2_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
INVxp67_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVxp67_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
CKINVDCx5p33_ASAP7_75t_R g1785 ( .A(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_SL g1786 ( .A(n_1787), .Y(n_1786) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
HB1xp67_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
NAND2xp5_ASAP7_75t_L g1792 ( .A(n_1793), .B(n_1810), .Y(n_1792) );
AND4x1_ASAP7_75t_L g1793 ( .A(n_1794), .B(n_1797), .C(n_1800), .D(n_1803), .Y(n_1793) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
CKINVDCx14_ASAP7_75t_R g1833 ( .A(n_1834), .Y(n_1833) );
INVx2_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
CKINVDCx5p33_ASAP7_75t_R g1835 ( .A(n_1836), .Y(n_1835) );
OAI21xp5_ASAP7_75t_L g1927 ( .A1(n_1837), .A2(n_1928), .B(n_1929), .Y(n_1927) );
CKINVDCx5p33_ASAP7_75t_R g1839 ( .A(n_1840), .Y(n_1839) );
INVx2_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
INVx2_ASAP7_75t_SL g1844 ( .A(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
NAND3xp33_ASAP7_75t_L g1848 ( .A(n_1849), .B(n_1873), .C(n_1904), .Y(n_1848) );
NOR2xp33_ASAP7_75t_L g1849 ( .A(n_1850), .B(n_1866), .Y(n_1849) );
AOI222xp33_ASAP7_75t_L g1884 ( .A1(n_1864), .A2(n_1885), .B1(n_1886), .B2(n_1890), .C1(n_1891), .C2(n_1892), .Y(n_1884) );
OAI31xp33_ASAP7_75t_SL g1873 ( .A1(n_1874), .A2(n_1883), .A3(n_1896), .B(n_1902), .Y(n_1873) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1877), .Y(n_1895) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1878), .Y(n_1877) );
INVx4_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
NAND2xp5_ASAP7_75t_SL g1883 ( .A(n_1884), .B(n_1893), .Y(n_1883) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1887), .B(n_1888), .Y(n_1886) );
INVx1_ASAP7_75t_SL g1901 ( .A(n_1887), .Y(n_1901) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
AOI22xp5_ASAP7_75t_L g1917 ( .A1(n_1890), .A2(n_1892), .B1(n_1918), .B2(n_1919), .Y(n_1917) );
CKINVDCx8_ASAP7_75t_R g1893 ( .A(n_1894), .Y(n_1893) );
CKINVDCx6p67_ASAP7_75t_R g1897 ( .A(n_1898), .Y(n_1897) );
INVx4_ASAP7_75t_L g1899 ( .A(n_1900), .Y(n_1899) );
OAI31xp33_ASAP7_75t_SL g1904 ( .A1(n_1905), .A2(n_1912), .A3(n_1921), .B(n_1924), .Y(n_1904) );
AND2x4_ASAP7_75t_L g1909 ( .A(n_1907), .B(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g1923 ( .A(n_1907), .Y(n_1923) );
INVx5_ASAP7_75t_SL g1908 ( .A(n_1909), .Y(n_1908) );
INVx1_ASAP7_75t_L g1910 ( .A(n_1911), .Y(n_1910) );
CKINVDCx11_ASAP7_75t_R g1913 ( .A(n_1914), .Y(n_1913) );
INVx1_ASAP7_75t_L g1915 ( .A(n_1916), .Y(n_1915) );
INVxp67_ASAP7_75t_L g1920 ( .A(n_1916), .Y(n_1920) );
CKINVDCx16_ASAP7_75t_R g1924 ( .A(n_1925), .Y(n_1924) );
HB1xp67_ASAP7_75t_L g1926 ( .A(n_1927), .Y(n_1926) );
endmodule