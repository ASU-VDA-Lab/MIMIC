module fake_jpeg_10_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_37),
.B1(n_33),
.B2(n_30),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_42),
.B1(n_30),
.B2(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_32),
.B(n_36),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_4),
.Y(n_69)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_15),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_7),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_6),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_57),
.B(n_8),
.C(n_7),
.D(n_11),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_86),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_84),
.C(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_78),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_97),
.B1(n_87),
.B2(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_95),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_94),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_96),
.B(n_88),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);


endmodule