module real_jpeg_29328_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_0),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_54),
.Y(n_94)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_3),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_109),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_109),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_242)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_5),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_120),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_120),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_120),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_28),
.B1(n_54),
.B2(n_55),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_28),
.B1(n_61),
.B2(n_62),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_114),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_114),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_114),
.Y(n_237)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_111),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_111),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_111),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_11),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_153)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_53)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_14),
.A2(n_37),
.B1(n_54),
.B2(n_55),
.Y(n_133)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_16),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_16),
.A2(n_30),
.B(n_34),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_124),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_16),
.B(n_32),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_16),
.A2(n_61),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_16),
.B(n_61),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_16),
.B(n_76),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_16),
.A2(n_93),
.B1(n_99),
.B2(n_248),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_16),
.A2(n_33),
.B(n_264),
.Y(n_263)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_17),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_22),
.B(n_43),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_24),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_30),
.Y(n_31)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_26),
.A2(n_35),
.B(n_124),
.C(n_125),
.Y(n_123)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_32),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_32),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_29),
.A2(n_32),
.B1(n_110),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_29),
.A2(n_32),
.B1(n_119),
.B2(n_192),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_32),
.Y(n_83)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_68),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_33),
.A2(n_62),
.A3(n_72),
.B1(n_265),
.B2(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_34),
.B(n_124),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_84),
.B(n_337),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_77),
.C(n_79),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_44),
.A2(n_45),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_65),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_46),
.B(n_321),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_48),
.A2(n_81),
.B1(n_83),
.B2(n_172),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_52),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_52),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_52),
.A2(n_65),
.B1(n_315),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_59),
.B1(n_102),
.B2(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_53),
.A2(n_59),
.B1(n_105),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_53),
.A2(n_59),
.B1(n_64),
.B2(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_53),
.A2(n_59),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_53),
.A2(n_59),
.B1(n_223),
.B2(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_53),
.B(n_124),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_53),
.A2(n_59),
.B1(n_190),
.B2(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_54),
.B(n_58),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_54),
.B(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_55),
.A2(n_61),
.A3(n_63),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_61),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_76),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_66),
.A2(n_76),
.B1(n_115),
.B2(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_66),
.A2(n_76),
.B1(n_186),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_66),
.A2(n_74),
.B1(n_76),
.B2(n_313),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_71),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_71),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_67),
.A2(n_71),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_67),
.A2(n_71),
.B1(n_129),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_67),
.A2(n_71),
.B1(n_198),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_72),
.Y(n_274)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_77),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_83),
.B1(n_118),
.B2(n_121),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_81),
.A2(n_83),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_330),
.B(n_336),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_306),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_85)
);

AOI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_156),
.A3(n_178),
.B1(n_300),
.B2(n_305),
.C(n_342),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_88),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_136),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_89),
.B(n_136),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_116),
.C(n_131),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_90),
.B(n_131),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_106),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_107),
.C(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_92),
.B(n_101),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_97),
.B1(n_100),
.B2(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_133),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_93),
.A2(n_148),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_93),
.A2(n_99),
.B1(n_242),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_93),
.A2(n_148),
.B1(n_237),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_94),
.A2(n_98),
.B1(n_127),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_94),
.A2(n_98),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_98),
.Y(n_148)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_103),
.A2(n_142),
.B1(n_145),
.B2(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_116),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_128),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_128),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_122),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_124),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_155),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_149),
.C(n_155),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_142),
.A2(n_145),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_147),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_146),
.A2(n_170),
.B(n_173),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_149),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.CI(n_154),
.CON(n_149),
.SN(n_149)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_157),
.B(n_158),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_176),
.B2(n_177),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_161),
.B(n_167),
.C(n_177),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B(n_166),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_165),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_164),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_166),
.B(n_308),
.C(n_317),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_166),
.B(n_308),
.CI(n_317),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_208),
.C(n_213),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_202),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_180),
.B(n_202),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.C(n_194),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_181),
.B(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_191),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_188),
.C(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_193),
.Y(n_298)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_201),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_196),
.B(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_199),
.B(n_201),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_200),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_209),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_210),
.B(n_211),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_294),
.B(n_299),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_280),
.B(n_293),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_258),
.B(n_279),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_238),
.B(n_257),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_218),
.B(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_245),
.B(n_256),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_240),
.B(n_244),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_250),
.B(n_255),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_260),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_271),
.B1(n_277),
.B2(n_278),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_261)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_270),
.C(n_278),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_268),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_289),
.C(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_318),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_316),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_310),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_312),
.C(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_323),
.C(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_327),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule