module fake_netlist_5_1447_n_1847 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1847);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1847;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_106),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_34),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_88),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_94),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_43),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_44),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_151),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_59),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_65),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_68),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_153),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_95),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_110),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_48),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_132),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_23),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_64),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_54),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_179),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_121),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_12),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_105),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_109),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_7),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_112),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_8),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_75),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_98),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_45),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_83),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_18),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_72),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_56),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_19),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_156),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_130),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_10),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_56),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_60),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_8),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_50),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_49),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_45),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_41),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_17),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_126),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_171),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_26),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_52),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_117),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_101),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_5),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_27),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_22),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_137),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_86),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_178),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_37),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_47),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_152),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_54),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_4),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_25),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_60),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_3),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_28),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_160),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_159),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_166),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_115),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_51),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_4),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_25),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_107),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_46),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_69),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_161),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_19),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_39),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_55),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_31),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_67),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_58),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_46),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_1),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_23),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_49),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_35),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_31),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_118),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_124),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_91),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_37),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_13),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_47),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_84),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_157),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_21),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_29),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_87),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_11),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_53),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_139),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_38),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_34),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_63),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_15),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_74),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_136),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_42),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_59),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_44),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_16),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_53),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_18),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_29),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_51),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_61),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_93),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_182),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_361),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_310),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_327),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_244),
.B(n_0),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_0),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_233),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_251),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_299),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_204),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_253),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_264),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_216),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_288),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_268),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_217),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_237),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_217),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_239),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_236),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_266),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_225),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_270),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_231),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_232),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_238),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_248),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_182),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_194),
.B(n_2),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_199),
.B(n_3),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_252),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_194),
.B(n_9),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_257),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_271),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_272),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_265),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_183),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_258),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_276),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_187),
.B(n_11),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_210),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_278),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_236),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_256),
.B(n_308),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_283),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_229),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_230),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_284),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_240),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_255),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_289),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_265),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_259),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_262),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_263),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_269),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_282),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_195),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_236),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_256),
.B(n_13),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_291),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_267),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_287),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_308),
.B(n_14),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_281),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_286),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_292),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_303),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_207),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_290),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_294),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_297),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_301),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_181),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_378),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_191),
.Y(n_461)
);

CKINVDCx8_ASAP7_75t_R g462 ( 
.A(n_366),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_452),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_181),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_399),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_402),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_403),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_362),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_404),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_372),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_405),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_374),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_383),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_362),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_441),
.B(n_185),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_185),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_374),
.B(n_207),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_370),
.B(n_321),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_411),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_413),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_367),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_419),
.B(n_195),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_396),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_421),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_437),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_371),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_384),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_445),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_446),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_409),
.B(n_226),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_448),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_368),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_449),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_426),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_450),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_376),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_392),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_345),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_533),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_461),
.A2(n_412),
.B1(n_447),
.B2(n_423),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_222),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_525),
.B(n_222),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_480),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_494),
.A2(n_410),
.B1(n_274),
.B2(n_277),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_345),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_462),
.B(n_389),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_519),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_382),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_516),
.B(n_376),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_470),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_365),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_386),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_L g563 ( 
.A(n_457),
.B(n_243),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_525),
.B(n_465),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_457),
.B(n_387),
.C(n_386),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_463),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_489),
.B(n_387),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_480),
.B(n_391),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_489),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_463),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_475),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_500),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_468),
.B(n_261),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_R g577 ( 
.A(n_466),
.B(n_368),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_468),
.B(n_391),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_525),
.B(n_401),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_525),
.B(n_243),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_525),
.B(n_401),
.Y(n_584)
);

BUFx10_ASAP7_75t_L g585 ( 
.A(n_520),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_484),
.Y(n_587)
);

AND3x4_ASAP7_75t_L g588 ( 
.A(n_462),
.B(n_369),
.C(n_410),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_484),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_530),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_460),
.A2(n_423),
.B1(n_314),
.B2(n_300),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_484),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_442),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_488),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_525),
.B(n_243),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_534),
.B(n_394),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_525),
.B(n_243),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_493),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_460),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_506),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_488),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_460),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_491),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_472),
.B(n_415),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_525),
.B(n_415),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_472),
.A2(n_300),
.B1(n_314),
.B2(n_287),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_493),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_491),
.B(n_417),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_488),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_477),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_472),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_492),
.B(n_422),
.C(n_417),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_521),
.B(n_243),
.Y(n_617)
);

NOR2x1p5_ASAP7_75t_L g618 ( 
.A(n_467),
.B(n_422),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_521),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_184),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_190),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_534),
.B(n_397),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_493),
.B(n_193),
.Y(n_624)
);

AO22x2_ASAP7_75t_L g625 ( 
.A1(n_522),
.A2(n_261),
.B1(n_254),
.B2(n_296),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_522),
.B(n_425),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_477),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_462),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_493),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_479),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_479),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_527),
.B(n_428),
.C(n_425),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_490),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_490),
.B(n_197),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_527),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_428),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_502),
.B(n_198),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_527),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_522),
.B(n_431),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_521),
.B(n_431),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_522),
.B(n_434),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_469),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_474),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_471),
.B(n_434),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_529),
.A2(n_330),
.B1(n_334),
.B2(n_349),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_496),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_471),
.B(n_444),
.Y(n_652)
);

AO22x2_ASAP7_75t_L g653 ( 
.A1(n_529),
.A2(n_202),
.B1(n_328),
.B2(n_359),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_531),
.B(n_200),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_496),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_496),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_515),
.B(n_390),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_476),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_507),
.B(n_393),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_531),
.B(n_203),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_509),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_478),
.B(n_444),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_497),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_509),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_478),
.B(n_451),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_481),
.B(n_451),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_481),
.B(n_234),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_482),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_499),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_499),
.B(n_400),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_496),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

NOR2x1p5_ASAP7_75t_L g673 ( 
.A(n_498),
.B(n_211),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_508),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_515),
.B(n_205),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_483),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_512),
.A2(n_305),
.B1(n_336),
.B2(n_343),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_502),
.B(n_208),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_515),
.B(n_273),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_565),
.A2(n_485),
.B(n_483),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_562),
.B(n_503),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_557),
.B(n_510),
.C(n_505),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_661),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_550),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_562),
.B(n_571),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_557),
.B(n_395),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_606),
.B(n_626),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_661),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_664),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_542),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_542),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_554),
.A2(n_398),
.B1(n_341),
.B2(n_220),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_485),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_638),
.B(n_486),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_539),
.B(n_654),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_664),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_550),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_638),
.B(n_641),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_539),
.A2(n_250),
.B1(n_215),
.B2(n_351),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_611),
.B(n_518),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_641),
.B(n_486),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_535),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_646),
.B(n_487),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_550),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_646),
.B(n_487),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_566),
.B(n_528),
.C(n_523),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_600),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_560),
.B(n_186),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_568),
.B(n_495),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_679),
.B(n_538),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_583),
.A2(n_495),
.B(n_246),
.C(n_348),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_569),
.B(n_186),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_538),
.A2(n_526),
.B(n_524),
.C(n_517),
.Y(n_715)
);

BUFx6f_ASAP7_75t_SL g716 ( 
.A(n_658),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_633),
.B(n_192),
.C(n_189),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_563),
.A2(n_526),
.B(n_524),
.C(n_517),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_535),
.B(n_524),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_558),
.B(n_189),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_607),
.B(n_192),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_668),
.B(n_495),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_546),
.B(n_526),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_536),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_658),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_657),
.B(n_211),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_668),
.B(n_509),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_649),
.B(n_196),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_652),
.B(n_196),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_676),
.B(n_224),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_582),
.A2(n_298),
.B1(n_295),
.B2(n_293),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_565),
.A2(n_242),
.B1(n_337),
.B2(n_332),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_608),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_662),
.B(n_206),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_651),
.A2(n_619),
.B(n_540),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_548),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_665),
.B(n_206),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_544),
.B(n_227),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_666),
.A2(n_657),
.B1(n_581),
.B2(n_590),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_555),
.B(n_228),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_637),
.B(n_235),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_605),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_597),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_546),
.B(n_532),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_549),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_640),
.B(n_247),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_546),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_563),
.B(n_249),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_549),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_572),
.B(n_209),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_657),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_532),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_654),
.A2(n_260),
.B1(n_309),
.B2(n_331),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_597),
.B(n_532),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_612),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_551),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_567),
.B(n_213),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_615),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_648),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_639),
.B(n_209),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_551),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_552),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_669),
.B(n_275),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_672),
.B(n_279),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_552),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_556),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_556),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_644),
.A2(n_218),
.B1(n_360),
.B2(n_350),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_574),
.B(n_212),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_674),
.B(n_280),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_212),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_540),
.A2(n_619),
.B(n_541),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_570),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_667),
.B(n_285),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_654),
.A2(n_356),
.B1(n_347),
.B2(n_354),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_586),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_639),
.B(n_218),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_644),
.B(n_587),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_587),
.B(n_496),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_678),
.B(n_219),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_570),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_678),
.B(n_219),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_576),
.B(n_221),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_594),
.B(n_213),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_573),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_573),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_559),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_589),
.B(n_504),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_575),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_654),
.A2(n_316),
.B1(n_504),
.B2(n_513),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_654),
.A2(n_316),
.B1(n_504),
.B2(n_513),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_660),
.A2(n_316),
.B1(n_504),
.B2(n_512),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_589),
.B(n_504),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_578),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_623),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_629),
.B(n_504),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_578),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_614),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_620),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_629),
.B(n_504),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_564),
.B(n_307),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_630),
.B(n_511),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_673),
.A2(n_323),
.B1(n_360),
.B2(n_338),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_564),
.B(n_307),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_591),
.A2(n_323),
.B1(n_313),
.B2(n_315),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_660),
.A2(n_325),
.B1(n_358),
.B2(n_357),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_592),
.B(n_313),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_L g810 ( 
.A1(n_650),
.A2(n_325),
.B1(n_358),
.B2(n_357),
.C(n_355),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_660),
.A2(n_322),
.B1(n_355),
.B2(n_353),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_273),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_541),
.A2(n_315),
.B1(n_333),
.B2(n_326),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_620),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_631),
.B(n_326),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_627),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_634),
.B(n_636),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_670),
.B(n_273),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_592),
.B(n_333),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_632),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_595),
.B(n_62),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_595),
.B(n_338),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_559),
.B(n_350),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_559),
.B(n_473),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_559),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_603),
.B(n_214),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_660),
.A2(n_214),
.B1(n_353),
.B2(n_352),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_658),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_599),
.B(n_473),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_599),
.Y(n_832)
);

INVxp33_ASAP7_75t_L g833 ( 
.A(n_659),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_650),
.A2(n_223),
.B1(n_352),
.B2(n_346),
.C(n_342),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_585),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_684),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_699),
.B(n_670),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_778),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_782),
.A2(n_613),
.B(n_603),
.C(n_545),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_687),
.B(n_537),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_784),
.B(n_577),
.C(n_547),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_690),
.B(n_625),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_693),
.B(n_647),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_585),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_716),
.B(n_647),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_712),
.B(n_625),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_734),
.A2(n_604),
.B(n_610),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_712),
.B(n_625),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_690),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_703),
.A2(n_577),
.B1(n_588),
.B2(n_618),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_826),
.A2(n_613),
.B(n_675),
.C(n_596),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_778),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_700),
.A2(n_609),
.B1(n_677),
.B2(n_653),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_685),
.B(n_663),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_737),
.A2(n_553),
.B(n_610),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_696),
.A2(n_553),
.B(n_610),
.Y(n_856)
);

OAI321xp33_ASAP7_75t_L g857 ( 
.A1(n_692),
.A2(n_677),
.A3(n_609),
.B1(n_594),
.B2(n_653),
.C(n_598),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_694),
.A2(n_702),
.B(n_695),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_696),
.A2(n_553),
.B(n_561),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_698),
.A2(n_660),
.B1(n_635),
.B2(n_653),
.Y(n_860)
);

CKINVDCx10_ASAP7_75t_R g861 ( 
.A(n_716),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_780),
.A2(n_617),
.B(n_621),
.Y(n_862)
);

INVx8_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_720),
.B(n_643),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_686),
.B(n_663),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_703),
.B(n_594),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_715),
.A2(n_645),
.B(n_643),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_704),
.A2(n_599),
.B(n_655),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_707),
.A2(n_319),
.B(n_241),
.C(n_245),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_724),
.B(n_635),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_774),
.A2(n_671),
.B(n_655),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_724),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_717),
.B(n_585),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_L g876 ( 
.A(n_681),
.B(n_340),
.C(n_304),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_746),
.B(n_635),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_741),
.A2(n_710),
.B(n_691),
.C(n_722),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_826),
.A2(n_223),
.B(n_346),
.C(n_304),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_746),
.A2(n_635),
.B1(n_622),
.B2(n_624),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_750),
.A2(n_588),
.B1(n_302),
.B2(n_628),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_711),
.A2(n_671),
.B(n_580),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_723),
.A2(n_580),
.B(n_593),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_753),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_789),
.A2(n_580),
.B(n_593),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_730),
.B(n_635),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_761),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_791),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_761),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_789),
.A2(n_580),
.B(n_593),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_773),
.A2(n_311),
.B(n_312),
.C(n_339),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_832),
.A2(n_593),
.B(n_656),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_736),
.B(n_624),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_832),
.A2(n_656),
.B(n_642),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_749),
.A2(n_656),
.B(n_642),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_745),
.A2(n_342),
.B(n_312),
.C(n_317),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_754),
.B(n_624),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_709),
.B(n_624),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_819),
.B(n_537),
.Y(n_899)
);

AOI22x1_ASAP7_75t_L g900 ( 
.A1(n_709),
.A2(n_757),
.B1(n_735),
.B2(n_744),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_735),
.B(n_624),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_754),
.A2(n_628),
.B1(n_622),
.B2(n_537),
.Y(n_902)
);

NOR2x1p5_ASAP7_75t_SL g903 ( 
.A(n_705),
.B(n_622),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_728),
.A2(n_656),
.B(n_642),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_744),
.B(n_622),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_762),
.B(n_602),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_SL g907 ( 
.A(n_725),
.B(n_622),
.Y(n_907)
);

AO21x1_ASAP7_75t_L g908 ( 
.A1(n_779),
.A2(n_14),
.B(n_16),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_750),
.A2(n_329),
.B1(n_317),
.B2(n_320),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_757),
.B(n_311),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_714),
.B(n_602),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_822),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_781),
.A2(n_473),
.B(n_575),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_752),
.B(n_320),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_790),
.A2(n_473),
.B(n_340),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_756),
.A2(n_339),
.B1(n_329),
.B2(n_322),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_830),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_701),
.B(n_20),
.C(n_21),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_795),
.A2(n_473),
.B(n_97),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_729),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_797),
.A2(n_100),
.B1(n_163),
.B2(n_162),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_718),
.B(n_92),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_776),
.B(n_28),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_822),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_30),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_835),
.B(n_99),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_760),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_927)
);

AO21x2_ASAP7_75t_L g928 ( 
.A1(n_680),
.A2(n_167),
.B(n_102),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_760),
.B(n_812),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_812),
.B(n_32),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_739),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_721),
.B(n_36),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_740),
.B(n_40),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_791),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_725),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_763),
.B(n_113),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_732),
.B(n_103),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_830),
.B(n_822),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_828),
.B(n_708),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_770),
.B(n_119),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_742),
.B(n_40),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_765),
.B(n_766),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_772),
.B(n_42),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_827),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_731),
.A2(n_50),
.B(n_55),
.C(n_57),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_759),
.B(n_57),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_805),
.B(n_66),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_798),
.A2(n_802),
.B(n_818),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_763),
.B(n_73),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_759),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_764),
.B(n_76),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_743),
.A2(n_78),
.B(n_80),
.C(n_82),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_682),
.B(n_123),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_824),
.A2(n_125),
.B(n_133),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_727),
.B(n_134),
.Y(n_956)
);

BUFx4f_ASAP7_75t_L g957 ( 
.A(n_786),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_803),
.B(n_135),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_748),
.A2(n_144),
.B(n_149),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_733),
.A2(n_829),
.B1(n_811),
.B2(n_808),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_764),
.A2(n_158),
.B(n_150),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_807),
.A2(n_154),
.B(n_834),
.C(n_810),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_825),
.A2(n_831),
.B(n_804),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_815),
.B(n_793),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_738),
.A2(n_814),
.B(n_801),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_792),
.A2(n_794),
.B1(n_777),
.B2(n_755),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_738),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_727),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_747),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_747),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_813),
.A2(n_767),
.B1(n_796),
.B2(n_788),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_806),
.B(n_823),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_751),
.A2(n_787),
.B(n_821),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_785),
.A2(n_719),
.B(n_809),
.C(n_820),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_833),
.B(n_783),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_767),
.A2(n_768),
.B1(n_796),
.B2(n_788),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_768),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_683),
.A2(n_688),
.B(n_689),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_751),
.A2(n_787),
.B(n_821),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_769),
.B(n_783),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_758),
.A2(n_799),
.B(n_817),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_758),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_775),
.A2(n_799),
.B(n_817),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_713),
.B(n_816),
.C(n_833),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_775),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_800),
.B(n_814),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_801),
.B(n_683),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_688),
.A2(n_689),
.B(n_697),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_697),
.A2(n_716),
.B1(n_726),
.B2(n_699),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_726),
.Y(n_990)
);

BUFx8_ASAP7_75t_L g991 ( 
.A(n_726),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_684),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_734),
.A2(n_737),
.B(n_619),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_791),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_699),
.A2(n_734),
.B(n_712),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_699),
.A2(n_687),
.B(n_685),
.C(n_560),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_694),
.A2(n_565),
.B(n_695),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_712),
.A2(n_699),
.B1(n_562),
.B2(n_703),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_699),
.B(n_687),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_694),
.A2(n_565),
.B(n_695),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_999),
.B(n_837),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_871),
.B1(n_947),
.B2(n_909),
.C(n_932),
.Y(n_1002)
);

OAI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_841),
.A2(n_850),
.B1(n_998),
.B2(n_951),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_846),
.B(n_848),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_844),
.B(n_899),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_855),
.B(n_847),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_874),
.B(n_929),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_960),
.A2(n_962),
.B(n_995),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_964),
.A2(n_893),
.B(n_886),
.C(n_862),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_975),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_924),
.B(n_867),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_914),
.B(n_854),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_L g1014 ( 
.A1(n_937),
.A2(n_948),
.B(n_858),
.C(n_972),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_863),
.B(n_889),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_939),
.A2(n_984),
.B1(n_960),
.B2(n_906),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_963),
.A2(n_949),
.B(n_870),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_882),
.A2(n_869),
.B(n_965),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_836),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_863),
.B(n_917),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_943),
.A2(n_864),
.B(n_995),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_869),
.A2(n_1000),
.B(n_997),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_973),
.A2(n_981),
.B(n_979),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_865),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_863),
.B(n_912),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_925),
.A2(n_853),
.B(n_878),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_868),
.B(n_938),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_SL g1028 ( 
.A1(n_908),
.A2(n_961),
.B(n_974),
.Y(n_1028)
);

INVx6_ASAP7_75t_SL g1029 ( 
.A(n_868),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_846),
.A2(n_848),
.B1(n_924),
.B2(n_853),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_838),
.B(n_852),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_983),
.A2(n_988),
.B(n_900),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_866),
.B(n_992),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_SL g1034 ( 
.A1(n_961),
.A2(n_842),
.B(n_920),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_872),
.A2(n_877),
.B(n_897),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_887),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_930),
.B(n_923),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_860),
.A2(n_966),
.B1(n_912),
.B2(n_958),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_967),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_980),
.B(n_910),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_967),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_980),
.B(n_910),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_968),
.B(n_875),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_971),
.A2(n_976),
.B(n_987),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_976),
.A2(n_883),
.B(n_904),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_843),
.B(n_940),
.Y(n_1047)
);

BUFx4f_ASAP7_75t_SL g1048 ( 
.A(n_991),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_939),
.B(n_958),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_912),
.B(n_956),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_884),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_945),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_986),
.A2(n_966),
.B(n_849),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_936),
.A2(n_898),
.A3(n_901),
.B(n_905),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_888),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_957),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_990),
.B(n_839),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_931),
.A2(n_913),
.B(n_955),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_950),
.A2(n_952),
.B(n_905),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_994),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_977),
.B(n_944),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_933),
.B(n_942),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_895),
.A2(n_880),
.B(n_894),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_SL g1064 ( 
.A1(n_954),
.A2(n_857),
.B(n_922),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_881),
.B(n_857),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_879),
.A2(n_891),
.B(n_935),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_934),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_892),
.A2(n_885),
.B(n_890),
.Y(n_1068)
);

CKINVDCx6p67_ASAP7_75t_R g1069 ( 
.A(n_861),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_957),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_970),
.A2(n_985),
.B(n_982),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_970),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_982),
.Y(n_1073)
);

AND3x4_ASAP7_75t_L g1074 ( 
.A(n_876),
.B(n_918),
.C(n_941),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_982),
.A2(n_985),
.B(n_926),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_946),
.A2(n_902),
.B(n_989),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_985),
.B(n_840),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_916),
.B(n_945),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_915),
.A2(n_953),
.B(n_927),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_959),
.A2(n_919),
.B(n_921),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_989),
.A2(n_903),
.B(n_907),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_845),
.B1(n_928),
.B2(n_991),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_928),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_899),
.B(n_716),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_841),
.A2(n_686),
.B1(n_557),
.B2(n_562),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_999),
.B(n_837),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_945),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_999),
.B(n_837),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_999),
.B(n_837),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_995),
.A2(n_998),
.B(n_699),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_999),
.B(n_837),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_999),
.B(n_837),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_868),
.B(n_938),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_996),
.A2(n_557),
.B(n_962),
.C(n_699),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_967),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_836),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_870),
.A2(n_882),
.B(n_993),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_995),
.A2(n_998),
.B(n_699),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_995),
.A2(n_998),
.B(n_699),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_964),
.A2(n_699),
.B(n_893),
.C(n_886),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_994),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_SL g1104 ( 
.A1(n_960),
.A2(n_557),
.B(n_881),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_841),
.B(n_693),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_870),
.A2(n_882),
.B(n_993),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_995),
.A2(n_998),
.B(n_699),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_975),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_844),
.B(n_543),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_889),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_994),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_SL g1116 ( 
.A1(n_908),
.A2(n_961),
.B(n_878),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_994),
.Y(n_1117)
);

NOR2xp67_ASAP7_75t_L g1118 ( 
.A(n_841),
.B(n_693),
.Y(n_1118)
);

AND3x4_ASAP7_75t_L g1119 ( 
.A(n_843),
.B(n_682),
.C(n_708),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_SL g1120 ( 
.A1(n_881),
.A2(n_686),
.B(n_867),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_889),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1122)
);

NOR2x1_ASAP7_75t_L g1123 ( 
.A(n_899),
.B(n_830),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_967),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_999),
.B(n_837),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_975),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_999),
.B(n_837),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_995),
.A2(n_998),
.B(n_699),
.Y(n_1129)
);

AO21x1_ASAP7_75t_L g1130 ( 
.A1(n_995),
.A2(n_699),
.B(n_961),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_960),
.A2(n_962),
.B(n_699),
.Y(n_1131)
);

NAND2x1_ASAP7_75t_L g1132 ( 
.A(n_969),
.B(n_789),
.Y(n_1132)
);

AND3x4_ASAP7_75t_L g1133 ( 
.A(n_843),
.B(n_682),
.C(n_708),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_999),
.B(n_837),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_999),
.B(n_837),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_978),
.A2(n_873),
.B(n_859),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_844),
.B(n_543),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_999),
.B(n_837),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1141)
);

NAND2x1_ASAP7_75t_L g1142 ( 
.A(n_969),
.B(n_789),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_862),
.A2(n_851),
.A3(n_976),
.B(n_699),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_993),
.A2(n_737),
.B(n_696),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1019),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_1131),
.A2(n_1009),
.B(n_1130),
.C(n_1096),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1113),
.B(n_1138),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1085),
.B(n_1013),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1002),
.A2(n_1065),
.B1(n_1049),
.B2(n_1074),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1151)
);

BUFx2_ASAP7_75t_SL g1152 ( 
.A(n_1060),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1038),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1024),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1122),
.A2(n_1139),
.B(n_1134),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1067),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1038),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1141),
.A2(n_1144),
.B(n_1021),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1098),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1103),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1016),
.A2(n_1026),
.B1(n_1030),
.B2(n_1003),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1011),
.B(n_1112),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_1115),
.B(n_1117),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1031),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1022),
.A2(n_1009),
.B(n_1028),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1126),
.B(n_1128),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1011),
.B(n_1112),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1120),
.B(n_1135),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1052),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1127),
.B(n_1136),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1140),
.B(n_1092),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1090),
.A2(n_1100),
.B(n_1101),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1114),
.Y(n_1174)
);

OR2x2_ASAP7_75t_SL g1175 ( 
.A(n_1004),
.B(n_1041),
.Y(n_1175)
);

INVx5_ASAP7_75t_SL g1176 ( 
.A(n_1069),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1127),
.B(n_1055),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1029),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1090),
.A2(n_1111),
.B(n_1129),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1036),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1043),
.B(n_1008),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1005),
.B(n_1062),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1037),
.B(n_1104),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1056),
.B(n_1044),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1100),
.A2(n_1129),
.B(n_1101),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1025),
.B(n_1050),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1121),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1033),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1191)
);

BUFx2_ASAP7_75t_SL g1192 ( 
.A(n_1114),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1052),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_1026),
.A2(n_1131),
.B(n_1116),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1025),
.B(n_1050),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_1095),
.B(n_1006),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1102),
.A2(n_1017),
.B(n_1014),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1029),
.Y(n_1198)
);

INVx6_ASAP7_75t_L g1199 ( 
.A(n_1020),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1070),
.B(n_1047),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1039),
.A2(n_1030),
.B1(n_1061),
.B2(n_1045),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1055),
.B(n_1051),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1087),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1039),
.B(n_1045),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1118),
.B(n_1123),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1015),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1048),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1025),
.B(n_1020),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1057),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1078),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1073),
.Y(n_1211)
);

OR2x2_ASAP7_75t_SL g1212 ( 
.A(n_1077),
.B(n_1119),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_SL g1213 ( 
.A(n_1012),
.B(n_1082),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1015),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1015),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1057),
.A2(n_1076),
.B1(n_1133),
.B2(n_1012),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1084),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1066),
.A2(n_1082),
.B1(n_1076),
.B2(n_1020),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1066),
.A2(n_1034),
.B1(n_1079),
.B2(n_1072),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1053),
.C(n_1075),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1087),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_L g1222 ( 
.A(n_1040),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1040),
.B(n_1124),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1110),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1097),
.B(n_1124),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1091),
.A2(n_1108),
.B(n_1137),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1042),
.B(n_1054),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1023),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1081),
.Y(n_1229)
);

CKINVDCx8_ASAP7_75t_R g1230 ( 
.A(n_1064),
.Y(n_1230)
);

BUFx2_ASAP7_75t_SL g1231 ( 
.A(n_1071),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1132),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1018),
.A2(n_1083),
.B(n_1058),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1142),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1054),
.B(n_1143),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1054),
.B(n_1143),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1059),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1109),
.B(n_863),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_1002),
.B1(n_1065),
.B2(n_1085),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1104),
.A2(n_1002),
.B1(n_1065),
.B2(n_1085),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1031),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1011),
.B(n_1112),
.Y(n_1242)
);

INVx3_ASAP7_75t_SL g1243 ( 
.A(n_1115),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1245)
);

AOI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_1085),
.B(n_1016),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1036),
.Y(n_1249)
);

INVx3_ASAP7_75t_SL g1250 ( 
.A(n_1115),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1002),
.A2(n_1065),
.B1(n_557),
.B2(n_784),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_1085),
.B(n_1002),
.C(n_1016),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1001),
.A2(n_1092),
.B1(n_1088),
.B2(n_1089),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1120),
.B(n_686),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1038),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1011),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1104),
.A2(n_1085),
.B(n_1002),
.C(n_1016),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1036),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1007),
.A2(n_696),
.B(n_1106),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1011),
.B(n_1112),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1031),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1011),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1019),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1038),
.B(n_1052),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1011),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1019),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1113),
.B(n_1138),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1038),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1027),
.B(n_1094),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1018),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1001),
.B(n_1088),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1145),
.Y(n_1285)
);

INVx8_ASAP7_75t_L g1286 ( 
.A(n_1188),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1154),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1202),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1156),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

BUFx10_ASAP7_75t_L g1291 ( 
.A(n_1207),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1268),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1226),
.A2(n_1228),
.B(n_1197),
.Y(n_1293)
);

INVx6_ASAP7_75t_L g1294 ( 
.A(n_1188),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1222),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1184),
.B(n_1146),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1151),
.B(n_1167),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1210),
.B(n_1208),
.Y(n_1298)
);

BUFx2_ASAP7_75t_R g1299 ( 
.A(n_1152),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1196),
.A2(n_1234),
.B(n_1233),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1244),
.B(n_1247),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1195),
.Y(n_1302)
);

AO21x2_ASAP7_75t_L g1303 ( 
.A1(n_1224),
.A2(n_1155),
.B(n_1194),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1213),
.A2(n_1257),
.B1(n_1204),
.B2(n_1201),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_SL g1305 ( 
.A(n_1174),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1254),
.A2(n_1213),
.B1(n_1150),
.B2(n_1239),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1243),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1195),
.B(n_1179),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1273),
.Y(n_1310)
);

CKINVDCx16_ASAP7_75t_R g1311 ( 
.A(n_1160),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1241),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1210),
.B(n_1191),
.Y(n_1313)
);

NAND2x1_ASAP7_75t_L g1314 ( 
.A(n_1232),
.B(n_1238),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

INVx8_ASAP7_75t_L g1316 ( 
.A(n_1208),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1171),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1177),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1162),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1238),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1204),
.A2(n_1201),
.B1(n_1169),
.B2(n_1217),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1253),
.B(n_1269),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1250),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1172),
.A2(n_1165),
.B1(n_1284),
.B2(n_1274),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1181),
.Y(n_1325)
);

INVx4_ASAP7_75t_SL g1326 ( 
.A(n_1199),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1168),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1153),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1161),
.A2(n_1246),
.B1(n_1239),
.B2(n_1240),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1260),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1242),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1240),
.A2(n_1149),
.B1(n_1216),
.B2(n_1275),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1264),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1265),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1238),
.B(n_1209),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1179),
.B(n_1187),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1165),
.B(n_1271),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1274),
.A2(n_1284),
.B1(n_1281),
.B2(n_1277),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1194),
.A2(n_1158),
.B(n_1263),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1277),
.A2(n_1281),
.B1(n_1256),
.B2(n_1212),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1256),
.B(n_1255),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1185),
.B(n_1246),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1261),
.A2(n_1218),
.B(n_1180),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1214),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1260),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1267),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1237),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1267),
.Y(n_1349)
);

BUFx12f_ASAP7_75t_L g1350 ( 
.A(n_1215),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1272),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1182),
.B(n_1183),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1175),
.A2(n_1230),
.B1(n_1218),
.B2(n_1272),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1148),
.B(n_1200),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1173),
.A2(n_1186),
.B1(n_1219),
.B2(n_1166),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1189),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1283),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1249),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1187),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1262),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1166),
.A2(n_1248),
.B1(n_1282),
.B2(n_1280),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1245),
.Y(n_1363)
);

AO21x1_ASAP7_75t_L g1364 ( 
.A1(n_1235),
.A2(n_1236),
.B(n_1227),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1245),
.A2(n_1252),
.B1(n_1282),
.B2(n_1280),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1223),
.Y(n_1366)
);

BUFx2_ASAP7_75t_SL g1367 ( 
.A(n_1163),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1248),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1225),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1147),
.A2(n_1232),
.B(n_1225),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1229),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1199),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1153),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1251),
.B(n_1279),
.Y(n_1374)
);

CKINVDCx6p67_ASAP7_75t_R g1375 ( 
.A(n_1192),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1251),
.A2(n_1279),
.B1(n_1252),
.B2(n_1276),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1270),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1258),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1203),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1193),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1178),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1220),
.A2(n_1205),
.B(n_1231),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1157),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1266),
.A2(n_1276),
.B1(n_1206),
.B2(n_1198),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1266),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1259),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1157),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1259),
.B(n_1278),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1221),
.A2(n_1203),
.B(n_1170),
.Y(n_1389)
);

INVx6_ASAP7_75t_L g1390 ( 
.A(n_1221),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1170),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1170),
.A2(n_1176),
.B(n_1099),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1176),
.A2(n_1002),
.B1(n_1161),
.B2(n_1254),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1176),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1156),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1202),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1238),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1161),
.A2(n_1002),
.B1(n_1254),
.B2(n_1246),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1145),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1145),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1188),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1145),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1204),
.B(n_1184),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1161),
.A2(n_1002),
.B1(n_1254),
.B2(n_1246),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1156),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1296),
.B(n_1342),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1329),
.A2(n_1307),
.B(n_1398),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1296),
.B(n_1342),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1320),
.B(n_1335),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1357),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1397),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1335),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1398),
.A2(n_1404),
.B(n_1329),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1330),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1403),
.B(n_1364),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1312),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1348),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1396),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1300),
.A2(n_1370),
.B(n_1314),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1293),
.A2(n_1303),
.B(n_1339),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1371),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1335),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1298),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1392),
.A2(n_1353),
.B(n_1382),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1343),
.B(n_1304),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1355),
.A2(n_1370),
.B(n_1364),
.Y(n_1428)
);

INVx4_ASAP7_75t_SL g1429 ( 
.A(n_1335),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1403),
.B(n_1340),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1320),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1306),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1320),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1382),
.Y(n_1434)
);

AO21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1404),
.A2(n_1362),
.B(n_1355),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1362),
.A2(n_1393),
.B(n_1341),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1382),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1298),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1324),
.A2(n_1338),
.B(n_1310),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1397),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1354),
.B(n_1313),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1358),
.B(n_1366),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1316),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1369),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1352),
.B(n_1297),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1308),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1319),
.B(n_1313),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1318),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1301),
.B(n_1322),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1321),
.A2(n_1332),
.B(n_1337),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1288),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1289),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1285),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1287),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1290),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1317),
.B(n_1331),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1292),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_1368),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1346),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1399),
.A2(n_1402),
.B(n_1400),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1315),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1327),
.B(n_1333),
.Y(n_1462)
);

AO222x2_ASAP7_75t_L g1463 ( 
.A1(n_1336),
.A2(n_1374),
.B1(n_1309),
.B2(n_1299),
.C1(n_1308),
.C2(n_1388),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1347),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1378),
.B(n_1385),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1377),
.A2(n_1386),
.B(n_1380),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1360),
.B(n_1401),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1395),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1378),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1360),
.B(n_1385),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1325),
.B(n_1294),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1389),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1373),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1294),
.Y(n_1475)
);

AO21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1384),
.A2(n_1394),
.B(n_1365),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1405),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1359),
.A2(n_1361),
.B(n_1372),
.Y(n_1478)
);

OAI222xp33_ASAP7_75t_L g1479 ( 
.A1(n_1365),
.A2(n_1376),
.B1(n_1372),
.B2(n_1309),
.C1(n_1363),
.C2(n_1374),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1309),
.B(n_1363),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1294),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1302),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1336),
.B(n_1374),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1336),
.B(n_1302),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1373),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1391),
.A2(n_1376),
.B(n_1383),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1427),
.B(n_1326),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1416),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1427),
.B(n_1326),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1428),
.B(n_1373),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1428),
.B(n_1410),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1415),
.B(n_1356),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1447),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1434),
.B(n_1437),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_L g1496 ( 
.A(n_1407),
.B(n_1328),
.C(n_1387),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1430),
.B(n_1356),
.Y(n_1497)
);

NOR2x1_ASAP7_75t_L g1498 ( 
.A(n_1467),
.B(n_1367),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1429),
.B(n_1326),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1422),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1434),
.B(n_1328),
.Y(n_1501)
);

AND2x4_ASAP7_75t_SL g1502 ( 
.A(n_1411),
.B(n_1323),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_SL g1503 ( 
.A(n_1413),
.B(n_1323),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1430),
.B(n_1375),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_SL g1505 ( 
.A(n_1435),
.B(n_1295),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1407),
.A2(n_1286),
.B1(n_1345),
.B2(n_1350),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1426),
.A2(n_1345),
.B1(n_1350),
.B2(n_1286),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1450),
.A2(n_1295),
.B1(n_1379),
.B2(n_1390),
.C(n_1381),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1426),
.B(n_1381),
.C(n_1286),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1409),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1422),
.B(n_1291),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1406),
.B(n_1291),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1408),
.B(n_1291),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1460),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1460),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1486),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1408),
.B(n_1305),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1460),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1431),
.B(n_1305),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1429),
.B(n_1409),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1431),
.B(n_1433),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1409),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1435),
.A2(n_1476),
.B1(n_1441),
.B2(n_1409),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1431),
.B(n_1433),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1503),
.A2(n_1445),
.B(n_1449),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1494),
.B(n_1448),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1451),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1488),
.B(n_1447),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1488),
.B(n_1414),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1532)
);

AOI21xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1508),
.A2(n_1446),
.B(n_1458),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_1478),
.C(n_1459),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_L g1536 ( 
.A(n_1506),
.B(n_1444),
.C(n_1438),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1523),
.B(n_1473),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1506),
.B(n_1424),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1508),
.A2(n_1438),
.B(n_1424),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1523),
.B(n_1429),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1522),
.B(n_1429),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1522),
.B(n_1429),
.Y(n_1542)
);

OAI221xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1524),
.A2(n_1419),
.B1(n_1452),
.B2(n_1463),
.C(n_1456),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1467),
.Y(n_1544)
);

NAND4xp25_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1465),
.C(n_1462),
.D(n_1464),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1496),
.B(n_1436),
.C(n_1464),
.Y(n_1546)
);

AND4x1_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1472),
.C(n_1485),
.D(n_1474),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1493),
.B(n_1469),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1496),
.B(n_1436),
.C(n_1423),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1477),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1509),
.A2(n_1479),
.B(n_1483),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1498),
.B(n_1436),
.C(n_1423),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1518),
.A2(n_1436),
.B1(n_1476),
.B2(n_1462),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1499),
.A2(n_1483),
.B(n_1425),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1504),
.A2(n_1457),
.B1(n_1453),
.B2(n_1454),
.C(n_1455),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1498),
.B(n_1423),
.C(n_1412),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1461),
.Y(n_1559)
);

NAND2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1499),
.B(n_1411),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1497),
.B(n_1461),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1512),
.B(n_1442),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1525),
.B(n_1425),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1512),
.B(n_1442),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1421),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1418),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_SL g1567 ( 
.A(n_1487),
.B(n_1484),
.C(n_1485),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1519),
.B(n_1423),
.C(n_1412),
.Y(n_1568)
);

OAI221xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1510),
.A2(n_1482),
.B1(n_1481),
.B2(n_1475),
.C(n_1457),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1510),
.A2(n_1439),
.B(n_1466),
.Y(n_1570)
);

OAI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1487),
.A2(n_1482),
.B1(n_1481),
.B2(n_1475),
.C(n_1412),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1510),
.B(n_1421),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1489),
.B(n_1475),
.C(n_1470),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1520),
.A2(n_1480),
.B1(n_1471),
.B2(n_1443),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1517),
.B(n_1486),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1515),
.A2(n_1420),
.B(n_1439),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1489),
.A2(n_1480),
.B1(n_1468),
.B2(n_1443),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1495),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1499),
.A2(n_1480),
.B(n_1440),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1518),
.A2(n_1480),
.B1(n_1468),
.B2(n_1443),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1563),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1565),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1578),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1578),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1575),
.B(n_1517),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1517),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1495),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1575),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1572),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1572),
.B(n_1490),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1556),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1552),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1535),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1541),
.B(n_1490),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1541),
.B(n_1490),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1542),
.B(n_1492),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1535),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1526),
.A2(n_1514),
.B1(n_1513),
.B2(n_1518),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1550),
.B(n_1495),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1537),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1537),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1576),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1559),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1576),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1540),
.B(n_1491),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_R g1611 ( 
.A(n_1567),
.B(n_1499),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1570),
.B(n_1491),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1531),
.B(n_1515),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1579),
.B(n_1515),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1554),
.B(n_1501),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1566),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1553),
.B(n_1516),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1554),
.B(n_1501),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1555),
.B(n_1516),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1560),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1598),
.B(n_1596),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1532),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1595),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1591),
.B(n_1589),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1591),
.B(n_1548),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1602),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1595),
.Y(n_1629)
);

AND3x2_ASAP7_75t_L g1630 ( 
.A(n_1601),
.B(n_1520),
.C(n_1514),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1631)
);

NOR3xp33_ASAP7_75t_L g1632 ( 
.A(n_1619),
.B(n_1543),
.C(n_1534),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1599),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1616),
.B(n_1549),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1616),
.B(n_1527),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1616),
.B(n_1528),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1582),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1598),
.B(n_1521),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.B(n_1596),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1602),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1601),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1603),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1585),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1606),
.B(n_1564),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1582),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1594),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1585),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1606),
.B(n_1529),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1596),
.B(n_1521),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1594),
.B(n_1546),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1585),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1582),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1594),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1653),
.B(n_1593),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1637),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1597),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1657),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1634),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1630),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1632),
.A2(n_1551),
.B1(n_1538),
.B2(n_1536),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1627),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1612),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1651),
.B(n_1597),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1631),
.B(n_1597),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1592),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1635),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1622),
.A2(n_1611),
.B1(n_1545),
.B2(n_1538),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1660),
.B(n_1593),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1584),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1584),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1622),
.A2(n_1611),
.B1(n_1626),
.B2(n_1574),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1627),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1612),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1623),
.A2(n_1533),
.B(n_1600),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1648),
.B(n_1610),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1633),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1584),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1621),
.B(n_1592),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1659),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1623),
.A2(n_1600),
.B(n_1547),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1659),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1621),
.B(n_1619),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1626),
.B(n_1613),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1623),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1656),
.B(n_1609),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1698),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1656),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1685),
.B(n_1625),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1667),
.A2(n_1625),
.B1(n_1568),
.B2(n_1588),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1666),
.B(n_1638),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1668),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1665),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1675),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1676),
.A2(n_1615),
.B1(n_1618),
.B2(n_1619),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1673),
.B(n_1646),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1665),
.A2(n_1615),
.B1(n_1618),
.B2(n_1619),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1673),
.B(n_1674),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1664),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1671),
.B(n_1650),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1701),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1701),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1669),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1669),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1687),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1696),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1696),
.B(n_1646),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1587),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1661),
.B(n_1654),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1687),
.B(n_1557),
.C(n_1539),
.Y(n_1729)
);

NOR2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1674),
.B(n_1615),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1670),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1661),
.B(n_1658),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1670),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1698),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1684),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1682),
.B(n_1587),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1700),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1677),
.Y(n_1739)
);

AOI222xp33_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1617),
.B1(n_1618),
.B2(n_1677),
.C1(n_1505),
.C2(n_1684),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1726),
.A2(n_1698),
.B1(n_1577),
.B2(n_1581),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_L g1742 ( 
.A(n_1713),
.B(n_1698),
.Y(n_1742)
);

AOI31xp33_ASAP7_75t_L g1743 ( 
.A1(n_1725),
.A2(n_1513),
.A3(n_1514),
.B(n_1520),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1725),
.A2(n_1617),
.B(n_1587),
.C(n_1663),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1663),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1718),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1708),
.B(n_1672),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1726),
.A2(n_1689),
.B(n_1688),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1713),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1717),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1729),
.A2(n_1617),
.B1(n_1672),
.B2(n_1678),
.Y(n_1752)
);

AOI211x1_ASAP7_75t_SL g1753 ( 
.A1(n_1707),
.A2(n_1679),
.B(n_1678),
.C(n_1662),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1733),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1711),
.A2(n_1679),
.B(n_1617),
.C(n_1689),
.Y(n_1755)
);

AOI322xp5_ASAP7_75t_L g1756 ( 
.A1(n_1712),
.A2(n_1702),
.A3(n_1699),
.B1(n_1694),
.B2(n_1703),
.C1(n_1590),
.C2(n_1604),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1710),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1703),
.Y(n_1758)
);

AO32x1_ASAP7_75t_L g1759 ( 
.A1(n_1704),
.A2(n_1688),
.A3(n_1691),
.B1(n_1697),
.B2(n_1695),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1721),
.A2(n_1716),
.B1(n_1730),
.B2(n_1738),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1713),
.Y(n_1762)
);

AOI311xp33_ASAP7_75t_L g1763 ( 
.A1(n_1709),
.A2(n_1691),
.A3(n_1633),
.B(n_1639),
.C(n_1641),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1719),
.B(n_1702),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1733),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1749),
.A2(n_1737),
.B1(n_1734),
.B2(n_1704),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1757),
.B(n_1739),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1762),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1757),
.B(n_1714),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1747),
.B(n_1727),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1754),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1749),
.A2(n_1734),
.B(n_1731),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1765),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1745),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1762),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1740),
.B(n_1728),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1750),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1764),
.B(n_1706),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1742),
.Y(n_1779)
);

INVxp33_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1751),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1728),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1706),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.B(n_1694),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1748),
.Y(n_1785)
);

OAI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1780),
.A2(n_1752),
.B1(n_1741),
.B2(n_1743),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1775),
.B(n_1753),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1780),
.A2(n_1743),
.B1(n_1744),
.B2(n_1755),
.Y(n_1788)
);

A2O1A1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1769),
.A2(n_1756),
.B(n_1732),
.C(n_1763),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1776),
.A2(n_1740),
.B1(n_1732),
.B2(n_1715),
.C(n_1735),
.Y(n_1790)
);

AOI311xp33_ASAP7_75t_L g1791 ( 
.A1(n_1774),
.A2(n_1722),
.A3(n_1723),
.B(n_1759),
.C(n_1639),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1776),
.A2(n_1715),
.B(n_1759),
.C(n_1736),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1770),
.B(n_1610),
.Y(n_1794)
);

XNOR2xp5_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1502),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1766),
.A2(n_1759),
.B1(n_1662),
.B2(n_1697),
.C(n_1695),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1779),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_L g1798 ( 
.A1(n_1777),
.A2(n_1681),
.B(n_1662),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1797),
.B(n_1768),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1789),
.B(n_1768),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1786),
.B(n_1771),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1788),
.B(n_1783),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1793),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1787),
.A2(n_1772),
.B(n_1773),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1794),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1795),
.Y(n_1806)
);

NOR2xp67_ASAP7_75t_L g1807 ( 
.A(n_1790),
.B(n_1782),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1792),
.A2(n_1781),
.B(n_1778),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_L g1809 ( 
.A(n_1798),
.B(n_1782),
.C(n_1784),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1796),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1800),
.A2(n_1784),
.B1(n_1791),
.B2(n_1680),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1799),
.B(n_1681),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_L g1813 ( 
.A(n_1802),
.B(n_1571),
.C(n_1681),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1683),
.Y(n_1814)
);

NOR2x1p5_ASAP7_75t_SL g1815 ( 
.A(n_1810),
.B(n_1683),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1692),
.C(n_1683),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1807),
.A2(n_1804),
.B(n_1803),
.C(n_1806),
.Y(n_1817)
);

OAI211xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1804),
.A2(n_1692),
.B(n_1697),
.C(n_1695),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1815),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1814),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1817),
.A2(n_1809),
.B1(n_1805),
.B2(n_1692),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1811),
.A2(n_1699),
.B1(n_1693),
.B2(n_1680),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1812),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1693),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1813),
.B(n_1641),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1818),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1819),
.B(n_1644),
.Y(n_1827)
);

NAND4xp75_ASAP7_75t_L g1828 ( 
.A(n_1821),
.B(n_1513),
.C(n_1614),
.D(n_1638),
.Y(n_1828)
);

NOR2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1820),
.B(n_1620),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1826),
.B(n_1645),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1823),
.B(n_1443),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1825),
.A2(n_1569),
.B1(n_1647),
.B2(n_1605),
.C(n_1607),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1828),
.A2(n_1822),
.B1(n_1824),
.B2(n_1620),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1829),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1830),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1834),
.A2(n_1831),
.B1(n_1827),
.B2(n_1832),
.Y(n_1836)
);

NOR3xp33_ASAP7_75t_L g1837 ( 
.A(n_1836),
.B(n_1835),
.C(n_1833),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1502),
.B(n_1620),
.Y(n_1838)
);

AOI221x1_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1605),
.B1(n_1607),
.B2(n_1608),
.C(n_1620),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1586),
.B1(n_1590),
.B2(n_1582),
.C(n_1583),
.Y(n_1840)
);

OAI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1607),
.B(n_1605),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1840),
.B(n_1583),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1841),
.B(n_1605),
.Y(n_1843)
);

AOI222xp33_ASAP7_75t_L g1844 ( 
.A1(n_1842),
.A2(n_1502),
.B1(n_1505),
.B2(n_1590),
.C1(n_1610),
.C2(n_1583),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1843),
.B1(n_1607),
.B2(n_1608),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1590),
.B1(n_1586),
.B2(n_1583),
.C(n_1604),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1573),
.B(n_1613),
.C(n_1588),
.Y(n_1847)
);


endmodule