module real_jpeg_24051_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_28),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_96),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_1),
.A2(n_25),
.B1(n_184),
.B2(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_64),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_83),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_37),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_2),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_157),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_5),
.A2(n_71),
.B1(n_78),
.B2(n_157),
.Y(n_265)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_7),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_54),
.B1(n_78),
.B2(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_9),
.A2(n_74),
.B1(n_81),
.B2(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_90),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_11),
.A2(n_71),
.B1(n_78),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_118),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_118),
.Y(n_261)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_166),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_166),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_13),
.A2(n_69),
.B1(n_78),
.B2(n_166),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_142),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_20),
.B(n_123),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_105),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_21),
.A2(n_85),
.B1(n_86),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_55),
.B2(n_84),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_22),
.A2(n_56),
.B(n_58),
.Y(n_141)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_24),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_24),
.A2(n_38),
.B1(n_56),
.B2(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_111),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_25),
.A2(n_32),
.B1(n_174),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_35),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_25),
.A2(n_211),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_26),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_26),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_26),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_27),
.B(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_32),
.Y(n_251)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_36),
.B(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_38),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_49),
.B(n_51),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_39),
.A2(n_48),
.B1(n_49),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_39),
.A2(n_48),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_39),
.A2(n_99),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_40),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_40),
.A2(n_100),
.B(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_40),
.A2(n_101),
.B1(n_156),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_40),
.A2(n_101),
.B1(n_165),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_40),
.A2(n_52),
.B(n_100),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_42),
.A2(n_43),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_42),
.B(n_94),
.Y(n_209)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_43),
.A2(n_47),
.B(n_154),
.C(n_159),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_43),
.A2(n_64),
.A3(n_93),
.B1(n_200),
.B2(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_48),
.B(n_154),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_48),
.A2(n_102),
.B(n_115),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_72),
.B(n_76),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_59),
.A2(n_117),
.B(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_59),
.A2(n_60),
.B1(n_117),
.B2(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_60),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_61),
.A2(n_65),
.A3(n_79),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_62),
.B(n_64),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_65),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_65),
.B(n_154),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_83),
.Y(n_119)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_74),
.B(n_154),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_130),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_78),
.A2(n_154),
.B(n_247),
.Y(n_264)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_83),
.A2(n_130),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_83),
.A2(n_130),
.B1(n_265),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_98),
.B(n_104),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_92),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_97),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_91),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_91),
.A2(n_96),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_91),
.A2(n_96),
.B1(n_224),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_91),
.A2(n_261),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_92),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_92),
.B(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_122),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_125),
.B1(n_139),
.B2(n_140),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_105),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_120),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_106),
.A2(n_107),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_108),
.B(n_114),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_109),
.A2(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_110),
.B(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_154),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_116),
.B(n_120),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_141),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_138),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_137),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_136),
.A2(n_201),
.B(n_276),
.Y(n_293)
);

AOI311xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_305),
.A3(n_317),
.B(n_321),
.C(n_322),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_267),
.C(n_300),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_241),
.B(n_266),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_217),
.B(n_240),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_193),
.B(n_216),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_170),
.B(n_192),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_152),
.B1(n_158),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_167),
.C(n_168),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_180),
.B(n_191),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_178),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_190),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_207),
.B1(n_214),
.B2(n_215),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_206),
.C(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_219),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_233),
.B2(n_234),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_236),
.C(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_243),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_258),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_257),
.C(n_258),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_253),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_249),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_268),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_285),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_269),
.B(n_285),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_280),
.C(n_281),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_271),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_281),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_295),
.B2(n_296),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_296),
.C(n_299),
.Y(n_319)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_318),
.B(n_323),
.C(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_314),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_314),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_311),
.CI(n_313),
.CON(n_320),
.SN(n_320)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_320),
.Y(n_328)
);


endmodule