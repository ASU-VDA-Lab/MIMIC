module fake_jpeg_28097_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_19),
.B1(n_17),
.B2(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_16),
.B1(n_13),
.B2(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_31),
.B1(n_17),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_50),
.B1(n_51),
.B2(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_33),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_21),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_17),
.B1(n_22),
.B2(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_12),
.B2(n_16),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_10),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_25),
.Y(n_63)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_10),
.C(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_74),
.B1(n_47),
.B2(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_55),
.B1(n_57),
.B2(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_14),
.B1(n_13),
.B2(n_20),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_73),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_52),
.C(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_87),
.C(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_0),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_102),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_28),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_97),
.B1(n_78),
.B2(n_82),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_81),
.C(n_82),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_85),
.B(n_86),
.C(n_80),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_28),
.B(n_24),
.C(n_29),
.D(n_44),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_34),
.C(n_40),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_78),
.C(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_1),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_1),
.B(n_3),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_97),
.B(n_4),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_54),
.A3(n_24),
.B1(n_18),
.B2(n_28),
.C1(n_72),
.C2(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_99),
.B1(n_95),
.B2(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_4),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_109),
.C(n_83),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_3),
.B(n_4),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_83),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_40),
.C(n_64),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_115),
.C(n_110),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_116),
.B(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_62),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_111),
.B(n_40),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_123),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_24),
.B(n_76),
.C(n_39),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_111),
.B1(n_109),
.B2(n_72),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.C(n_121),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_6),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_7),
.B(n_76),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_130),
.C(n_18),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_39),
.B(n_132),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_39),
.Y(n_134)
);


endmodule