module real_jpeg_6238_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_1),
.B(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_2),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_3),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_4),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_4),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_5),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_5),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_5),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_5),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_5),
.B(n_397),
.Y(n_396)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_7),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_7),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_7),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_8),
.B(n_35),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_164),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_8),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_8),
.B(n_77),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_8),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_8),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_8),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_8),
.B(n_431),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_11),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_11),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_11),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_95),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_13),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_13),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_13),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_14),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_14),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_14),
.B(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_15),
.Y(n_147)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_15),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g431 ( 
.A(n_15),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_183),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_181),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_155),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_19),
.B(n_155),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.C(n_117),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_20),
.B(n_100),
.CI(n_117),
.CON(n_475),
.SN(n_475)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_59),
.B1(n_98),
.B2(n_99),
.Y(n_20)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_41),
.C(n_99),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.C(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_23),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.C(n_30),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_49),
.C(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_24),
.A2(n_30),
.B1(n_71),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_24),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_24),
.A2(n_126),
.B1(n_132),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_24),
.A2(n_132),
.B1(n_383),
.B2(n_384),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_25),
.B(n_143),
.Y(n_142)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_25),
.B(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_28),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_28),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_30),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_30),
.B(n_61),
.C(n_68),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_30),
.B(n_320),
.C(n_324),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_30),
.A2(n_71),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_34),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_36),
.A2(n_37),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_36),
.A2(n_37),
.B1(n_148),
.B2(n_149),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_37),
.B(n_135),
.C(n_148),
.Y(n_134)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_39),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_39),
.Y(n_281)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_40),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_49),
.C(n_54),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_48),
.A2(n_49),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_52),
.Y(n_266)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_53),
.Y(n_386)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_72),
.C(n_84),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_60),
.B(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_68),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_67),
.B(n_103),
.C(n_109),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_67),
.A2(n_68),
.B1(n_126),
.B2(n_296),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_68),
.B(n_126),
.C(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_69),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_70),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_72),
.B(n_84),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_79),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_73),
.A2(n_122),
.B1(n_247),
.B2(n_252),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_73),
.B(n_109),
.C(n_247),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_75),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_76),
.B(n_79),
.Y(n_123)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_78),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_83),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_94),
.B2(n_97),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_93),
.C(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_89),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_89),
.B(n_276),
.C(n_278),
.Y(n_288)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_113),
.B2(n_114),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_115),
.C(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_107),
.Y(n_307)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_109),
.A2(n_112),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_109),
.A2(n_112),
.B1(n_246),
.B2(n_253),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_110),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_111),
.Y(n_373)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_134),
.C(n_152),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_118),
.A2(n_119),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.C(n_129),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_125),
.Y(n_339)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_128),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_129),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_132),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_134),
.B(n_152),
.Y(n_356)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_136),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.C(n_145),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_138),
.B(n_146),
.Y(n_291)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_142),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_155),
.Y(n_480)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.CI(n_158),
.CON(n_155),
.SN(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_169),
.B2(n_180),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_165),
.B(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_174),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_174),
.B(n_220),
.C(n_225),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_473),
.B(n_476),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_349),
.B(n_358),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_333),
.B(n_348),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_310),
.B(n_332),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_188),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_283),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_189),
.B(n_283),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_244),
.C(n_271),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_190),
.B(n_331),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_190),
.Y(n_478)
);

FAx1_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_217),
.CI(n_227),
.CON(n_190),
.SN(n_190)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_191),
.B(n_217),
.C(n_227),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.C(n_210),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_192),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_201),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_197),
.C(n_201),
.Y(n_282)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_204),
.A2(n_210),
.B1(n_211),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_204),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_205),
.B(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_326)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_220),
.A2(n_226),
.B1(n_259),
.B2(n_260),
.Y(n_391)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_235),
.C(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_233),
.B(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_242),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_239),
.Y(n_407)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_240),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_243),
.B(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_243),
.B(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_243),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_271),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.C(n_256),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_245),
.A2(n_254),
.B1(n_255),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_256),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_262),
.C(n_267),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_257),
.A2(n_258),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_262),
.A2(n_263),
.B1(n_267),
.B2(n_268),
.Y(n_461)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_282),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_274),
.C(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_286),
.C(n_309),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_297),
.B1(n_308),
.B2(n_309),
.Y(n_285)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_289),
.C(n_293),
.Y(n_341)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_306),
.C(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_330),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_311),
.B(n_330),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_327),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_312),
.A2(n_313),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_316),
.B(n_327),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_326),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_317),
.B(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_319),
.B(n_326),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_320),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_334),
.B(n_349),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_336),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_350),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_336),
.B(n_350),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_340),
.CI(n_347),
.CON(n_336),
.SN(n_336)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_343),
.C(n_345),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_351),
.B(n_353),
.C(n_355),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

OAI31xp33_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_469),
.A3(n_470),
.B(n_472),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_463),
.B(n_468),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_448),
.B(n_462),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_402),
.B(n_447),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_392),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_363),
.B(n_392),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_381),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_378),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_365),
.B(n_378),
.C(n_381),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.C(n_374),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_367),
.B1(n_369),
.B2(n_370),
.Y(n_394)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_457),
.C(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_401),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_401),
.B1(n_439),
.B2(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_399),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_441),
.B(n_446),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_427),
.B(n_440),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_412),
.B(n_426),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_423),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_423),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_418),
.B(n_422),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_418),
.Y(n_422)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_429),
.B1(n_434),
.B2(n_435),
.Y(n_428)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_422),
.Y(n_434)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_436),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_436),
.Y(n_440)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_429),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_430),
.A2(n_432),
.B(n_434),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B(n_439),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_443),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_450),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_456),
.C(n_459),
.Y(n_464)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_465),
.Y(n_468)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_474),
.B(n_475),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_475),
.Y(n_477)
);


endmodule