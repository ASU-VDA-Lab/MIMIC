module fake_jpeg_26131_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_34),
.B1(n_23),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_34),
.B1(n_29),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_52),
.B1(n_62),
.B2(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_29),
.B1(n_31),
.B2(n_19),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_32),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_41),
.C(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_0),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_77),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_81),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_32),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_97),
.B1(n_50),
.B2(n_33),
.Y(n_123)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_80),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_32),
.Y(n_81)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_41),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_35),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_87),
.B(n_27),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_35),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_46),
.A2(n_21),
.B1(n_20),
.B2(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2x1p5_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_39),
.Y(n_100)
);

AND2x4_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_46),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_48),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_103),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_63),
.Y(n_109)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_116),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_85),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_85),
.B(n_96),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_58),
.C(n_50),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_100),
.C(n_83),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_74),
.B1(n_76),
.B2(n_80),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_87),
.B1(n_86),
.B2(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_136),
.B1(n_122),
.B2(n_127),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_126),
.C(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_83),
.B(n_91),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_144),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_71),
.Y(n_141)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_159),
.B1(n_119),
.B2(n_111),
.Y(n_166)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_71),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_119),
.B(n_117),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_102),
.B(n_95),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_115),
.B(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_1),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_107),
.A2(n_89),
.B1(n_90),
.B2(n_67),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_171),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_180),
.B(n_181),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_185),
.B1(n_16),
.B2(n_4),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_188),
.B1(n_140),
.B2(n_156),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_119),
.B1(n_128),
.B2(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_147),
.B(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_129),
.B1(n_105),
.B2(n_90),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_105),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_67),
.C(n_125),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_125),
.C(n_116),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_68),
.B1(n_79),
.B2(n_125),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_30),
.B(n_24),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_24),
.B(n_27),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_22),
.C(n_68),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_27),
.B1(n_22),
.B2(n_0),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_1),
.Y(n_189)
);

FAx1_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_133),
.CI(n_144),
.CON(n_191),
.SN(n_191)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_192),
.B(n_180),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_137),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_195),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_145),
.B1(n_150),
.B2(n_159),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_201),
.B1(n_212),
.B2(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_135),
.Y(n_198)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_204),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_149),
.B1(n_156),
.B2(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_143),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_174),
.B1(n_185),
.B2(n_172),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_196),
.B1(n_210),
.B2(n_212),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_200),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_199),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_224),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_178),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_162),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_209),
.Y(n_236)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_194),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_193),
.B(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_164),
.C(n_171),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_177),
.C(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_186),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_169),
.B(n_192),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_191),
.B(n_193),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_190),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_182),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.C(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_166),
.C(n_187),
.Y(n_249)
);

OA21x2_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_233),
.B(n_224),
.Y(n_251)
);

OA21x2_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_235),
.B(n_222),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_219),
.B1(n_217),
.B2(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_254),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_229),
.B1(n_216),
.B2(n_220),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_214),
.B(n_236),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_229),
.CI(n_216),
.CON(n_260),
.SN(n_260)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_6),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_255),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_267),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_257),
.B1(n_260),
.B2(n_258),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_266),
.A2(n_252),
.B1(n_259),
.B2(n_12),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_235),
.C(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_6),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_259),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_222),
.C(n_7),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_9),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_267),
.B(n_268),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_282),
.B(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_274),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_284),
.C(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_288),
.B(n_285),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_289),
.B1(n_13),
.B2(n_14),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_10),
.C(n_14),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_15),
.C(n_16),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_15),
.B(n_195),
.Y(n_294)
);


endmodule