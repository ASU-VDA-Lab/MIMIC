module fake_aes_5555_n_10 (n_1, n_2, n_0, n_10);
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_2), .B(n_1), .Y(n_4) );
OA21x2_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_3), .B(n_0), .Y(n_5) );
INVx5_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
OAI22xp33_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_5), .B1(n_3), .B2(n_2), .Y(n_7) );
NAND3xp33_ASAP7_75t_L g8 ( .A(n_7), .B(n_6), .C(n_0), .Y(n_8) );
OA22x2_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_1), .B1(n_2), .B2(n_0), .Y(n_9) );
AOI22xp33_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_1), .B1(n_6), .B2(n_8), .Y(n_10) );
endmodule