module fake_jpeg_17932_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_39),
.C(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_32),
.C(n_35),
.Y(n_55)
);

CKINVDCx12_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_65),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_8),
.B(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_4),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_5),
.Y(n_66)
);

BUFx24_ASAP7_75t_SL g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_7),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_71),
.B(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_12),
.B(n_13),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_14),
.Y(n_77)
);

CKINVDCx10_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_20),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_24),
.C(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_72),
.B1(n_74),
.B2(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_82),
.A3(n_83),
.B1(n_89),
.B2(n_84),
.C1(n_88),
.C2(n_31),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_27),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_30),
.Y(n_96)
);


endmodule