module fake_jpeg_18496_n_290 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_6),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_23),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_50),
.B1(n_62),
.B2(n_37),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_51),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.C(n_43),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_25),
.B(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_22),
.B1(n_44),
.B2(n_18),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_72),
.B1(n_22),
.B2(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_74),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_59),
.B1(n_62),
.B2(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_39),
.B1(n_37),
.B2(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_37),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_44),
.A3(n_38),
.B1(n_34),
.B2(n_30),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_59),
.B(n_52),
.C(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_54),
.C(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_55),
.C(n_59),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_43),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_15),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_70),
.B(n_75),
.Y(n_103)
);

OAI22x1_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_34),
.B1(n_32),
.B2(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_75),
.B1(n_68),
.B2(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_100),
.B1(n_91),
.B2(n_84),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_81),
.B1(n_64),
.B2(n_70),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_108),
.B1(n_115),
.B2(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_27),
.C(n_28),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_64),
.A3(n_74),
.B1(n_72),
.B2(n_58),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_68),
.B1(n_71),
.B2(n_44),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_36),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_99),
.B1(n_97),
.B2(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_99),
.B1(n_85),
.B2(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_57),
.B1(n_66),
.B2(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_136),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_135),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_15),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_91),
.B(n_92),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_134),
.B(n_137),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_89),
.B1(n_92),
.B2(n_84),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_18),
.B(n_13),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_88),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_155),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_148),
.C(n_56),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_88),
.B1(n_73),
.B2(n_66),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_66),
.B1(n_56),
.B2(n_47),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_43),
.C(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_0),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_18),
.B1(n_13),
.B2(n_38),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_17),
.B1(n_56),
.B2(n_15),
.Y(n_171)
);

NOR4xp25_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_13),
.C(n_21),
.D(n_16),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_109),
.B(n_21),
.C(n_16),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_36),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_151),
.A2(n_114),
.B1(n_121),
.B2(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_170),
.B(n_178),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_156),
.B1(n_137),
.B2(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_17),
.Y(n_173)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_28),
.B(n_32),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_141),
.B1(n_142),
.B2(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_9),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_20),
.B1(n_12),
.B2(n_19),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_147),
.B1(n_130),
.B2(n_134),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_150),
.B(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_8),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_133),
.A2(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_128),
.A2(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_176),
.B1(n_172),
.B2(n_180),
.Y(n_211)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_148),
.C(n_144),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_191),
.C(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_189),
.B1(n_194),
.B2(n_156),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_134),
.B1(n_135),
.B2(n_145),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_130),
.C(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_132),
.B1(n_152),
.B2(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_171),
.B1(n_169),
.B2(n_10),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_140),
.C(n_131),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_131),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_170),
.B1(n_179),
.B2(n_174),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_8),
.C(n_11),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_8),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_197),
.C(n_224),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_187),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_163),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_222),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_164),
.C(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_217),
.C(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_181),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_223),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_164),
.C(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_159),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_172),
.C(n_157),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_190),
.B1(n_169),
.B2(n_10),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_201),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_15),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_193),
.B(n_189),
.C(n_184),
.D(n_194),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_7),
.B(n_9),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_232),
.Y(n_247)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_199),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_203),
.B(n_197),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_215),
.B1(n_209),
.B2(n_10),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_245),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_211),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_6),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_208),
.B1(n_217),
.B2(n_220),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_14),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_237),
.C(n_236),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_19),
.B(n_20),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_29),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_4),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_29),
.C(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_29),
.C(n_6),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_5),
.B(n_10),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_263),
.B(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_4),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_4),
.C(n_9),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_247),
.C(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_241),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_270),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_271),
.B(n_272),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_274),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_4),
.C(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_0),
.C(n_1),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_259),
.B(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_278),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_11),
.C2(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_1),
.C(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_275),
.C(n_280),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_285),
.A2(n_282),
.B(n_1),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_1),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_3),
.Y(n_290)
);


endmodule