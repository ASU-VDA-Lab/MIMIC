module fake_jpeg_13009_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_1),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_13),
.B1(n_15),
.B2(n_10),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_35),
.B1(n_43),
.B2(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_13),
.B1(n_12),
.B2(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_10),
.B1(n_27),
.B2(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_17),
.B1(n_21),
.B2(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_50),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_27),
.C(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_3),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_42),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_45),
.B1(n_35),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_64),
.B1(n_51),
.B2(n_49),
.Y(n_67)
);

OAI21x1_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_51),
.B(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_68),
.B1(n_58),
.B2(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_51),
.B1(n_53),
.B2(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_63),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_39),
.C(n_38),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_39),
.B(n_36),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_59),
.B(n_36),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_79),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_58),
.B(n_63),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_67),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_83),
.B(n_5),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_79),
.A3(n_83),
.B1(n_68),
.B2(n_73),
.C1(n_21),
.C2(n_6),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.C(n_85),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_4),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_84),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_6),
.C(n_4),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_5),
.Y(n_93)
);


endmodule