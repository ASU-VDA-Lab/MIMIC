module fake_jpeg_31289_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_12),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_19),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_28),
.B1(n_14),
.B2(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_28),
.B1(n_13),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_15),
.B1(n_14),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_15),
.B1(n_14),
.B2(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_50)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_31),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_31),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_34),
.B(n_37),
.Y(n_54)
);

AO21x1_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_62),
.B(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_61),
.B1(n_51),
.B2(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_33),
.C(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_16),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_73),
.Y(n_89)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_43),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_62),
.C(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_55),
.B1(n_68),
.B2(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_82),
.B1(n_62),
.B2(n_45),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_47),
.B(n_50),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_46),
.B1(n_50),
.B2(n_45),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_54),
.C(n_56),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.C(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_59),
.C(n_64),
.Y(n_85)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_90),
.B1(n_94),
.B2(n_82),
.C(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_78),
.C(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_73),
.B(n_26),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_23),
.A3(n_10),
.B1(n_9),
.B2(n_7),
.C(n_6),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_80),
.C(n_77),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_101),
.B(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_69),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_102),
.B(n_23),
.C(n_22),
.D(n_16),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_71),
.C(n_59),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_71),
.B(n_72),
.C(n_52),
.D(n_27),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_58),
.B1(n_67),
.B2(n_52),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_104),
.B1(n_101),
.B2(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_13),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_102),
.C(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_23),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_105),
.B1(n_39),
.B2(n_36),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_103),
.B(n_11),
.C(n_10),
.D(n_9),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_2),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_117),
.B(n_7),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_40),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_115),
.B(n_6),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_114),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_23),
.B(n_21),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_123),
.C(n_7),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);


endmodule