module fake_jpeg_20134_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_23),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_9),
.B(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_11),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.C(n_18),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_40),
.C(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_50),
.B1(n_43),
.B2(n_37),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_10),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_43),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_19),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_22),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_25),
.C(n_27),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_25),
.C(n_13),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_50),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_19),
.B(n_2),
.C(n_5),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_61),
.C(n_62),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_60),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_60),
.Y(n_68)
);

OAI311xp33_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_25),
.A3(n_46),
.B1(n_6),
.C1(n_4),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_5),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_69),
.Y(n_72)
);


endmodule