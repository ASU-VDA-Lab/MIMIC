module fake_ariane_1466_n_791 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_791);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_791;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_52),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_20),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_19),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_41),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_48),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_25),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_33),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx11_ASAP7_75t_R g179 ( 
.A(n_138),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

INVx4_ASAP7_75t_R g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_39),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_68),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_96),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_146),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_93),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_24),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_69),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_59),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_62),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_36),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_37),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_123),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_9),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_149),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_105),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_118),
.Y(n_219)
);

INVx4_ASAP7_75t_R g220 ( 
.A(n_136),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_54),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_214),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_210),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_0),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_191),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_3),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_179),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_13),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_201),
.B(n_180),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_7),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_169),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_173),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_176),
.A2(n_7),
.B(n_8),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_226),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_185),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_262),
.B(n_261),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_223),
.B1(n_221),
.B2(n_186),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_188),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_257),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_266),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_243),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_244),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_189),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_244),
.B(n_197),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_242),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_248),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_239),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_239),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_229),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_231),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_247),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_249),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_253),
.C(n_246),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_274),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_237),
.Y(n_329)
);

BUFx6f_ASAP7_75t_SL g330 ( 
.A(n_303),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_202),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_237),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_203),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_232),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_232),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_281),
.B(n_241),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_233),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_298),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_306),
.B(n_249),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_307),
.B(n_249),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_288),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_205),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_L g348 ( 
.A(n_278),
.B(n_233),
.C(n_236),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_236),
.Y(n_349)
);

BUFx8_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

BUFx6f_ASAP7_75t_SL g353 ( 
.A(n_275),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_305),
.B(n_240),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_240),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_250),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_276),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_272),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_282),
.B(n_250),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_284),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_300),
.B(n_251),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_256),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_300),
.B(n_251),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_251),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_254),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_297),
.B(n_254),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_290),
.B(n_254),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_268),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_286),
.B(n_206),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_290),
.B(n_225),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_290),
.B(n_207),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_L g379 ( 
.A(n_270),
.B(n_219),
.C(n_212),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_290),
.B(n_234),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_271),
.B(n_268),
.C(n_238),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_286),
.B(n_208),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

O2A1O1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_323),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_386)
);

AND2x6_ASAP7_75t_SL g387 ( 
.A(n_354),
.B(n_10),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_215),
.B1(n_213),
.B2(n_11),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_238),
.B(n_234),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_327),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_321),
.B(n_180),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_346),
.A2(n_352),
.B1(n_356),
.B2(n_353),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_344),
.B(n_180),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_361),
.A2(n_12),
.B1(n_220),
.B2(n_238),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

AND2x6_ASAP7_75t_SL g400 ( 
.A(n_339),
.B(n_12),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_332),
.A2(n_234),
.B(n_15),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_164),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_14),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_336),
.B(n_17),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_325),
.B(n_360),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_379),
.B(n_18),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_337),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_364),
.B(n_26),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_353),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_324),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_361),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_324),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_338),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_348),
.B(n_45),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_322),
.A2(n_46),
.B(n_47),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_359),
.B(n_49),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_378),
.B(n_50),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_322),
.B(n_53),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_55),
.Y(n_434)
);

OR2x6_ASAP7_75t_L g435 ( 
.A(n_358),
.B(n_56),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_320),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_377),
.B(n_63),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

BUFx12f_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

NOR2x1p5_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_162),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_331),
.B(n_64),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_370),
.B(n_347),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_160),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_340),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_365),
.B(n_65),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_368),
.B(n_159),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_330),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_342),
.B(n_67),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_381),
.B(n_71),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_390),
.B(n_330),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_455),
.A2(n_72),
.B(n_74),
.Y(n_459)
);

BUFx8_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_390),
.B(n_75),
.Y(n_461)
);

CKINVDCx8_ASAP7_75t_R g462 ( 
.A(n_423),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_388),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_83),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_405),
.A2(n_84),
.B(n_86),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_431),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_403),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_158),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_418),
.B(n_87),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_88),
.Y(n_471)
);

BUFx4f_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_391),
.A2(n_89),
.B(n_90),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_407),
.A2(n_92),
.B(n_94),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_435),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_95),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_452),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_406),
.Y(n_482)
);

A2O1A1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_444),
.A2(n_97),
.B(n_98),
.C(n_100),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

O2A1O1Ixp5_ASAP7_75t_L g485 ( 
.A1(n_395),
.A2(n_101),
.B(n_102),
.C(n_104),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_435),
.B(n_106),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_107),
.Y(n_487)
);

OA22x2_ASAP7_75t_L g488 ( 
.A1(n_398),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_114),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_406),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_396),
.B(n_115),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_396),
.B(n_116),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_396),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_433),
.A2(n_117),
.B(n_119),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_427),
.B(n_157),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_426),
.A2(n_120),
.B(n_121),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_410),
.A2(n_451),
.B(n_442),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_122),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_406),
.B(n_124),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_387),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_456),
.B(n_445),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_430),
.A2(n_125),
.B(n_126),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_436),
.A2(n_128),
.B(n_130),
.C(n_131),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_415),
.A2(n_132),
.B(n_133),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_134),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_417),
.B(n_135),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_416),
.A2(n_140),
.B(n_143),
.C(n_144),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_439),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_459),
.A2(n_429),
.B(n_438),
.Y(n_515)
);

BUFx4f_ASAP7_75t_L g516 ( 
.A(n_470),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_463),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

INVx5_ASAP7_75t_SL g519 ( 
.A(n_512),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_499),
.A2(n_402),
.B(n_446),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_412),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_465),
.A2(n_481),
.B(n_471),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_495),
.A2(n_454),
.B(n_421),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_487),
.A2(n_432),
.B(n_389),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g525 ( 
.A1(n_464),
.A2(n_425),
.B(n_386),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_408),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_458),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_450),
.B(n_449),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

AOI22x1_ASAP7_75t_L g533 ( 
.A1(n_497),
.A2(n_441),
.B1(n_412),
.B2(n_408),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_420),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_509),
.A2(n_424),
.B(n_417),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_482),
.Y(n_537)
);

OAI21x1_ASAP7_75t_SL g538 ( 
.A1(n_508),
.A2(n_400),
.B(n_151),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_494),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_475),
.A2(n_150),
.B(n_152),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_505),
.B(n_153),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_467),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_466),
.A2(n_154),
.B(n_156),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

BUFx8_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_462),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_501),
.B(n_488),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_474),
.A2(n_485),
.B(n_506),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_493),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_513),
.A2(n_489),
.B(n_496),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_528),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_529),
.Y(n_560)
);

INVx11_ASAP7_75t_L g561 ( 
.A(n_530),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_520),
.A2(n_510),
.B(n_492),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_555),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_515),
.A2(n_491),
.B(n_457),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_552),
.A2(n_486),
.B1(n_504),
.B2(n_478),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_516),
.A2(n_478),
.B1(n_476),
.B2(n_480),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_547),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_527),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_528),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_550),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_558),
.A2(n_536),
.B(n_522),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_469),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_534),
.B(n_483),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_524),
.A2(n_502),
.B(n_526),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_527),
.Y(n_581)
);

AO21x1_ASAP7_75t_SL g582 ( 
.A1(n_516),
.A2(n_544),
.B(n_549),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_550),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_545),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_534),
.A2(n_516),
.B1(n_549),
.B2(n_538),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_547),
.Y(n_586)
);

CKINVDCx12_ASAP7_75t_R g587 ( 
.A(n_530),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_544),
.A2(n_549),
.B1(n_557),
.B2(n_551),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_520),
.A2(n_515),
.B(n_553),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_555),
.B(n_551),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_535),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_528),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_514),
.A2(n_555),
.B1(n_554),
.B2(n_521),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_514),
.A2(n_542),
.B1(n_525),
.B2(n_521),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_558),
.A2(n_523),
.B(n_531),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_519),
.B(n_556),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_519),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_528),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_540),
.B(n_556),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_576),
.Y(n_602)
);

NOR2x1_ASAP7_75t_SL g603 ( 
.A(n_582),
.B(n_540),
.Y(n_603)
);

INVx3_ASAP7_75t_SL g604 ( 
.A(n_575),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_578),
.B(n_519),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_579),
.A2(n_556),
.B1(n_519),
.B2(n_533),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_567),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_543),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_R g609 ( 
.A(n_598),
.B(n_541),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_562),
.B(n_543),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_581),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_533),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_570),
.B(n_548),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_562),
.B(n_548),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_540),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_591),
.B(n_538),
.Y(n_620)
);

AO31x2_ASAP7_75t_L g621 ( 
.A1(n_597),
.A2(n_525),
.A3(n_558),
.B(n_536),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_537),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_561),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_574),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_580),
.B(n_537),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_584),
.B(n_569),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_600),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_591),
.B(n_537),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_601),
.B(n_548),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_584),
.B(n_541),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_569),
.B(n_541),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_587),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_597),
.A2(n_546),
.B(n_553),
.Y(n_635)
);

AO31x2_ASAP7_75t_L g636 ( 
.A1(n_595),
.A2(n_536),
.A3(n_523),
.B(n_531),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_SL g637 ( 
.A(n_585),
.B(n_523),
.C(n_541),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_594),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_583),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_R g640 ( 
.A(n_599),
.B(n_546),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_580),
.B(n_531),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_565),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_566),
.B(n_571),
.Y(n_643)
);

INVxp33_ASAP7_75t_SL g644 ( 
.A(n_583),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_573),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_SL g646 ( 
.A(n_564),
.B(n_601),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_559),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_588),
.A2(n_570),
.B1(n_593),
.B2(n_573),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_626),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_610),
.B(n_576),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_622),
.B(n_593),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_628),
.A2(n_559),
.B1(n_589),
.B2(n_563),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_589),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_607),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_589),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_620),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_619),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_590),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_614),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_643),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_641),
.B(n_610),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_616),
.Y(n_663)
);

OA21x2_ASAP7_75t_L g664 ( 
.A1(n_642),
.A2(n_602),
.B(n_627),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_629),
.Y(n_665)
);

INVx4_ASAP7_75t_R g666 ( 
.A(n_618),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_621),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_611),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_621),
.B(n_627),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_620),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_621),
.B(n_645),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_636),
.B(n_605),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_612),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_630),
.B(n_624),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_624),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_649),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_647),
.B(n_617),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_649),
.Y(n_679)
);

AO21x1_ASAP7_75t_SL g680 ( 
.A1(n_613),
.A2(n_609),
.B(n_620),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_608),
.B(n_637),
.Y(n_681)
);

AO21x2_ASAP7_75t_L g682 ( 
.A1(n_637),
.A2(n_615),
.B(n_606),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_608),
.B(n_647),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_650),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_677),
.B(n_604),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_655),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_660),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_678),
.B(n_648),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_654),
.B(n_635),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_676),
.B(n_606),
.C(n_646),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_677),
.B(n_623),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_654),
.B(n_623),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_662),
.B(n_631),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_673),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_661),
.B(n_639),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_656),
.B(n_635),
.C(n_634),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_673),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_674),
.B(n_603),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_667),
.Y(n_701)
);

NAND2x1_ASAP7_75t_SL g702 ( 
.A(n_670),
.B(n_644),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_668),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_667),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_675),
.Y(n_705)
);

BUFx2_ASAP7_75t_SL g706 ( 
.A(n_678),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_664),
.Y(n_707)
);

OAI221xp5_ASAP7_75t_SL g708 ( 
.A1(n_679),
.A2(n_625),
.B1(n_681),
.B2(n_663),
.C(n_669),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_662),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_689),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_685),
.B(n_674),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_669),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_701),
.B(n_663),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_686),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_696),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_687),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_688),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_684),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_693),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_696),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_703),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_707),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_703),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_709),
.B(n_680),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_701),
.B(n_651),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_699),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_689),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_680),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_671),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_704),
.B(n_651),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_694),
.B(n_659),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_712),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_712),
.B(n_698),
.C(n_691),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_714),
.Y(n_734)
);

XNOR2x2_ASAP7_75t_L g735 ( 
.A(n_729),
.B(n_681),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_719),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_L g737 ( 
.A1(n_722),
.A2(n_690),
.B(n_691),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_713),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_711),
.B(n_706),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_729),
.B(n_690),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_725),
.A2(n_670),
.B1(n_657),
.B2(n_695),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_722),
.B(n_707),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_SL g743 ( 
.A(n_727),
.B(n_657),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_738),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_733),
.A2(n_730),
.B1(n_670),
.B2(n_657),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_737),
.A2(n_708),
.B1(n_736),
.B2(n_727),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_742),
.A2(n_718),
.B(n_717),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_734),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_744),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_748),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_747),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_746),
.Y(n_752)
);

NOR3x1_ASAP7_75t_L g753 ( 
.A(n_750),
.B(n_710),
.C(n_742),
.Y(n_753)
);

NOR3x1_ASAP7_75t_L g754 ( 
.A(n_750),
.B(n_740),
.C(n_732),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_751),
.B(n_716),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_756),
.Y(n_757)
);

NOR2x1p5_ASAP7_75t_L g758 ( 
.A(n_755),
.B(n_727),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_753),
.A2(n_752),
.B(n_735),
.C(n_724),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_757),
.B(n_745),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_758),
.A2(n_682),
.B1(n_741),
.B2(n_754),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_759),
.B(n_697),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_758),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_739),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_763),
.Y(n_766)
);

NOR2x1_ASAP7_75t_L g767 ( 
.A(n_761),
.B(n_666),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_682),
.B1(n_728),
.B2(n_672),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_766),
.B(n_765),
.Y(n_769)
);

NOR5xp2_ASAP7_75t_L g770 ( 
.A(n_764),
.B(n_702),
.C(n_743),
.D(n_723),
.E(n_721),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_768),
.B(n_731),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_767),
.B(n_700),
.Y(n_772)
);

OR5x1_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_652),
.C(n_653),
.D(n_682),
.E(n_659),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_765),
.Y(n_774)
);

XOR2xp5_ASAP7_75t_L g775 ( 
.A(n_769),
.B(n_683),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_774),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_770),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_772),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_776),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_777),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

OAI31xp33_ASAP7_75t_SL g783 ( 
.A1(n_781),
.A2(n_782),
.A3(n_780),
.B(n_779),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_779),
.Y(n_784)
);

AOI31xp33_ASAP7_75t_L g785 ( 
.A1(n_779),
.A2(n_773),
.A3(n_771),
.B(n_652),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_784),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_786),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_787),
.B(n_783),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_785),
.B1(n_672),
.B2(n_671),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_789),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_790),
.A2(n_726),
.B1(n_720),
.B2(n_715),
.Y(n_791)
);


endmodule