module fake_jpeg_10400_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_35),
.B(n_45),
.CON(n_67),
.SN(n_67)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_16),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B(n_17),
.C(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_47),
.B(n_63),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_64),
.B1(n_23),
.B2(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_18),
.B1(n_26),
.B2(n_17),
.Y(n_90)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_81),
.B1(n_60),
.B2(n_46),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_45),
.B1(n_35),
.B2(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_38),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_19),
.C(n_37),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_93),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_58),
.B1(n_32),
.B2(n_22),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_19),
.B1(n_17),
.B2(n_38),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_68),
.B1(n_49),
.B2(n_61),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_97),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_43),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_19),
.B(n_17),
.C(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_106),
.B(n_110),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_109),
.Y(n_148)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_37),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_78),
.C(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_54),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

AO21x1_ASAP7_75t_SL g153 ( 
.A1(n_113),
.A2(n_118),
.B(n_22),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_119),
.B1(n_124),
.B2(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_88),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_9),
.Y(n_142)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_46),
.B(n_57),
.C(n_27),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_18),
.B1(n_34),
.B2(n_78),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_60),
.B1(n_18),
.B2(n_43),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_20),
.B1(n_77),
.B2(n_25),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_81),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_132),
.C(n_137),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_142),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_153),
.B1(n_32),
.B2(n_22),
.Y(n_180)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_50),
.B(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_108),
.B1(n_124),
.B2(n_104),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_97),
.C(n_80),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_37),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_147),
.C(n_118),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_139),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_18),
.B1(n_34),
.B2(n_95),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_87),
.B(n_27),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_151),
.B(n_102),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_87),
.C(n_44),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_125),
.Y(n_158)
);

OR2x6_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_18),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_164),
.B1(n_152),
.B2(n_143),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_177),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_156),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_178),
.B(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_163),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_119),
.B1(n_110),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_161),
.A2(n_167),
.B1(n_170),
.B2(n_32),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_153),
.B1(n_135),
.B2(n_136),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_175),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_114),
.B1(n_118),
.B2(n_95),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_169),
.C(n_171),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_105),
.B1(n_120),
.B2(n_109),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_107),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_116),
.B1(n_77),
.B2(n_84),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_107),
.C(n_22),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_31),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_50),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_70),
.C(n_66),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_34),
.B1(n_84),
.B2(n_86),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_152),
.B1(n_141),
.B2(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_183),
.B(n_32),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_149),
.B(n_146),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_186),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_135),
.B(n_134),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_143),
.C(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_198),
.B1(n_201),
.B2(n_181),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_130),
.B(n_140),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_200),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_129),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_202),
.C(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_205),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_164),
.B1(n_179),
.B2(n_160),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_141),
.B(n_139),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_33),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_33),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_55),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_219),
.B1(n_231),
.B2(n_14),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_221),
.B(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_165),
.B1(n_171),
.B2(n_66),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_201),
.B(n_186),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_48),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_225),
.C(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_55),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_185),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_232),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_189),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_29),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_25),
.C(n_1),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.C(n_184),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_16),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_202),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_245),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_200),
.B(n_208),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_0),
.B(n_2),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_244),
.B1(n_234),
.B2(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_206),
.B1(n_182),
.B2(n_197),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_207),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_190),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.C(n_253),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_204),
.B1(n_196),
.B2(n_199),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_252),
.B(n_255),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_210),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_196),
.B1(n_183),
.B2(n_195),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_257),
.B1(n_231),
.B2(n_224),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_182),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_183),
.C(n_1),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_214),
.B(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_15),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_14),
.C(n_12),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_264),
.B1(n_273),
.B2(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_240),
.A2(n_225),
.B1(n_223),
.B2(n_235),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_9),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_0),
.C(n_2),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_270),
.C(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_276),
.B(n_237),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_245),
.C(n_236),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_272),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_9),
.B(n_11),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_284),
.C(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_260),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_254),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_250),
.B(n_253),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_291),
.B(n_267),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_249),
.C(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_262),
.B1(n_276),
.B2(n_259),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_304),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_259),
.B1(n_274),
.B2(n_264),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_289),
.B1(n_284),
.B2(n_277),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_296),
.A2(n_285),
.B(n_288),
.C(n_8),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_266),
.B(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_263),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_263),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_291),
.B(n_280),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_5),
.B(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_304),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_313),
.B(n_306),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_281),
.B1(n_285),
.B2(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_312),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_6),
.B(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_298),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_316),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_300),
.B1(n_303),
.B2(n_295),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_321),
.B(n_323),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_320),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_7),
.C(n_8),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_312),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_324),
.A2(n_307),
.B(n_322),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.C(n_326),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_325),
.A3(n_328),
.B1(n_318),
.B2(n_7),
.C(n_8),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_7),
.Y(n_334)
);


endmodule