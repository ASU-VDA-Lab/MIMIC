module fake_jpeg_30268_n_446 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_446);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_2),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_62),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_7),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_20),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_8),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_90),
.Y(n_101)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_8),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_35),
.B1(n_30),
.B2(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_142),
.B1(n_43),
.B2(n_23),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_26),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_26),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_47),
.A2(n_41),
.B1(n_34),
.B2(n_27),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_19),
.B1(n_23),
.B2(n_39),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_34),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_18),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_18),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_48),
.B(n_45),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_144),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_51),
.A2(n_35),
.B1(n_39),
.B2(n_19),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_56),
.B(n_44),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_71),
.B1(n_70),
.B2(n_30),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_149),
.B1(n_174),
.B2(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_148),
.B(n_162),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_42),
.B1(n_32),
.B2(n_30),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_150),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_19),
.B(n_39),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_184),
.B(n_120),
.Y(n_201)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_139),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_165),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_111),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_168),
.A2(n_118),
.B1(n_98),
.B2(n_136),
.Y(n_204)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_101),
.A2(n_90),
.B1(n_89),
.B2(n_64),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_84),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_183),
.Y(n_193)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_119),
.A2(n_60),
.B1(n_77),
.B2(n_75),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_123),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_23),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_188),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_97),
.A2(n_42),
.B(n_32),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_118),
.C(n_43),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_131),
.A2(n_67),
.B1(n_92),
.B2(n_43),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_105),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_114),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_94),
.B1(n_136),
.B2(n_114),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_190),
.A2(n_204),
.B1(n_153),
.B2(n_165),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_134),
.C(n_138),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_134),
.C(n_138),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_113),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_150),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_162),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_161),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_128),
.B(n_119),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_189),
.B(n_166),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_146),
.B1(n_108),
.B2(n_132),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_108),
.B1(n_146),
.B2(n_102),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_229),
.B1(n_231),
.B2(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_156),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_242),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_170),
.B1(n_188),
.B2(n_102),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_208),
.B1(n_204),
.B2(n_210),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_221),
.B(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_253),
.B1(n_189),
.B2(n_211),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_237),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_170),
.B1(n_188),
.B2(n_173),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_110),
.B1(n_107),
.B2(n_128),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_248),
.Y(n_266)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_222),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_160),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_155),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_193),
.A2(n_110),
.B1(n_132),
.B2(n_107),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_260),
.A2(n_278),
.B1(n_237),
.B2(n_269),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_193),
.B(n_200),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_264),
.B(n_269),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_203),
.C(n_202),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_242),
.C(n_227),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_221),
.B1(n_209),
.B2(n_199),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_198),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_196),
.B1(n_216),
.B2(n_198),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_282),
.B(n_296),
.Y(n_317)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_231),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_288),
.Y(n_319)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_284),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_259),
.B1(n_270),
.B2(n_206),
.Y(n_333)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_293),
.C(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_229),
.B1(n_234),
.B2(n_225),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_292),
.A2(n_297),
.B1(n_279),
.B2(n_254),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_230),
.C(n_228),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_230),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_239),
.C(n_253),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_243),
.B1(n_238),
.B2(n_241),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_262),
.C(n_256),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_216),
.C(n_196),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_303),
.C(n_308),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_280),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_191),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_223),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_275),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_226),
.B1(n_244),
.B2(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_223),
.C(n_191),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_278),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_296),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_266),
.B(n_260),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_320),
.A2(n_330),
.B1(n_335),
.B2(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_288),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_325),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_268),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_323),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_258),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_254),
.C(n_258),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_318),
.C(n_317),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_328),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_301),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_268),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_297),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_292),
.A2(n_259),
.B1(n_270),
.B2(n_276),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_334),
.Y(n_345)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_220),
.B1(n_212),
.B2(n_214),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_338),
.B(n_343),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_355),
.C(n_357),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_291),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_340),
.B(n_312),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_319),
.B(n_291),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_307),
.C(n_306),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_348),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_286),
.B1(n_294),
.B2(n_284),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_349),
.B(n_351),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_352),
.B(n_354),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_212),
.B1(n_169),
.B2(n_214),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_309),
.C(n_326),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_330),
.A2(n_177),
.B1(n_176),
.B2(n_158),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_356),
.B(n_333),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_206),
.C(n_219),
.Y(n_357)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_10),
.C(n_3),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_358),
.A2(n_329),
.B1(n_314),
.B2(n_322),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_372),
.B1(n_374),
.B2(n_10),
.Y(n_389)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_342),
.A2(n_335),
.B(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_365),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_331),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_367),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_324),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_324),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_377),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_219),
.C(n_186),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_375),
.C(n_357),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_152),
.B1(n_181),
.B2(n_184),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_137),
.C(n_63),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_157),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_376),
.B(n_37),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_337),
.A2(n_137),
.B(n_2),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_388),
.Y(n_404)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_341),
.B(n_353),
.C(n_347),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_359),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_360),
.A2(n_348),
.B(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_354),
.C(n_356),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_386),
.C(n_387),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_38),
.C(n_42),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_38),
.C(n_32),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_32),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_393),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_37),
.C(n_0),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_367),
.C(n_375),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_37),
.C(n_3),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_371),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_361),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_403),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_374),
.Y(n_399)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_410),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_405),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_383),
.C(n_382),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_394),
.C(n_393),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_395),
.B(n_373),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_384),
.A2(n_369),
.B(n_373),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_406),
.B(n_407),
.Y(n_411)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_361),
.B1(n_4),
.B2(n_5),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_408),
.A2(n_409),
.B1(n_13),
.B2(n_4),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_390),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_416),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_388),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_401),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_396),
.A2(n_386),
.B(n_387),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_418),
.B(n_422),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_37),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_421),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_37),
.C(n_0),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_5),
.C(n_6),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_400),
.B(n_4),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_423),
.B(n_430),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_398),
.B(n_408),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_425),
.A2(n_413),
.B(n_418),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_422),
.A2(n_398),
.B1(n_410),
.B2(n_409),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_429),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_5),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_412),
.B(n_6),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_431),
.B(n_9),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_435),
.B(n_436),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_12),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_420),
.B(n_415),
.Y(n_435)
);

OAI21x1_ASAP7_75t_SL g436 ( 
.A1(n_424),
.A2(n_9),
.B(n_11),
.Y(n_436)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_438),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_439),
.A2(n_433),
.B1(n_428),
.B2(n_423),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_440),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_430),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_444),
.A2(n_441),
.B(n_429),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_49),
.Y(n_446)
);


endmodule