module real_jpeg_30069_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_57;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_0),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_18),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_14),
.Y(n_13)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_2),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_4),
.A2(n_12),
.B1(n_16),
.B2(n_21),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_4),
.A2(n_46),
.B(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_46),
.Y(n_48)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_14),
.B1(n_17),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_34),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_29),
.B(n_33),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_24),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_11),
.B(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_36)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_14),
.B(n_27),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI32xp33_ASAP7_75t_L g52 ( 
.A1(n_17),
.A2(n_26),
.A3(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_28),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_25),
.B(n_50),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_56),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_52),
.B2(n_55),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);


endmodule