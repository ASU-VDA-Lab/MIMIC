module fake_jpeg_7002_n_263 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_25),
.B1(n_18),
.B2(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_61),
.B(n_65),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_59),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_74),
.B1(n_78),
.B2(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_29),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_67),
.Y(n_109)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_63),
.B(n_66),
.Y(n_104)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_27),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_26),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_34),
.A2(n_20),
.B1(n_14),
.B2(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_34),
.A2(n_20),
.B1(n_22),
.B2(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_1),
.Y(n_107)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_35),
.A2(n_17),
.B1(n_22),
.B2(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_34),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_31),
.B1(n_30),
.B2(n_4),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_49),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_115),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_12),
.B1(n_13),
.B2(n_68),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_31),
.B(n_30),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_110),
.B(n_117),
.C(n_12),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_2),
.B(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_2),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_9),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_7),
.B(n_9),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_53),
.B1(n_65),
.B2(n_61),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_134),
.B1(n_143),
.B2(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_48),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_135),
.B(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_144),
.B1(n_145),
.B2(n_149),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_92),
.A2(n_86),
.B(n_88),
.C(n_77),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_132),
.B(n_121),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_10),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_62),
.B1(n_48),
.B2(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_10),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_59),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_83),
.B1(n_77),
.B2(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_13),
.B1(n_102),
.B2(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_117),
.B1(n_114),
.B2(n_96),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_115),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_135),
.B(n_148),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_98),
.B(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_96),
.B1(n_94),
.B2(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_160),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_93),
.B1(n_121),
.B2(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_164),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_98),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_166),
.Y(n_190)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_127),
.B1(n_146),
.B2(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_174),
.B(n_176),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_143),
.B1(n_134),
.B2(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_150),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_129),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_180),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_125),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_138),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_164),
.C(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_197),
.Y(n_204)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_152),
.B1(n_156),
.B2(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_188),
.C(n_192),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_177),
.B(n_191),
.C(n_181),
.D(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_206),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_167),
.B(n_161),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_193),
.B(n_182),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_156),
.A3(n_157),
.B1(n_172),
.B2(n_152),
.C1(n_165),
.C2(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_221),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_199),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_225),
.B(n_198),
.Y(n_234)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_201),
.C(n_215),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_230),
.C(n_236),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_203),
.C(n_213),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_237),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_219),
.C(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_204),
.B1(n_205),
.B2(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_204),
.B1(n_200),
.B2(n_214),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_246),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_227),
.C(n_222),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_222),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_200),
.Y(n_255)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_207),
.C(n_214),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_239),
.B(n_185),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_255),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_247),
.B1(n_235),
.B2(n_252),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_155),
.C(n_250),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_240),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_259),
.C(n_253),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_250),
.Y(n_263)
);


endmodule