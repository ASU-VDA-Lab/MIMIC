module real_aes_7019_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g490 ( .A(n_1), .Y(n_490) );
INVx1_ASAP7_75t_L g269 ( .A(n_2), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_3), .A2(n_37), .B1(n_188), .B2(n_518), .Y(n_517) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_4), .A2(n_177), .B(n_178), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_5), .B(n_175), .Y(n_467) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_7), .A2(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_10), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g147 ( .A(n_11), .Y(n_147) );
INVx1_ASAP7_75t_L g486 ( .A(n_12), .Y(n_486) );
INVx1_ASAP7_75t_L g251 ( .A(n_13), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_14), .B(n_153), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_15), .B(n_143), .Y(n_495) );
AO32x2_ASAP7_75t_L g515 ( .A1(n_16), .A2(n_142), .A3(n_175), .B1(n_478), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_17), .B(n_188), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_18), .B(n_196), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_19), .B(n_143), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_20), .A2(n_50), .B1(n_188), .B2(n_518), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_21), .B(n_177), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_22), .A2(n_76), .B1(n_153), .B2(n_188), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_23), .B(n_188), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_24), .B(n_173), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_25), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_26), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_27), .B(n_190), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_28), .B(n_183), .Y(n_270) );
INVx1_ASAP7_75t_L g161 ( .A(n_29), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_30), .B(n_190), .Y(n_512) );
INVx2_ASAP7_75t_L g155 ( .A(n_31), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_32), .B(n_188), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_33), .B(n_190), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_34), .A2(n_104), .B1(n_115), .B2(n_751), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_35), .A2(n_42), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_35), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_36), .A2(n_150), .B(n_162), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g159 ( .A(n_39), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_40), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_41), .B(n_183), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_42), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_43), .B(n_188), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_44), .A2(n_87), .B1(n_213), .B2(n_518), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_45), .B(n_188), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_46), .B(n_188), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_47), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_48), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_49), .B(n_177), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_51), .A2(n_60), .B1(n_153), .B2(n_188), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_52), .A2(n_153), .B1(n_156), .B2(n_162), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_53), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_54), .B(n_188), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_55), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_56), .B(n_188), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_57), .A2(n_182), .B(n_184), .C(n_187), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_58), .Y(n_226) );
INVx1_ASAP7_75t_L g179 ( .A(n_59), .Y(n_179) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_62), .B(n_188), .Y(n_491) );
INVx1_ASAP7_75t_L g146 ( .A(n_63), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_65), .A2(n_175), .A3(n_231), .B1(n_478), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g475 ( .A(n_66), .Y(n_475) );
INVx1_ASAP7_75t_L g507 ( .A(n_67), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_68), .A2(n_745), .B1(n_746), .B2(n_749), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_68), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_SL g195 ( .A1(n_69), .A2(n_187), .B(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g198 ( .A(n_70), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_71), .B(n_153), .Y(n_508) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_73), .Y(n_170) );
INVx1_ASAP7_75t_L g219 ( .A(n_74), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_75), .A2(n_101), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_75), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_77), .A2(n_150), .B(n_162), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_78), .B(n_518), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_79), .B(n_153), .Y(n_511) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_80), .A2(n_126), .B1(n_127), .B2(n_133), .C1(n_734), .C2(n_737), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_81), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_83), .B(n_196), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_84), .B(n_153), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_85), .A2(n_150), .B(n_162), .C(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g110 ( .A(n_86), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g449 ( .A(n_86), .B(n_112), .Y(n_449) );
INVx2_ASAP7_75t_L g733 ( .A(n_86), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_88), .A2(n_102), .B1(n_153), .B2(n_154), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_89), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_90), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_91), .A2(n_150), .B(n_162), .C(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_92), .Y(n_241) );
INVx1_ASAP7_75t_L g194 ( .A(n_93), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_94), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_95), .B(n_209), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_96), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_96), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_97), .B(n_153), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_98), .B(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_99), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_100), .A2(n_177), .B(n_193), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_101), .Y(n_132) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g752 ( .A(n_105), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g123 ( .A(n_110), .Y(n_123) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_110), .Y(n_750) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_111), .B(n_733), .Y(n_739) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g732 ( .A(n_112), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_125), .B1(n_740), .B2(n_741), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g740 ( .A(n_119), .Y(n_740) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_122), .A2(n_742), .B(n_750), .Y(n_741) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_447), .B1(n_450), .B2(n_730), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_134), .A2(n_135), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_135), .A2(n_447), .B1(n_735), .B2(n_736), .Y(n_734) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_372), .C(n_421), .Y(n_135) );
NOR3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_279), .C(n_317), .Y(n_136) );
OAI222xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_200), .B1(n_254), .B2(n_260), .C1(n_274), .C2(n_277), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_139), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_139), .B(n_322), .Y(n_413) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g290 ( .A(n_140), .B(n_191), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_140), .B(n_172), .Y(n_298) );
AND2x2_ASAP7_75t_L g333 ( .A(n_140), .B(n_310), .Y(n_333) );
OR2x2_ASAP7_75t_L g357 ( .A(n_140), .B(n_172), .Y(n_357) );
OR2x2_ASAP7_75t_L g365 ( .A(n_140), .B(n_264), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_140), .B(n_191), .Y(n_368) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g262 ( .A(n_141), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_141), .B(n_191), .Y(n_276) );
AND2x2_ASAP7_75t_L g326 ( .A(n_141), .B(n_264), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_141), .B(n_172), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_141), .B(n_425), .Y(n_446) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_169), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_142), .A2(n_265), .B(n_272), .Y(n_264) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_144), .B(n_145), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B1(n_165), .B2(n_166), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_180), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_149), .A2(n_180), .B(n_247), .C(n_248), .Y(n_246) );
INVx4_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_150), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g177 ( .A(n_150), .B(n_167), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_150), .A2(n_459), .B(n_462), .Y(n_458) );
BUFx3_ASAP7_75t_L g478 ( .A(n_150), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_150), .A2(n_485), .B(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_150), .A2(n_506), .B(n_509), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_522), .B(n_526), .Y(n_521) );
INVx2_ASAP7_75t_L g271 ( .A(n_153), .Y(n_271) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx4_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
AND2x2_ASAP7_75t_L g167 ( .A(n_158), .B(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx3_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx1_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx5_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
AND2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
BUFx3_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
INVx1_ASAP7_75t_L g518 ( .A(n_163), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_166), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_166), .A2(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g465 ( .A(n_168), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_171), .A2(n_365), .B(n_366), .C(n_369), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_171), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_171), .B(n_309), .Y(n_431) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_191), .Y(n_171) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_172), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_172), .B(n_310), .Y(n_316) );
INVx1_ASAP7_75t_SL g324 ( .A(n_172), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_172), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g425 ( .A(n_172), .Y(n_425) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_189), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_174), .B(n_216), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_174), .B(n_478), .C(n_497), .Y(n_496) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_174), .A2(n_497), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_175), .A2(n_192), .B(n_199), .Y(n_191) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_175), .A2(n_458), .B(n_467), .Y(n_457) );
BUFx2_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_182), .A2(n_475), .B(n_476), .C(n_477), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_182), .A2(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx4_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_183), .A2(n_466), .B1(n_498), .B2(n_499), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_183), .A2(n_466), .B1(n_517), .B2(n_519), .Y(n_516) );
OAI22xp5_ASAP7_75t_SL g536 ( .A1(n_183), .A2(n_186), .B1(n_537), .B2(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_186), .B(n_198), .Y(n_197) );
INVx5_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_SL g506 ( .A1(n_187), .A2(n_209), .B(n_507), .C(n_508), .Y(n_506) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
INVx1_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_244), .B(n_253), .Y(n_243) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_190), .A2(n_505), .B(n_512), .Y(n_504) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_190), .A2(n_521), .B(n_529), .Y(n_520) );
BUFx2_ASAP7_75t_L g261 ( .A(n_191), .Y(n_261) );
INVx1_ASAP7_75t_L g323 ( .A(n_191), .Y(n_323) );
INVx3_ASAP7_75t_L g348 ( .A(n_191), .Y(n_348) );
INVx1_ASAP7_75t_L g525 ( .A(n_196), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_200), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_228), .Y(n_200) );
INVx1_ASAP7_75t_L g344 ( .A(n_201), .Y(n_344) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_201), .A2(n_289), .A3(n_351), .B1(n_352), .B2(n_353), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_201), .A2(n_355), .B1(n_358), .B2(n_363), .Y(n_354) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g292 ( .A(n_202), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g370 ( .A(n_202), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g440 ( .A(n_202), .B(n_386), .Y(n_440) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g255 ( .A(n_203), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
INVx1_ASAP7_75t_L g304 ( .A(n_203), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_203), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_203), .B(n_293), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_203), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_203), .B(n_258), .Y(n_340) );
INVx3_ASAP7_75t_L g362 ( .A(n_203), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_203), .B(n_259), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_203), .B(n_352), .Y(n_435) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_214), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_211), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_209), .A2(n_269), .B(n_270), .C(n_271), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_209), .A2(n_460), .B(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g466 ( .A(n_209), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_209), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g252 ( .A(n_213), .Y(n_252) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_214), .A2(n_470), .B(n_479), .Y(n_469) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_214), .A2(n_484), .B(n_492), .Y(n_483) );
INVx2_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
AND2x2_ASAP7_75t_L g391 ( .A(n_217), .B(n_229), .Y(n_391) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_227), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_227), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g433 ( .A(n_228), .Y(n_433) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_229), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_229), .B(n_259), .Y(n_313) );
AND2x2_ASAP7_75t_L g371 ( .A(n_229), .B(n_294), .Y(n_371) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g257 ( .A(n_230), .Y(n_257) );
AND2x2_ASAP7_75t_L g284 ( .A(n_230), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_230), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_230), .B(n_259), .Y(n_359) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_240), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_242), .B(n_259), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_242), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g386 ( .A(n_242), .Y(n_386) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_243), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_249), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g488 ( .A(n_249), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_249), .A2(n_510), .B(n_511), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_264), .B1(n_423), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_256), .A2(n_367), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_257), .B(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g404 ( .A(n_257), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_258), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g331 ( .A(n_258), .B(n_284), .Y(n_331) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_412), .B1(n_429), .B2(n_432), .C(n_434), .Y(n_428) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_261), .B(n_310), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_262), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g353 ( .A(n_262), .B(n_299), .Y(n_353) );
INVx3_ASAP7_75t_SL g394 ( .A(n_262), .Y(n_394) );
AND2x2_ASAP7_75t_L g338 ( .A(n_263), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_263), .B(n_276), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_263), .B(n_322), .Y(n_408) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
OAI322xp33_ASAP7_75t_L g405 ( .A1(n_264), .A2(n_336), .A3(n_358), .B1(n_406), .B2(n_408), .C1(n_409), .C2(n_410), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_271), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_275), .A2(n_278), .B(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_276), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g377 ( .A(n_276), .B(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_276), .B(n_316), .Y(n_392) );
INVxp67_ASAP7_75t_L g343 ( .A(n_278), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_278), .A2(n_350), .B(n_354), .C(n_364), .Y(n_349) );
OAI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_288), .B1(n_291), .B2(n_295), .C(n_300), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g303 ( .A(n_287), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_288), .A2(n_437), .B1(n_442), .B2(n_443), .C(n_445), .Y(n_436) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_289), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g336 ( .A(n_289), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_289), .B(n_367), .Y(n_374) );
AND2x2_ASAP7_75t_L g416 ( .A(n_289), .B(n_394), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_290), .B(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_290), .A2(n_302), .B1(n_412), .B2(n_413), .Y(n_411) );
OR2x2_ASAP7_75t_L g442 ( .A(n_290), .B(n_310), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g419 ( .A(n_293), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_293), .B(n_387), .Y(n_444) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_298), .B(n_309), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B1(n_311), .B2(n_314), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g375 ( .A(n_303), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_303), .B(n_343), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g334 ( .A1(n_305), .A2(n_335), .A3(n_337), .B1(n_338), .B2(n_340), .C1(n_341), .C2(n_345), .Y(n_334) );
INVxp67_ASAP7_75t_L g328 ( .A(n_306), .Y(n_328) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_308), .A2(n_313), .B1(n_330), .B2(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_309), .B(n_322), .Y(n_409) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_310), .B(n_348), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_334), .C(n_349), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_325), .B2(n_327), .C(n_329), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_321), .B(n_326), .Y(n_325) );
INVx3_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_328), .Y(n_407) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_333), .B(n_347), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_336), .B(n_394), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_337), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g412 ( .A(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g427 ( .A(n_340), .B(n_404), .Y(n_427) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_351), .A2(n_422), .B(n_428), .C(n_436), .Y(n_421) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_391), .Y(n_390) );
NAND2x1_ASAP7_75t_SL g432 ( .A(n_362), .B(n_433), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_387), .Y(n_401) );
NOR5xp2_ASAP7_75t_L g372 ( .A(n_373), .B(n_388), .C(n_405), .D(n_411), .E(n_414), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_378), .C(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_377), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_387), .B(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_392), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AOI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_417), .B(n_419), .C(n_420), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g735 ( .A(n_450), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_451), .B(n_654), .Y(n_450) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_612), .Y(n_451) );
NOR4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_552), .C(n_588), .D(n_602), .Y(n_452) );
OAI221xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_500), .B1(n_530), .B2(n_539), .C(n_543), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_454), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_480), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
AND2x2_ASAP7_75t_L g549 ( .A(n_457), .B(n_469), .Y(n_549) );
INVx3_ASAP7_75t_L g557 ( .A(n_457), .Y(n_557) );
AND2x2_ASAP7_75t_L g611 ( .A(n_457), .B(n_483), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_457), .B(n_482), .Y(n_647) );
AND2x2_ASAP7_75t_L g705 ( .A(n_457), .B(n_567), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_466), .Y(n_462) );
INVx2_ASAP7_75t_L g476 ( .A(n_465), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_466), .A2(n_476), .B(n_490), .C(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g540 ( .A(n_468), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g554 ( .A(n_468), .B(n_483), .Y(n_554) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_469), .B(n_483), .Y(n_569) );
AND2x2_ASAP7_75t_L g581 ( .A(n_469), .B(n_557), .Y(n_581) );
OR2x2_ASAP7_75t_L g583 ( .A(n_469), .B(n_541), .Y(n_583) );
AND2x2_ASAP7_75t_L g618 ( .A(n_469), .B(n_541), .Y(n_618) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_469), .Y(n_663) );
INVx1_ASAP7_75t_L g671 ( .A(n_469), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B(n_478), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_480), .A2(n_589), .B1(n_593), .B2(n_597), .C(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g548 ( .A(n_481), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
INVx2_ASAP7_75t_L g547 ( .A(n_482), .Y(n_547) );
AND2x2_ASAP7_75t_L g600 ( .A(n_482), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g619 ( .A(n_482), .B(n_557), .Y(n_619) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g682 ( .A(n_483), .B(n_557), .Y(n_682) );
AND2x2_ASAP7_75t_L g604 ( .A(n_493), .B(n_549), .Y(n_604) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_493), .A2(n_628), .A3(n_673), .B1(n_675), .B2(n_678), .C1(n_680), .C2(n_684), .Y(n_672) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_494), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g568 ( .A(n_494), .Y(n_568) );
AND2x2_ASAP7_75t_L g677 ( .A(n_494), .B(n_557), .Y(n_677) );
AND2x2_ASAP7_75t_L g709 ( .A(n_494), .B(n_581), .Y(n_709) );
OR2x2_ASAP7_75t_L g712 ( .A(n_494), .B(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g542 ( .A(n_495), .Y(n_542) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
INVx1_ASAP7_75t_L g725 ( .A(n_502), .Y(n_725) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g532 ( .A(n_503), .B(n_520), .Y(n_532) );
INVx2_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_504), .Y(n_595) );
OR2x2_ASAP7_75t_L g719 ( .A(n_504), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g544 ( .A(n_513), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g584 ( .A(n_513), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g636 ( .A(n_513), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
AND2x2_ASAP7_75t_L g533 ( .A(n_514), .B(n_534), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g591 ( .A(n_514), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g645 ( .A(n_514), .B(n_535), .Y(n_645) );
OR2x2_ASAP7_75t_L g653 ( .A(n_514), .B(n_587), .Y(n_653) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_515), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g596 ( .A(n_515), .B(n_520), .Y(n_596) );
AND2x2_ASAP7_75t_L g660 ( .A(n_515), .B(n_535), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_520), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_520), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
INVx1_ASAP7_75t_L g578 ( .A(n_520), .Y(n_578) );
AND2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_591), .Y(n_590) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_520), .Y(n_668) );
INVx1_ASAP7_75t_L g720 ( .A(n_520), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g697 ( .A(n_531), .B(n_606), .Y(n_697) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g624 ( .A(n_533), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g723 ( .A(n_533), .B(n_658), .Y(n_723) );
INVx1_ASAP7_75t_L g545 ( .A(n_534), .Y(n_545) );
AND2x2_ASAP7_75t_L g571 ( .A(n_534), .B(n_565), .Y(n_571) );
BUFx2_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
INVx1_ASAP7_75t_L g561 ( .A(n_535), .Y(n_561) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_539), .B(n_546), .Y(n_699) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI32xp33_ASAP7_75t_L g543 ( .A1(n_540), .A2(n_544), .A3(n_546), .B1(n_548), .B2(n_550), .Y(n_543) );
AND2x2_ASAP7_75t_L g683 ( .A(n_540), .B(n_556), .Y(n_683) );
AND2x2_ASAP7_75t_L g721 ( .A(n_540), .B(n_619), .Y(n_721) );
INVx1_ASAP7_75t_L g601 ( .A(n_541), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_545), .B(n_607), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_546), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_546), .B(n_549), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_546), .B(n_618), .Y(n_700) );
OR2x2_ASAP7_75t_L g714 ( .A(n_546), .B(n_583), .Y(n_714) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g641 ( .A(n_547), .B(n_549), .Y(n_641) );
OR2x2_ASAP7_75t_L g650 ( .A(n_547), .B(n_637), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_549), .B(n_600), .Y(n_622) );
INVx2_ASAP7_75t_L g637 ( .A(n_551), .Y(n_637) );
OR2x2_ASAP7_75t_L g652 ( .A(n_551), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g667 ( .A(n_551), .B(n_668), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_551), .A2(n_644), .B(n_725), .C(n_726), .Y(n_724) );
OAI321xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_558), .A3(n_563), .B1(n_566), .B2(n_570), .C(n_574), .Y(n_552) );
INVx1_ASAP7_75t_L g665 ( .A(n_553), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g676 ( .A(n_554), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g628 ( .A(n_556), .Y(n_628) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_557), .B(n_671), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_558), .A2(n_696), .B1(n_698), .B2(n_700), .C(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x2_ASAP7_75t_L g633 ( .A(n_560), .B(n_607), .Y(n_633) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_561), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g606 ( .A(n_562), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_563), .A2(n_604), .B(n_649), .C(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g615 ( .A(n_565), .B(n_572), .Y(n_615) );
BUFx2_ASAP7_75t_L g625 ( .A(n_565), .Y(n_625) );
INVx1_ASAP7_75t_L g640 ( .A(n_565), .Y(n_640) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g646 ( .A(n_568), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g729 ( .A(n_568), .Y(n_729) );
INVx1_ASAP7_75t_L g722 ( .A(n_569), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g575 ( .A(n_571), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g679 ( .A(n_571), .B(n_596), .Y(n_679) );
INVx1_ASAP7_75t_L g608 ( .A(n_572), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B1(n_582), .B2(n_584), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_576), .B(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g644 ( .A(n_577), .B(n_645), .Y(n_644) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_578), .B(n_587), .Y(n_607) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g599 ( .A(n_581), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g609 ( .A(n_583), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_586), .A2(n_704), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_703) );
INVx1_ASAP7_75t_L g592 ( .A(n_587), .Y(n_592) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_590), .B(n_709), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_591), .A2(n_596), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_594), .B(n_604), .Y(n_701) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g670 ( .A(n_595), .Y(n_670) );
AND2x2_ASAP7_75t_L g629 ( .A(n_596), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g718 ( .A(n_596), .Y(n_718) );
INVx1_ASAP7_75t_L g634 ( .A(n_599), .Y(n_634) );
INVx1_ASAP7_75t_L g689 ( .A(n_600), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_606), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g674 ( .A(n_607), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_607), .B(n_645), .Y(n_711) );
OR2x2_ASAP7_75t_L g684 ( .A(n_608), .B(n_637), .Y(n_684) );
INVx1_ASAP7_75t_L g623 ( .A(n_609), .Y(n_623) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_611), .B(n_662), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_631), .C(n_642), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_620), .C(n_626), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_615), .A2(n_686), .B1(n_690), .B2(n_693), .C(n_695), .Y(n_685) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g627 ( .A(n_618), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g681 ( .A(n_618), .B(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_619), .A2(n_667), .B(n_669), .C(n_671), .Y(n_666) );
INVx2_ASAP7_75t_L g713 ( .A(n_619), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_623), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g692 ( .A(n_625), .B(n_645), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_634), .B(n_635), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_638), .B(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_636), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_641), .B(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B(n_648), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g669 ( .A(n_645), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND4x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_685), .C(n_702), .D(n_724), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_672), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_661), .B(n_664), .C(n_666), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_660), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_671), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g706 ( .A(n_681), .Y(n_706) );
INVx2_ASAP7_75t_SL g694 ( .A(n_682), .Y(n_694) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g707 ( .A(n_692), .Y(n_707) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_SL g702 ( .A(n_703), .B(n_710), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_712), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g736 ( .A(n_731), .Y(n_736) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
endmodule