module fake_jpeg_8913_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_14),
.B1(n_15),
.B2(n_10),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_33),
.B1(n_13),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_14),
.B1(n_10),
.B2(n_15),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_35),
.B1(n_39),
.B2(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_18),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_49),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_12),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_35),
.B1(n_41),
.B2(n_29),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_40),
.C(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_2),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_51),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_51),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_59),
.C(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_77),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_65),
.B(n_57),
.C(n_66),
.D(n_67),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_57),
.B(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_77),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_59),
.C(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_79),
.B1(n_70),
.B2(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_73),
.C(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_56),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_86),
.B1(n_87),
.B2(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_69),
.B(n_57),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_17),
.B(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_25),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_103),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_98),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B(n_3),
.C(n_25),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_3),
.Y(n_108)
);


endmodule