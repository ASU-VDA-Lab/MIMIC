module fake_jpeg_613_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_20),
.B1(n_22),
.B2(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_19),
.B1(n_18),
.B2(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_34),
.B1(n_29),
.B2(n_23),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_19),
.B1(n_13),
.B2(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_33),
.B1(n_30),
.B2(n_14),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_26),
.C(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.C(n_17),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_29),
.C(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_39),
.B1(n_30),
.B2(n_42),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.C(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_43),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_31),
.B(n_14),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_14),
.B(n_2),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_14),
.Y(n_54)
);


endmodule