module fake_jpeg_29345_n_119 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_38),
.B(n_5),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_2),
.C(n_4),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_5),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_5),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_49),
.B(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_26),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_28),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_23),
.B1(n_20),
.B2(n_11),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_27),
.A2(n_20),
.B1(n_11),
.B2(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_11),
.B1(n_17),
.B2(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_29),
.A2(n_17),
.B1(n_7),
.B2(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_7),
.B1(n_17),
.B2(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_59),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_57),
.A3(n_60),
.B1(n_47),
.B2(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_60),
.B1(n_45),
.B2(n_47),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_74),
.B1(n_73),
.B2(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_69),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_68),
.B(n_75),
.Y(n_99)
);

AOI21x1_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_81),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_102),
.B(n_100),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_95),
.C(n_80),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_109),
.B(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_97),
.B1(n_94),
.B2(n_92),
.Y(n_108)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_106),
.A3(n_102),
.B1(n_105),
.B2(n_84),
.C(n_76),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.C(n_65),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_87),
.C(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_78),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.C(n_85),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_115),
.B(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_78),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_52),
.Y(n_119)
);


endmodule