module real_jpeg_6938_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_1),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_2),
.B(n_60),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_2),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_2),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_2),
.B(n_429),
.Y(n_428)
);

NAND2x1_ASAP7_75t_SL g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_3),
.B(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_4),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_4),
.Y(n_408)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_7),
.Y(n_134)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_7),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_10),
.B(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_10),
.B(n_114),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_10),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_10),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_10),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_10),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_10),
.B(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_42),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_12),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_12),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_12),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_13),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_13),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_13),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_13),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_13),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_13),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_13),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_14),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_14),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_14),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_14),
.B(n_419),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_162),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_161),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_96),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_20),
.B(n_96),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_20),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_43),
.CI(n_80),
.CON(n_20),
.SN(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.C(n_38),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_22),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.C(n_31),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_47),
.C(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_23),
.A2(n_47),
.B1(n_48),
.B2(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_23),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_23),
.A2(n_95),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_23),
.A2(n_95),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_23),
.B(n_172),
.C(n_177),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_33),
.Y(n_32)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_26),
.Y(n_387)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_27),
.Y(n_289)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_27),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_28),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_31),
.A2(n_32),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_31),
.A2(n_32),
.B1(n_183),
.B2(n_300),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_32),
.B(n_103),
.C(n_108),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_32),
.B(n_182),
.C(n_183),
.Y(n_181)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_37),
.B(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_42),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_43)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_59),
.B2(n_63),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_58),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_47),
.A2(n_48),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_48),
.B(n_201),
.C(n_206),
.Y(n_290)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_50),
.Y(n_312)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_51),
.Y(n_228)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_51),
.Y(n_345)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_51),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_52),
.B(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_56),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_56),
.Y(n_255)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_58),
.B(n_265),
.C(n_270),
.Y(n_326)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_63),
.B1(n_118),
.B2(n_126),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_59),
.B(n_119),
.C(n_125),
.Y(n_157)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_69),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_103),
.C(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_68),
.A2(n_69),
.B1(n_112),
.B2(n_113),
.Y(n_329)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_73),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_92),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_81),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_92),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.C(n_91),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_88),
.A2(n_89),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_89),
.B(n_133),
.C(n_188),
.Y(n_346)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_151),
.C(n_159),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_97),
.B(n_151),
.CI(n_159),
.CON(n_487),
.SN(n_487)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_127),
.C(n_130),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_98),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.C(n_117),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_99),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_108),
.B2(n_110),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_102),
.A2(n_103),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_103),
.B(n_202),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_103),
.B(n_202),
.Y(n_381)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_111),
.B(n_117),
.Y(n_354)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_116),
.Y(n_307)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_122),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_122),
.B(n_249),
.C(n_254),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_127),
.B(n_130),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_142),
.C(n_146),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g361 ( 
.A1(n_131),
.A2(n_132),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_133),
.A2(n_188),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_133),
.A2(n_141),
.B1(n_277),
.B2(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_133),
.B(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_133),
.A2(n_277),
.B1(n_372),
.B2(n_373),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_135),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_223),
.C(n_226),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_135),
.A2(n_229),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_139),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_140),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_141),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_146),
.A2(n_147),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_147),
.B(n_342),
.C(n_346),
.Y(n_360)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_158),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_152),
.A2(n_153),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_157),
.B(n_158),
.Y(n_485)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_478),
.B(n_492),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_349),
.B(n_364),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_320),
.B(n_348),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_291),
.B(n_319),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_166),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_257),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_167),
.B(n_257),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_221),
.C(n_245),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_168),
.B(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_197),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_198),
.C(n_208),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_181),
.C(n_186),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_170),
.B(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_181),
.A2(n_186),
.B1(n_187),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_181),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_182),
.B(n_299),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_183),
.Y(n_300)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_188),
.A2(n_193),
.B1(n_194),
.B2(n_278),
.Y(n_313)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_191),
.Y(n_431)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g375 ( 
.A(n_192),
.Y(n_375)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_204),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_208),
.Y(n_498)
);

FAx1_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.CI(n_218),
.CON(n_208),
.SN(n_208)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_210),
.B(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_213),
.C(n_218),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_219),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_221),
.B(n_245),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.C(n_233),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_222),
.A2(n_231),
.B1(n_232),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_224),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_224),
.B(n_424),
.Y(n_444)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_233),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_241),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_234),
.A2(n_235),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_236),
.A2(n_237),
.B1(n_241),
.B2(n_242),
.Y(n_466)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_239),
.Y(n_411)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_256),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_248),
.C(n_256),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_260),
.C(n_279),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_279),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_274),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_263),
.C(n_274),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_287),
.C(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_317),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_292),
.B(n_317),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.C(n_314),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_293),
.A2(n_294),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_297),
.B(n_314),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.C(n_313),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_298),
.B(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_301),
.B(n_313),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.C(n_308),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_302),
.A2(n_303),
.B1(n_308),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_305),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_309),
.B(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_321),
.B(n_349),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_323),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_350),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_323),
.B(n_350),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_334),
.CI(n_347),
.CON(n_323),
.SN(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_327),
.C(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_337),
.C(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_351),
.B(n_353),
.C(n_355),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_356),
.B(n_360),
.C(n_361),
.Y(n_486)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OAI31xp33_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_474),
.A3(n_475),
.B(n_477),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_468),
.B(n_473),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_455),
.B(n_467),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_413),
.B(n_454),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_399),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_369),
.B(n_399),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_382),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_370),
.B(n_383),
.C(n_396),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_371),
.B(n_377),
.C(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_396),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.C(n_393),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_384),
.B(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_388),
.A2(n_389),
.B1(n_393),
.B2(n_394),
.Y(n_401)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.C(n_412),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_451),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_403),
.B1(n_412),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_405),
.B1(n_409),
.B2(n_410),
.Y(n_425)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_448),
.B(n_453),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_435),
.B(n_447),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_426),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_426),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_425),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_422),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_422),
.C(n_425),
.Y(n_449)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_428),
.B1(n_432),
.B2(n_433),
.Y(n_445)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_443),
.B(n_446),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_444),
.B(n_445),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_450),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_457),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_462),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_463),
.C(n_464),
.Y(n_472)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_472),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_472),
.Y(n_473)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_488),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_479),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_487),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_487),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.C(n_486),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_483),
.Y(n_491)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_491),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_487),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_490),
.Y(n_493)
);


endmodule