module fake_jpeg_911_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_24),
.B1(n_13),
.B2(n_14),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_17),
.B1(n_14),
.B2(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_27),
.B1(n_22),
.B2(n_13),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_50),
.B1(n_20),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_53),
.B1(n_28),
.B2(n_39),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_17),
.B1(n_40),
.B2(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_16),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_26),
.B1(n_20),
.B2(n_28),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_73),
.B(n_46),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_44),
.B(n_43),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_43),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_9),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_36),
.C(n_20),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_57),
.B1(n_46),
.B2(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_80),
.B1(n_88),
.B2(n_67),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_84),
.C(n_86),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_43),
.B1(n_54),
.B2(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_72),
.C(n_71),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_98),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_60),
.C(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_101),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_77),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_61),
.C(n_64),
.Y(n_100)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_87),
.A3(n_78),
.B1(n_84),
.B2(n_88),
.C(n_76),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_66),
.B1(n_70),
.B2(n_67),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_70),
.B1(n_89),
.B2(n_101),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_97),
.C(n_100),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_91),
.C(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_65),
.B(n_75),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_106),
.B(n_58),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_111),
.C(n_108),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_110),
.B(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_115),
.B(n_114),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.C(n_58),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_120),
.B1(n_119),
.B2(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_89),
.B1(n_65),
.B2(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_3),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_129),
.B(n_131),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_3),
.Y(n_134)
);


endmodule