module fake_netlist_6_2700_n_1217 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1217);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1217;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_1212;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_1209;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1099;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_1120;
wire n_369;
wire n_894;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1216;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_953;
wire n_1094;
wire n_1004;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_1213;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_1211;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_172;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_1215;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_1152;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1041;
wire n_279;
wire n_686;
wire n_796;
wire n_1000;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_1090;
wire n_395;
wire n_813;
wire n_592;
wire n_912;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1207;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_121),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_77),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_8),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_62),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_74),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_119),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_113),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_149),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_107),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_70),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_82),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_22),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_108),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_8),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_31),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_26),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_63),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_110),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_157),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_26),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_20),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_111),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_76),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_52),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_128),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_47),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_20),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_4),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_167),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_130),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_122),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_109),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_90),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_80),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_116),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_45),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_155),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_129),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_12),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_106),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_127),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_150),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_100),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_17),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_81),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_112),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_97),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_43),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_44),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_131),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_42),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_145),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_40),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_168),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_40),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_0),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_0),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_160),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_171),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_173),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_171),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_179),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_180),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_173),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_171),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_171),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_191),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_210),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_191),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_219),
.B(n_2),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_217),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_217),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_206),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_213),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_228),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_2),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_237),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_180),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_249),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_218),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_218),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_238),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_182),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_182),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_257),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_238),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_284),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_278),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_243),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_212),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_286),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_212),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_190),
.B(n_214),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_174),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_190),
.B(n_3),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_288),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_262),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_243),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_186),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_196),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_208),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_214),
.B(n_3),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_263),
.B(n_4),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_252),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_255),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_263),
.B(n_5),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_255),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_209),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_221),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_223),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_229),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_247),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_188),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_267),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_178),
.B(n_5),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_177),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_248),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_267),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_178),
.B(n_9),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_254),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_261),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_188),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_172),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_279),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_252),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_279),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_200),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_265),
.Y(n_382)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_266),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_274),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_290),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_282),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_297),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_285),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_175),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_302),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_216),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_176),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_216),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_303),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_294),
.B(n_289),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

NAND2x1_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_177),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_315),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_242),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_294),
.B(n_289),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_353),
.B(n_177),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_375),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_330),
.B(n_289),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_183),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_319),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_347),
.B(n_184),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_185),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_348),
.B(n_192),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_355),
.B(n_193),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_319),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_355),
.B(n_195),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_312),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_327),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_374),
.B(n_287),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_359),
.B(n_197),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_291),
.B(n_296),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_293),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_304),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_354),
.B1(n_308),
.B2(n_177),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_369),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_405),
.B(n_366),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_L g455 ( 
.A1(n_448),
.A2(n_181),
.B1(n_227),
.B2(n_225),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_366),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_381),
.B(n_376),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_398),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_449),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_429),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_418),
.B(n_376),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_301),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_449),
.B(n_330),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

CKINVDCx12_ASAP7_75t_R g469 ( 
.A(n_409),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_293),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_295),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_251),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_427),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_429),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_449),
.B(n_295),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_436),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_442),
.A2(n_251),
.B1(n_275),
.B2(n_227),
.Y(n_485)
);

AO21x2_ASAP7_75t_L g486 ( 
.A1(n_389),
.A2(n_281),
.B(n_277),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_444),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_300),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_444),
.A2(n_251),
.B1(n_275),
.B2(n_181),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_436),
.B(n_251),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_275),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_382),
.B(n_385),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_449),
.A2(n_275),
.B1(n_225),
.B2(n_281),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_384),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_430),
.B(n_300),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_446),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_383),
.A2(n_385),
.B1(n_382),
.B2(n_421),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_384),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_437),
.B(n_313),
.Y(n_509)
);

NOR3xp33_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_447),
.C(n_441),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_395),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_440),
.A2(n_344),
.B1(n_321),
.B2(n_334),
.Y(n_515)
);

BUFx8_ASAP7_75t_SL g516 ( 
.A(n_431),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_403),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_434),
.B(n_313),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_451),
.B(n_460),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_454),
.A2(n_382),
.B1(n_385),
.B2(n_439),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_491),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_454),
.B(n_435),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_472),
.B(n_378),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_491),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_451),
.B(n_382),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_485),
.A2(n_383),
.B1(n_385),
.B2(n_421),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_497),
.B(n_409),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_445),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_485),
.A2(n_397),
.B1(n_412),
.B2(n_400),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_489),
.B(n_419),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_419),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

AND2x6_ASAP7_75t_SL g539 ( 
.A(n_474),
.B(n_440),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_515),
.B(n_317),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_474),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_403),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_403),
.Y(n_543)
);

AOI221xp5_ASAP7_75t_L g544 ( 
.A1(n_455),
.A2(n_378),
.B1(n_344),
.B2(n_339),
.C(n_317),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_404),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_492),
.A2(n_404),
.B1(n_407),
.B2(n_406),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_492),
.A2(n_407),
.B1(n_406),
.B2(n_413),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_509),
.B(n_403),
.Y(n_549)
);

NAND3xp33_ASAP7_75t_L g550 ( 
.A(n_499),
.B(n_321),
.C(n_320),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_320),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_406),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_474),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_451),
.B(n_406),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_455),
.B(n_299),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_451),
.B(n_406),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_490),
.A2(n_336),
.B1(n_339),
.B2(n_323),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_461),
.A2(n_415),
.B(n_401),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_451),
.B(n_413),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_452),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_459),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_505),
.A2(n_337),
.B1(n_305),
.B2(n_307),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_472),
.A2(n_326),
.B1(n_356),
.B2(n_358),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_481),
.B(n_413),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_460),
.B(n_323),
.Y(n_568)
);

BUFx6f_ASAP7_75t_SL g569 ( 
.A(n_501),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_460),
.B(n_372),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_460),
.B(n_198),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_465),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_490),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

NOR2x1p5_ASAP7_75t_L g577 ( 
.A(n_472),
.B(n_441),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_437),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_499),
.A2(n_415),
.B1(n_401),
.B2(n_417),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_476),
.A2(n_415),
.B1(n_417),
.B2(n_420),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_477),
.B(n_437),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_490),
.B(n_324),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_477),
.B(n_437),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_487),
.B(n_199),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

INVx8_ASAP7_75t_L g589 ( 
.A(n_479),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_487),
.B(n_201),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_452),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_483),
.B(n_417),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_484),
.A2(n_325),
.B1(n_332),
.B2(n_346),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_484),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_452),
.B(n_487),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_458),
.B(n_402),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_463),
.B(n_482),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_487),
.B(n_202),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_470),
.B(n_420),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_464),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_470),
.B(n_423),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_450),
.B(n_433),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_470),
.B(n_204),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_456),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_450),
.B(n_433),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_464),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_470),
.B(n_423),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_525),
.A2(n_510),
.B(n_467),
.C(n_520),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_521),
.A2(n_496),
.B(n_494),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_532),
.B(n_496),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_592),
.A2(n_504),
.B(n_510),
.C(n_486),
.Y(n_614)
);

A2O1A1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_522),
.A2(n_495),
.B(n_475),
.C(n_512),
.Y(n_615)
);

OA22x2_ASAP7_75t_L g616 ( 
.A1(n_541),
.A2(n_553),
.B1(n_575),
.B2(n_561),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_531),
.B(n_496),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_531),
.B(n_486),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_SL g619 ( 
.A1(n_528),
.A2(n_543),
.B(n_542),
.C(n_549),
.Y(n_619)
);

BUFx12f_ASAP7_75t_L g620 ( 
.A(n_539),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_528),
.A2(n_495),
.B(n_475),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_524),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_534),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_561),
.B(n_486),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_547),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_535),
.B(n_511),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_598),
.A2(n_608),
.B1(n_604),
.B2(n_545),
.Y(n_628)
);

NOR2x1_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_511),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_402),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_599),
.A2(n_545),
.B1(n_596),
.B2(n_537),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_588),
.A2(n_552),
.B(n_554),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_604),
.B(n_512),
.Y(n_634)
);

AO21x1_ASAP7_75t_L g635 ( 
.A1(n_572),
.A2(n_591),
.B(n_585),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_538),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_556),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_588),
.A2(n_517),
.B(n_500),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

CKINVDCx10_ASAP7_75t_R g641 ( 
.A(n_589),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_523),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_588),
.A2(n_517),
.B(n_500),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_608),
.B(n_519),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_588),
.A2(n_517),
.B(n_500),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_546),
.B(n_367),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_577),
.B(n_380),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_554),
.A2(n_517),
.B(n_514),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_530),
.B(n_519),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_557),
.A2(n_517),
.B(n_514),
.Y(n_650)
);

CKINVDCx10_ASAP7_75t_R g651 ( 
.A(n_589),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_533),
.B(n_513),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_583),
.B(n_432),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_548),
.B(n_513),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_567),
.B(n_513),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_567),
.B(n_518),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_597),
.B(n_514),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_529),
.B(n_516),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_518),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_557),
.A2(n_514),
.B(n_506),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_560),
.A2(n_514),
.B(n_506),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_560),
.A2(n_514),
.B(n_506),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_550),
.B(n_555),
.Y(n_663)
);

BUFx4f_ASAP7_75t_SL g664 ( 
.A(n_571),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_503),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_568),
.A2(n_518),
.B(n_410),
.C(n_428),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_558),
.B(n_469),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_574),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_544),
.B(n_410),
.C(n_408),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_595),
.B(n_471),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_593),
.A2(n_478),
.B(n_480),
.C(n_488),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_L g673 ( 
.A1(n_579),
.A2(n_411),
.B(n_408),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_582),
.B(n_471),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_527),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_607),
.B(n_471),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_569),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

NAND2x1_ASAP7_75t_L g680 ( 
.A(n_586),
.B(n_502),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_562),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_540),
.A2(n_508),
.B(n_416),
.C(n_411),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_562),
.B(n_502),
.Y(n_683)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_559),
.A2(n_488),
.B(n_480),
.C(n_478),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_573),
.B(n_462),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_551),
.A2(n_432),
.B1(n_438),
.B2(n_433),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_601),
.A2(n_498),
.B(n_473),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_603),
.A2(n_498),
.B(n_473),
.Y(n_688)
);

O2A1O1Ixp5_ASAP7_75t_L g689 ( 
.A1(n_581),
.A2(n_480),
.B(n_473),
.C(n_462),
.Y(n_689)
);

O2A1O1Ixp5_ASAP7_75t_L g690 ( 
.A1(n_584),
.A2(n_576),
.B(n_610),
.C(n_605),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_576),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_594),
.B(n_414),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_586),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_569),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_590),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_580),
.B(n_462),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_566),
.A2(n_498),
.B(n_423),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_578),
.A2(n_422),
.B(n_428),
.C(n_426),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_571),
.B(n_414),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_605),
.A2(n_498),
.B(n_422),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_590),
.B(n_395),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_565),
.B(n_569),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_624),
.Y(n_703)
);

BUFx2_ASAP7_75t_SL g704 ( 
.A(n_636),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_613),
.B(n_585),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_617),
.A2(n_600),
.B(n_591),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_611),
.A2(n_600),
.B(n_526),
.C(n_416),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_646),
.B(n_602),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_631),
.B(n_606),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_628),
.A2(n_606),
.B1(n_602),
.B2(n_609),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_628),
.B(n_387),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_649),
.A2(n_609),
.B1(n_564),
.B2(n_260),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_633),
.A2(n_619),
.B(n_612),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_618),
.A2(n_256),
.B1(n_207),
.B2(n_211),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_663),
.A2(n_424),
.B1(n_426),
.B2(n_438),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_SL g719 ( 
.A(n_702),
.B(n_253),
.C(n_215),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_653),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_625),
.B(n_387),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_630),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_625),
.B(n_390),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_699),
.B(n_390),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_630),
.B(n_589),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_678),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_635),
.B(n_220),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_637),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_663),
.B(n_589),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_638),
.B(n_498),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_621),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_692),
.B(n_424),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_614),
.A2(n_699),
.B(n_673),
.C(n_669),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_664),
.B(n_222),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_638),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_642),
.B(n_230),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_642),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_616),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_668),
.B(n_396),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_640),
.B(n_391),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_668),
.A2(n_259),
.B1(n_232),
.B2(n_280),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_666),
.A2(n_394),
.B(n_234),
.C(n_235),
.Y(n_744)
);

BUFx8_ASAP7_75t_SL g745 ( 
.A(n_620),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_664),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_678),
.B(n_498),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_629),
.B(n_634),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_644),
.A2(n_271),
.B1(n_270),
.B2(n_269),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_623),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_652),
.A2(n_264),
.B(n_246),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_694),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_694),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_632),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_627),
.B(n_245),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_622),
.A2(n_241),
.B(n_231),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_SL g758 ( 
.A(n_702),
.B(n_9),
.C(n_10),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_654),
.A2(n_657),
.B1(n_696),
.B2(n_615),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_670),
.B(n_10),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_670),
.B(n_11),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_679),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_691),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_677),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_SL g765 ( 
.A1(n_667),
.A2(n_69),
.B(n_164),
.C(n_163),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_682),
.B(n_48),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_SL g767 ( 
.A(n_658),
.B(n_12),
.C(n_13),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_686),
.B(n_14),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_SL g769 ( 
.A(n_686),
.B(n_16),
.C(n_17),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_715),
.A2(n_665),
.B(n_690),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_709),
.B(n_681),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_733),
.B(n_693),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_706),
.A2(n_639),
.B(n_645),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_705),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_759),
.A2(n_643),
.B(n_659),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_733),
.B(n_695),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_707),
.A2(n_655),
.B(n_656),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_710),
.A2(n_672),
.B(n_689),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_722),
.B(n_698),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_725),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_745),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_741),
.B(n_701),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_732),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_760),
.B(n_700),
.C(n_697),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_734),
.A2(n_648),
.B(n_650),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_704),
.Y(n_786)
);

AOI31xp67_ASAP7_75t_L g787 ( 
.A1(n_727),
.A2(n_676),
.A3(n_671),
.B(n_674),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_768),
.A2(n_683),
.B(n_684),
.C(n_685),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_732),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_749),
.A2(n_662),
.B(n_661),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_749),
.A2(n_660),
.B(n_684),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_727),
.A2(n_756),
.B(n_752),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_726),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_726),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_703),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_708),
.A2(n_688),
.B(n_687),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_751),
.A2(n_75),
.B(n_169),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_755),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_729),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_711),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_721),
.A2(n_73),
.B(n_159),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_746),
.Y(n_802)
);

AO31x2_ASAP7_75t_L g803 ( 
.A1(n_723),
.A2(n_16),
.A3(n_18),
.B(n_19),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_761),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_728),
.Y(n_805)
);

BUFx12f_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_767),
.B(n_641),
.C(n_651),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_764),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_724),
.A2(n_72),
.B(n_136),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_756),
.A2(n_68),
.B(n_135),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_736),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_720),
.B(n_21),
.Y(n_812)
);

AO31x2_ASAP7_75t_L g813 ( 
.A1(n_744),
.A2(n_22),
.A3(n_23),
.B(n_24),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_709),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_712),
.B(n_25),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_766),
.A2(n_84),
.B(n_125),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_714),
.B(n_735),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_713),
.A2(n_83),
.B(n_124),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_744),
.A2(n_79),
.B(n_123),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_737),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_806),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_817),
.A2(n_766),
.B1(n_729),
.B2(n_740),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_793),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_781),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_774),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_814),
.A2(n_772),
.B1(n_776),
.B2(n_815),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_771),
.A2(n_743),
.B1(n_735),
.B2(n_722),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_793),
.Y(n_828)
);

INVx6_ASAP7_75t_L g829 ( 
.A(n_793),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_819),
.A2(n_718),
.B1(n_742),
.B2(n_716),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_818),
.A2(n_738),
.B1(n_750),
.B2(n_718),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_794),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_SL g833 ( 
.A1(n_816),
.A2(n_769),
.B1(n_758),
.B2(n_753),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_795),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_779),
.A2(n_820),
.B1(n_816),
.B2(n_782),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_802),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_783),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_779),
.A2(n_738),
.B1(n_762),
.B2(n_763),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_820),
.A2(n_762),
.B1(n_739),
.B2(n_757),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_799),
.A2(n_762),
.B1(n_717),
.B2(n_730),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_786),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_794),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_811),
.A2(n_754),
.B1(n_719),
.B2(n_739),
.Y(n_843)
);

BUFx10_ASAP7_75t_L g844 ( 
.A(n_794),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_804),
.A2(n_736),
.B1(n_762),
.B2(n_765),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_800),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_812),
.A2(n_730),
.B1(n_717),
.B2(n_748),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_805),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_808),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_799),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_SL g852 ( 
.A1(n_804),
.A2(n_765),
.B1(n_28),
.B2(n_29),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_789),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_807),
.Y(n_854)
);

CKINVDCx11_ASAP7_75t_R g855 ( 
.A(n_798),
.Y(n_855)
);

BUFx4f_ASAP7_75t_L g856 ( 
.A(n_811),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_810),
.Y(n_857)
);

BUFx4_ASAP7_75t_SL g858 ( 
.A(n_813),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_803),
.Y(n_859)
);

BUFx2_ASAP7_75t_SL g860 ( 
.A(n_810),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_792),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_809),
.A2(n_748),
.B1(n_747),
.B2(n_29),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_803),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_809),
.Y(n_865)
);

CKINVDCx11_ASAP7_75t_R g866 ( 
.A(n_813),
.Y(n_866)
);

INVx6_ASAP7_75t_L g867 ( 
.A(n_801),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_801),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_790),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_777),
.B(n_748),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_777),
.B(n_27),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_785),
.A2(n_731),
.B1(n_30),
.B2(n_31),
.Y(n_873)
);

CKINVDCx11_ASAP7_75t_R g874 ( 
.A(n_803),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_803),
.Y(n_875)
);

BUFx10_ASAP7_75t_L g876 ( 
.A(n_797),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_775),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_775),
.B(n_773),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_824),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_878),
.A2(n_796),
.B(n_770),
.Y(n_880)
);

BUFx12f_ASAP7_75t_L g881 ( 
.A(n_855),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_859),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_830),
.A2(n_770),
.B(n_788),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_871),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_869),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_864),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_875),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_876),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_858),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_862),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_862),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_870),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_862),
.Y(n_893)
);

OA21x2_ASAP7_75t_L g894 ( 
.A1(n_872),
.A2(n_791),
.B(n_778),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_876),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_858),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_867),
.Y(n_897)
);

CKINVDCx11_ASAP7_75t_R g898 ( 
.A(n_854),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_874),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_856),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_867),
.Y(n_901)
);

BUFx8_ASAP7_75t_SL g902 ( 
.A(n_842),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_834),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_877),
.A2(n_788),
.B1(n_33),
.B2(n_34),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_846),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_850),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_866),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_867),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_853),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_868),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_837),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_877),
.B(n_32),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_860),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_SL g915 ( 
.A1(n_852),
.A2(n_787),
.B1(n_35),
.B2(n_36),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_904),
.A2(n_865),
.B(n_861),
.Y(n_916)
);

NOR2x1_ASAP7_75t_SL g917 ( 
.A(n_900),
.B(n_843),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_903),
.B(n_907),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_904),
.A2(n_827),
.B(n_831),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_884),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_881),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_883),
.A2(n_856),
.B(n_830),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_903),
.B(n_835),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_904),
.A2(n_857),
.B(n_863),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_906),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_903),
.B(n_822),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_903),
.B(n_822),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_892),
.B(n_825),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_913),
.A2(n_915),
.B1(n_908),
.B2(n_852),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_883),
.A2(n_863),
.B(n_833),
.C(n_873),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_898),
.B(n_836),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_892),
.B(n_826),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_883),
.A2(n_913),
.B(n_833),
.C(n_899),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_887),
.B(n_841),
.Y(n_934)
);

AND2x4_ASAP7_75t_SL g935 ( 
.A(n_900),
.B(n_844),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_906),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_907),
.B(n_845),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_898),
.B(n_848),
.Y(n_938)
);

AO32x1_ASAP7_75t_L g939 ( 
.A1(n_913),
.A2(n_845),
.A3(n_832),
.B1(n_826),
.B2(n_851),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_888),
.Y(n_940)
);

NOR2x1_ASAP7_75t_SL g941 ( 
.A(n_900),
.B(n_828),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_907),
.B(n_851),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_887),
.B(n_851),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_911),
.B(n_851),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_907),
.B(n_851),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_913),
.A2(n_838),
.B(n_839),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_915),
.A2(n_911),
.B(n_880),
.Y(n_947)
);

OAI211xp5_ASAP7_75t_L g948 ( 
.A1(n_899),
.A2(n_847),
.B(n_840),
.C(n_821),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_905),
.B(n_851),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_SL g950 ( 
.A1(n_899),
.A2(n_823),
.B(n_821),
.C(n_828),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_905),
.B(n_823),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_900),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_889),
.B(n_828),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_890),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_915),
.A2(n_821),
.B1(n_829),
.B2(n_832),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_900),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_929),
.A2(n_908),
.B1(n_896),
.B2(n_889),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_918),
.B(n_882),
.Y(n_958)
);

NOR2x1p5_ASAP7_75t_L g959 ( 
.A(n_932),
.B(n_908),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_918),
.B(n_882),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_942),
.B(n_882),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_942),
.B(n_886),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_920),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_920),
.B(n_887),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_925),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_SL g967 ( 
.A1(n_919),
.A2(n_908),
.B(n_889),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_925),
.B(n_905),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_945),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_954),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_951),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_945),
.B(n_886),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_934),
.B(n_884),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_949),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_937),
.B(n_886),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_937),
.B(n_880),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_949),
.B(n_880),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_940),
.Y(n_978)
);

OAI222xp33_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_890),
.B1(n_891),
.B2(n_896),
.C1(n_893),
.C2(n_900),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_951),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_923),
.B(n_914),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_916),
.A2(n_893),
.B1(n_897),
.B2(n_901),
.Y(n_982)
);

OAI211xp5_ASAP7_75t_SL g983 ( 
.A1(n_967),
.A2(n_933),
.B(n_930),
.C(n_924),
.Y(n_983)
);

AND2x4_ASAP7_75t_SL g984 ( 
.A(n_958),
.B(n_952),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_978),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_969),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_964),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_969),
.B(n_947),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_958),
.Y(n_989)
);

AO21x2_ASAP7_75t_L g990 ( 
.A1(n_979),
.A2(n_944),
.B(n_895),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_957),
.A2(n_946),
.B1(n_890),
.B2(n_891),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_969),
.B(n_977),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_977),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_961),
.Y(n_994)
);

INVx5_ASAP7_75t_SL g995 ( 
.A(n_979),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_977),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_961),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_981),
.B(n_923),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_976),
.B(n_974),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_958),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_976),
.B(n_940),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_981),
.B(n_926),
.Y(n_1002)
);

OR2x6_ASAP7_75t_L g1003 ( 
.A(n_978),
.B(n_952),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_978),
.B(n_940),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_983),
.A2(n_967),
.B1(n_959),
.B2(n_957),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_959),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_986),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_989),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_985),
.B(n_961),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_1002),
.B(n_973),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_996),
.B(n_976),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_983),
.A2(n_982),
.B(n_955),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_989),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_989),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_987),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_1016),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1010),
.B(n_996),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1015),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1005),
.B(n_988),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1015),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_996),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_1010),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_1011),
.B(n_1002),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1019),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1019),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1020),
.B(n_1007),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_1017),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1025),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1028),
.B(n_1013),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1026),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_991),
.B1(n_1021),
.B2(n_931),
.C(n_921),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_879),
.Y(n_1034)
);

AO21x1_ASAP7_75t_L g1035 ( 
.A1(n_1025),
.A2(n_1021),
.B(n_1018),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1028),
.A2(n_995),
.B1(n_991),
.B2(n_988),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1025),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1025),
.Y(n_1038)
);

INVxp33_ASAP7_75t_L g1039 ( 
.A(n_1028),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_1035),
.A2(n_1022),
.B(n_1018),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1039),
.A2(n_938),
.B(n_879),
.Y(n_1041)
);

OAI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_1036),
.A2(n_1023),
.B1(n_1024),
.B2(n_985),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1029),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1031),
.A2(n_950),
.B(n_1023),
.C(n_1024),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1033),
.A2(n_995),
.B1(n_1023),
.B2(n_1022),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1030),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1034),
.B(n_881),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1037),
.Y(n_1048)
);

OAI32xp33_ASAP7_75t_L g1049 ( 
.A1(n_1038),
.A2(n_987),
.A3(n_995),
.B1(n_993),
.B2(n_1011),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1032),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1033),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1029),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1033),
.A2(n_995),
.B1(n_988),
.B2(n_990),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1039),
.A2(n_948),
.B(n_928),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1029),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_1048),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1041),
.B(n_1012),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_881),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_1040),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1043),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1046),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1051),
.B(n_1012),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1052),
.Y(n_1063)
);

AOI211xp5_ASAP7_75t_L g1064 ( 
.A1(n_1041),
.A2(n_928),
.B(n_934),
.C(n_995),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_1050),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_1044),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1045),
.B(n_1053),
.Y(n_1067)
);

NAND5xp2_ASAP7_75t_L g1068 ( 
.A(n_1054),
.B(n_896),
.C(n_881),
.D(n_902),
.E(n_914),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1054),
.A2(n_939),
.B(n_1008),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1055),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1042),
.B(n_902),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1049),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1043),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1041),
.Y(n_1074)
);

NOR4xp25_ASAP7_75t_L g1075 ( 
.A(n_1059),
.B(n_1008),
.C(n_1006),
.D(n_1014),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_993),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1072),
.B(n_993),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1056),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1065),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1059),
.B(n_995),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1058),
.B(n_987),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_1059),
.B(n_828),
.C(n_985),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1065),
.B(n_987),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_1006),
.Y(n_1084)
);

NAND4xp75_ASAP7_75t_L g1085 ( 
.A(n_1056),
.B(n_995),
.C(n_1009),
.D(n_999),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1057),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1072),
.B(n_993),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1066),
.B(n_993),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1057),
.B(n_993),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1060),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_1061),
.B(n_33),
.C(n_35),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1080),
.A2(n_1067),
.B1(n_1062),
.B2(n_1070),
.C(n_1073),
.Y(n_1092)
);

AOI221x1_ASAP7_75t_L g1093 ( 
.A1(n_1078),
.A2(n_1073),
.B1(n_1070),
.B2(n_1061),
.C(n_1063),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1086),
.B(n_1063),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1081),
.A2(n_1071),
.B1(n_1064),
.B2(n_1069),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_1083),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1079),
.B(n_998),
.Y(n_1097)
);

NAND4xp25_ASAP7_75t_SL g1098 ( 
.A(n_1077),
.B(n_1068),
.C(n_973),
.D(n_999),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_SL g1099 ( 
.A(n_1091),
.B(n_829),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_952),
.C(n_901),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_1089),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_1090),
.B(n_36),
.Y(n_1102)
);

AOI321xp33_ASAP7_75t_L g1103 ( 
.A1(n_1075),
.A2(n_953),
.A3(n_890),
.B1(n_891),
.B2(n_966),
.C(n_914),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1082),
.B(n_985),
.C(n_963),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_1088),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1076),
.A2(n_939),
.B(n_941),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_SL g1107 ( 
.A1(n_1087),
.A2(n_37),
.B(n_38),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_1084),
.A2(n_37),
.B(n_38),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1085),
.A2(n_985),
.B(n_963),
.Y(n_1109)
);

AOI211xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1078),
.A2(n_953),
.B(n_966),
.C(n_42),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1086),
.B(n_992),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1086),
.A2(n_984),
.B1(n_1003),
.B2(n_953),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1086),
.A2(n_984),
.B1(n_1003),
.B2(n_990),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_1081),
.A2(n_984),
.B(n_1003),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1086),
.A2(n_984),
.B1(n_1003),
.B2(n_990),
.Y(n_1115)
);

AO22x2_ASAP7_75t_L g1116 ( 
.A1(n_1093),
.A2(n_986),
.B1(n_997),
.B2(n_994),
.Y(n_1116)
);

OAI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_1092),
.A2(n_1095),
.B1(n_1094),
.B2(n_1114),
.C(n_1105),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1101),
.Y(n_1118)
);

OAI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1110),
.A2(n_1003),
.B1(n_956),
.B2(n_964),
.C(n_985),
.Y(n_1119)
);

AOI211xp5_ASAP7_75t_L g1120 ( 
.A1(n_1108),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_1120)
);

AOI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1096),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1098),
.A2(n_990),
.B1(n_974),
.B2(n_970),
.C(n_986),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1101),
.B(n_999),
.Y(n_1123)
);

OAI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1100),
.A2(n_1003),
.B1(n_956),
.B2(n_985),
.C(n_891),
.Y(n_1124)
);

OAI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1112),
.A2(n_985),
.B1(n_1003),
.B2(n_956),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1101),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1099),
.Y(n_1127)
);

OAI211xp5_ASAP7_75t_L g1128 ( 
.A1(n_1107),
.A2(n_985),
.B(n_47),
.C(n_46),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1102),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1097),
.A2(n_990),
.B1(n_970),
.B2(n_1004),
.C(n_1001),
.Y(n_1130)
);

OAI221xp5_ASAP7_75t_L g1131 ( 
.A1(n_1109),
.A2(n_1003),
.B1(n_956),
.B2(n_985),
.C(n_829),
.Y(n_1131)
);

AOI211xp5_ASAP7_75t_L g1132 ( 
.A1(n_1111),
.A2(n_1004),
.B(n_1001),
.C(n_965),
.Y(n_1132)
);

AOI222xp33_ASAP7_75t_L g1133 ( 
.A1(n_1104),
.A2(n_917),
.B1(n_941),
.B2(n_1001),
.C1(n_1000),
.C2(n_1004),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1113),
.A2(n_50),
.B(n_51),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1103),
.B(n_965),
.C(n_840),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1106),
.B(n_968),
.C(n_895),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1115),
.A2(n_997),
.B(n_994),
.C(n_1000),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1098),
.A2(n_956),
.B1(n_935),
.B2(n_897),
.Y(n_1138)
);

XOR2xp5_ASAP7_75t_L g1139 ( 
.A(n_1095),
.B(n_917),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1126),
.B(n_1004),
.Y(n_1140)
);

NOR4xp25_ASAP7_75t_L g1141 ( 
.A(n_1117),
.B(n_968),
.C(n_1000),
.D(n_994),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1118),
.B(n_895),
.C(n_1004),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1128),
.B(n_54),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1129),
.A2(n_1004),
.B1(n_935),
.B2(n_975),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1127),
.B(n_997),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1120),
.B(n_997),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1123),
.B(n_994),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_L g1148 ( 
.A(n_1139),
.B(n_992),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1116),
.Y(n_1149)
);

NOR2x1_ASAP7_75t_L g1150 ( 
.A(n_1119),
.B(n_992),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1121),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1138),
.A2(n_975),
.B1(n_980),
.B2(n_972),
.Y(n_1152)
);

NAND4xp75_ASAP7_75t_L g1153 ( 
.A(n_1122),
.B(n_975),
.C(n_844),
.D(n_972),
.Y(n_1153)
);

NOR2x1_ASAP7_75t_L g1154 ( 
.A(n_1136),
.B(n_888),
.Y(n_1154)
);

NOR2x1_ASAP7_75t_L g1155 ( 
.A(n_1131),
.B(n_888),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1116),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1134),
.B(n_980),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1135),
.B(n_888),
.Y(n_1158)
);

AND2x2_ASAP7_75t_SL g1159 ( 
.A(n_1130),
.B(n_909),
.Y(n_1159)
);

XOR2xp5_ASAP7_75t_L g1160 ( 
.A(n_1125),
.B(n_55),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1137),
.B(n_895),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1151),
.B(n_1133),
.C(n_1124),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1156),
.B(n_1132),
.C(n_909),
.Y(n_1163)
);

AOI322xp5_ASAP7_75t_L g1164 ( 
.A1(n_1148),
.A2(n_971),
.A3(n_884),
.B1(n_962),
.B2(n_972),
.C1(n_939),
.C2(n_926),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1149),
.B(n_888),
.C(n_909),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1143),
.B(n_962),
.Y(n_1166)
);

XNOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1141),
.B(n_57),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1160),
.B(n_909),
.C(n_943),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_L g1169 ( 
.A(n_1146),
.B(n_897),
.C(n_901),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1140),
.A2(n_939),
.B(n_888),
.Y(n_1170)
);

NAND3x1_ASAP7_75t_SL g1171 ( 
.A(n_1158),
.B(n_59),
.C(n_60),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1145),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1157),
.Y(n_1173)
);

NAND4xp25_ASAP7_75t_L g1174 ( 
.A(n_1155),
.B(n_897),
.C(n_901),
.D(n_927),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_L g1175 ( 
.A(n_1157),
.B(n_897),
.C(n_901),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1142),
.Y(n_1176)
);

AOI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_1159),
.B1(n_1154),
.B2(n_1161),
.C1(n_1150),
.C2(n_1147),
.Y(n_1177)
);

OAI222xp33_ASAP7_75t_L g1178 ( 
.A1(n_1173),
.A2(n_1176),
.B1(n_1167),
.B2(n_1172),
.C1(n_1166),
.C2(n_1144),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1175),
.B(n_1152),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1162),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1165),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1168),
.A2(n_1153),
.B1(n_962),
.B2(n_901),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1171),
.Y(n_1183)
);

INVxp33_ASAP7_75t_SL g1184 ( 
.A(n_1169),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1174),
.Y(n_1185)
);

NOR3xp33_ASAP7_75t_L g1186 ( 
.A(n_1170),
.B(n_897),
.C(n_910),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1164),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1162),
.A2(n_943),
.B1(n_910),
.B2(n_912),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1173),
.A2(n_910),
.B(n_912),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1163),
.A2(n_910),
.B1(n_912),
.B2(n_960),
.C(n_927),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1173),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1180),
.A2(n_912),
.B1(n_960),
.B2(n_894),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1187),
.A2(n_1183),
.B1(n_1191),
.B2(n_1185),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1181),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1179),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1177),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1184),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1186),
.A2(n_960),
.B1(n_894),
.B2(n_885),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1182),
.A2(n_894),
.B1(n_65),
.B2(n_67),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1190),
.A2(n_894),
.B1(n_885),
.B2(n_87),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1188),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1196),
.A2(n_1189),
.B1(n_1178),
.B2(n_894),
.Y(n_1202)
);

OAI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1193),
.A2(n_894),
.B1(n_86),
.B2(n_89),
.Y(n_1203)
);

XOR2x1_ASAP7_75t_L g1204 ( 
.A(n_1195),
.B(n_64),
.Y(n_1204)
);

OR3x1_ASAP7_75t_L g1205 ( 
.A(n_1194),
.B(n_93),
.C(n_95),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1197),
.B(n_96),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1201),
.A2(n_894),
.B1(n_885),
.B2(n_102),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1206),
.A2(n_1199),
.B(n_1192),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1204),
.B(n_1198),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1205),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1203),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1209),
.A2(n_1202),
.B(n_1207),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1212),
.Y(n_1213)
);

XOR2xp5_ASAP7_75t_L g1214 ( 
.A(n_1213),
.B(n_1210),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1214),
.Y(n_1215)
);

OAI221xp5_ASAP7_75t_R g1216 ( 
.A1(n_1215),
.A2(n_1211),
.B1(n_1208),
.B2(n_1200),
.C(n_105),
.Y(n_1216)
);

AOI211xp5_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_98),
.B(n_99),
.C(n_103),
.Y(n_1217)
);


endmodule