module fake_jpeg_10112_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2x1_ASAP7_75t_R g43 ( 
.A(n_40),
.B(n_20),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_77),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_23),
.B1(n_42),
.B2(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_52),
.B1(n_42),
.B2(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_16),
.B1(n_25),
.B2(n_74),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_89),
.B1(n_97),
.B2(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_54),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_98),
.Y(n_118)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_99),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_48),
.B1(n_53),
.B2(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_81),
.B1(n_75),
.B2(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_16),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_62),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_115),
.C(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_13),
.C(n_14),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_125),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_71),
.C(n_45),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_76),
.B(n_78),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_103),
.B(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_98),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_23),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_106),
.C(n_23),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_87),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_141),
.C(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_135),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_105),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_99),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_105),
.B1(n_97),
.B2(n_89),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_128),
.B1(n_147),
.B2(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_44),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_47),
.C(n_95),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_76),
.C(n_79),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_116),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_163),
.C(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_122),
.B1(n_117),
.B2(n_139),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_160),
.B1(n_78),
.B2(n_7),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_133),
.C(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_6),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_117),
.B1(n_109),
.B2(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_72),
.C(n_82),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_23),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_23),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_132),
.B1(n_145),
.B2(n_141),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_170),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_160),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_0),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_6),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_157),
.B1(n_150),
.B2(n_3),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_149),
.C(n_152),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_193),
.C(n_5),
.Y(n_201)
);

AOI321xp33_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_152),
.A3(n_162),
.B1(n_165),
.B2(n_159),
.C(n_164),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_177),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_1),
.CI(n_4),
.CON(n_192),
.SN(n_192)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_8),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_10),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_172),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_195),
.B(n_199),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_167),
.B(n_170),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_176),
.B(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_201),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_192),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_190),
.B(n_184),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_182),
.B(n_187),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_195),
.B(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_213),
.C(n_8),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_204),
.B(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_13),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_10),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

OAI311xp33_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_218),
.A3(n_219),
.B1(n_12),
.C1(n_11),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_222),
.B(n_12),
.C(n_1),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule