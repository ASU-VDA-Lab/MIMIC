module fake_ariane_2659_n_1390 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1390);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1390;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_1121;
wire n_461;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

INVxp67_ASAP7_75t_L g310 ( 
.A(n_110),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_224),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_132),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_176),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_11),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_137),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_127),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_188),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_126),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_104),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_243),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_212),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_118),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_218),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_163),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_113),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_260),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_292),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_152),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_65),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_150),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_264),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_13),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_189),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_194),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_167),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_42),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_97),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_3),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_47),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_123),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_74),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_299),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_85),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_35),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_38),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_205),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_280),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_147),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_50),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_304),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_275),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_98),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_209),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_265),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_286),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_293),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_155),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_219),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_186),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_254),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_273),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_228),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_87),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_195),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_111),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_169),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_211),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_2),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_86),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_139),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_282),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_102),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_203),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_236),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_16),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_56),
.B(n_73),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_138),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_160),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_200),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_285),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_92),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_266),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_231),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_287),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_24),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_172),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_133),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_128),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_262),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_165),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_112),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_206),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_121),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_81),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_28),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_301),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_75),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_53),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_168),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_100),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_134),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_302),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_234),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_252),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_20),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_261),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_18),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_197),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_276),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_1),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_114),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_143),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_269),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_106),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_233),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_199),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_36),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_181),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_216),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_309),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_283),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_32),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_140),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_290),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_149),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_193),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_294),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_250),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_96),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_124),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_105),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_235),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_229),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_153),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_31),
.B(n_291),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_24),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_103),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_198),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_40),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_135),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_129),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_42),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_178),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_210),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_237),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_170),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_45),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_38),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_159),
.Y(n_461)
);

INVxp33_ASAP7_75t_R g462 ( 
.A(n_156),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_222),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_14),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_145),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_183),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_142),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_136),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_277),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_162),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_249),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_204),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_232),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_84),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_247),
.Y(n_475)
);

BUFx5_ASAP7_75t_L g476 ( 
.A(n_1),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_41),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_180),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_297),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_7),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_29),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_151),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_308),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_213),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_240),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_305),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_161),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_109),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_177),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_148),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_158),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_90),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_6),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_49),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_201),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_255),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_91),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_154),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_274),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_239),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_196),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_131),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_130),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_306),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_202),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_175),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_44),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_267),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_48),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_241),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_215),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_108),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_248),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_190),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_226),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_125),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_217),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_253),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_69),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_214),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_303),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_166),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_296),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_94),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_173),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_50),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_182),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_208),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_89),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_238),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_11),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_17),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_284),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_21),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_227),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_174),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_53),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_60),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_242),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_58),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_220),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_120),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_363),
.Y(n_543)
);

OAI22x1_ASAP7_75t_L g544 ( 
.A1(n_451),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_544)
);

NOR2x1_ASAP7_75t_L g545 ( 
.A(n_342),
.B(n_55),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_341),
.Y(n_546)
);

OAI22x1_ASAP7_75t_SL g547 ( 
.A1(n_417),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_354),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_354),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_344),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_362),
.A2(n_59),
.B(n_57),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_469),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_316),
.B(n_5),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_313),
.A2(n_7),
.B(n_8),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_316),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_379),
.A2(n_62),
.B(n_61),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_343),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_383),
.B(n_8),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_383),
.B(n_542),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_314),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_9),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_451),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_480),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_315),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_469),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_354),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_415),
.B(n_10),
.Y(n_570)
);

BUFx8_ASAP7_75t_SL g571 ( 
.A(n_434),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_354),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_354),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_436),
.B(n_13),
.Y(n_574)
);

OA21x2_ASAP7_75t_L g575 ( 
.A1(n_317),
.A2(n_14),
.B(n_15),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_484),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_476),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_326),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_342),
.B(n_364),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

BUFx12f_ASAP7_75t_L g582 ( 
.A(n_371),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_322),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_315),
.Y(n_584)
);

CKINVDCx6p67_ASAP7_75t_R g585 ( 
.A(n_371),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_476),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_315),
.Y(n_587)
);

AOI22x1_ASAP7_75t_SL g588 ( 
.A1(n_429),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_412),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_476),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_364),
.B(n_19),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_22),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_319),
.B(n_22),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_484),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_351),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_336),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_323),
.B(n_23),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_376),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_412),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_484),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_484),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_315),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_332),
.B(n_23),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_25),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_389),
.A2(n_64),
.B(n_63),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_384),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_402),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_402),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_402),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_535),
.B(n_25),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_480),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_437),
.B(n_26),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_370),
.A2(n_490),
.B1(n_361),
.B2(n_367),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_311),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_402),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_505),
.B(n_26),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_391),
.B(n_27),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_349),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_505),
.Y(n_619)
);

OA21x2_ASAP7_75t_L g620 ( 
.A1(n_333),
.A2(n_27),
.B(n_28),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_459),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_350),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_395),
.B(n_29),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_396),
.Y(n_624)
);

CKINVDCx6p67_ASAP7_75t_R g625 ( 
.A(n_355),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_340),
.B(n_30),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_377),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_459),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_346),
.B(n_30),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_419),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_440),
.A2(n_67),
.B(n_66),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_459),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_399),
.B(n_31),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_459),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_373),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_477),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_507),
.B(n_33),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_435),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_531),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_452),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_353),
.B(n_36),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_374),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_407),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_345),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_359),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_410),
.B(n_37),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_365),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_422),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_369),
.Y(n_650)
);

BUFx12f_ASAP7_75t_L g651 ( 
.A(n_448),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_378),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_382),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_387),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_393),
.Y(n_655)
);

BUFx12f_ASAP7_75t_L g656 ( 
.A(n_454),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_460),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_397),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_398),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_474),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_464),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_400),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_406),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_408),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_380),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_420),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_423),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_426),
.Y(n_668)
);

BUFx8_ASAP7_75t_SL g669 ( 
.A(n_504),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_433),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_481),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_493),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_447),
.B(n_68),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_388),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_494),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_442),
.Y(n_676)
);

OAI22x1_ASAP7_75t_SL g677 ( 
.A1(n_509),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_462),
.B(n_43),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_443),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_445),
.Y(n_680)
);

BUFx8_ASAP7_75t_SL g681 ( 
.A(n_511),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_449),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_455),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_463),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_472),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_409),
.B(n_45),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_312),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_526),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_516),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_473),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_537),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_475),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_457),
.B(n_46),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_478),
.B(n_49),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_521),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_467),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_488),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_525),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_583),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_549),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_621),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_489),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_643),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_669),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_549),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_681),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_613),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_595),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_695),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_578),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_625),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_550),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_571),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_578),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_581),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_559),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_621),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_581),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_644),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_567),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_638),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_590),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_698),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_585),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_599),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_543),
.B(n_432),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_627),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_580),
.B(n_458),
.Y(n_728)
);

XOR2xp5_ASAP7_75t_L g729 ( 
.A(n_678),
.B(n_320),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_618),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_651),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_656),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_582),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_L g736 ( 
.A(n_589),
.B(n_310),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_619),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_621),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_572),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_554),
.B(n_310),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_614),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_614),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_687),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_687),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_657),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_661),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_671),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_691),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_573),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_622),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_R g751 ( 
.A(n_655),
.B(n_321),
.Y(n_751)
);

AND3x2_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_318),
.C(n_483),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_672),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_598),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_675),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_553),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_632),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_649),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_688),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_616),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_658),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_564),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_624),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_659),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_630),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_632),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_641),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_664),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_690),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_565),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_638),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_640),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_640),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_584),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_662),
.B(n_324),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_640),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_587),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_645),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_R g781 ( 
.A(n_556),
.B(n_325),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_645),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_645),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_566),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_611),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_587),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_665),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_665),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_607),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_SL g790 ( 
.A1(n_562),
.A2(n_318),
.B1(n_538),
.B2(n_495),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_636),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_665),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_674),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_674),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_663),
.B(n_541),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_561),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_636),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_700),
.B(n_705),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_762),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_728),
.B(n_686),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_767),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_792),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_710),
.B(n_548),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_741),
.B(n_574),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_742),
.B(n_674),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_799),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_577),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_715),
.B(n_586),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_673),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_743),
.B(n_673),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_767),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_722),
.A2(n_558),
.B(n_551),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_725),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_755),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_744),
.B(n_570),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_764),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_766),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_720),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_765),
.B(n_686),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_770),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_716),
.B(n_579),
.C(n_593),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_739),
.B(n_667),
.Y(n_825)
);

BUFx6f_ASAP7_75t_SL g826 ( 
.A(n_740),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_733),
.B(n_749),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_769),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_789),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_732),
.B(n_670),
.Y(n_830)
);

BUFx2_ASAP7_75t_R g831 ( 
.A(n_713),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_776),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_779),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_702),
.B(n_673),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_SL g835 ( 
.A(n_707),
.B(n_673),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_732),
.B(n_676),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_771),
.B(n_591),
.Y(n_837)
);

AO221x1_ASAP7_75t_L g838 ( 
.A1(n_712),
.A2(n_544),
.B1(n_606),
.B2(n_588),
.C(n_677),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_726),
.B(n_546),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_763),
.B(n_604),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_763),
.B(n_647),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_786),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_757),
.B(n_604),
.Y(n_843)
);

NOR3xp33_ASAP7_75t_L g844 ( 
.A(n_719),
.B(n_603),
.C(n_597),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_724),
.B(n_610),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_791),
.B(n_637),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_702),
.B(n_650),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_721),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_701),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_759),
.B(n_653),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_790),
.B(n_679),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_793),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_783),
.B(n_623),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_760),
.B(n_637),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_701),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_745),
.B(n_626),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_736),
.B(n_617),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_751),
.A2(n_631),
.B(n_605),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_773),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_784),
.B(n_546),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_701),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_777),
.B(n_797),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_717),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_774),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_780),
.B(n_682),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_781),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_717),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_730),
.B(n_685),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_782),
.B(n_697),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_708),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_787),
.B(n_693),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_775),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_788),
.B(n_633),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_794),
.B(n_795),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_746),
.B(n_696),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_796),
.B(n_552),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_747),
.B(n_646),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_778),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_717),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_738),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_723),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_748),
.B(n_646),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_738),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_753),
.B(n_646),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_738),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_758),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_752),
.B(n_552),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_756),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_758),
.B(n_560),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_648),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_798),
.B(n_648),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_758),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_875),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_870),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_866),
.B(n_727),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_816),
.B(n_617),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_835),
.A2(n_761),
.B1(n_729),
.B2(n_642),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_801),
.B(n_823),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_881),
.B(n_711),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_804),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_849),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_821),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_850),
.B(n_731),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_813),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_817),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_888),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_831),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_890),
.B(n_734),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_847),
.B(n_839),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_872),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_849),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_847),
.B(n_629),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_849),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_841),
.B(n_563),
.Y(n_915)
);

AO22x1_ASAP7_75t_L g916 ( 
.A1(n_824),
.A2(n_703),
.B1(n_706),
.B2(n_704),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_857),
.B(n_639),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_819),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_820),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_818),
.B(n_891),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_828),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_SL g922 ( 
.A1(n_802),
.A2(n_660),
.B(n_635),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_800),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_860),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_840),
.B(n_639),
.Y(n_926)
);

OR2x2_ASAP7_75t_SL g927 ( 
.A(n_838),
.B(n_547),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_835),
.A2(n_694),
.B1(n_689),
.B2(n_592),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_800),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_830),
.B(n_735),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_854),
.B(n_750),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_SL g932 ( 
.A(n_844),
.B(n_785),
.C(n_772),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_836),
.A2(n_856),
.B1(n_834),
.B2(n_826),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_884),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_833),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_842),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_883),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_877),
.B(n_737),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_827),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_857),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_882),
.B(n_648),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_868),
.B(n_845),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_883),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_827),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_829),
.Y(n_945)
);

AND2x2_ASAP7_75t_SL g946 ( 
.A(n_845),
.B(n_555),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_859),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_832),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_652),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_803),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_855),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_848),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_SL g953 ( 
.A1(n_864),
.A2(n_699),
.B1(n_588),
.B2(n_575),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_825),
.B(n_652),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_861),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_807),
.B(n_851),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_851),
.B(n_652),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_871),
.B(n_654),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_814),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_862),
.B(n_654),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_871),
.B(n_654),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_865),
.B(n_869),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_805),
.A2(n_668),
.B1(n_680),
.B2(n_666),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_873),
.B(n_865),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_852),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_834),
.A2(n_575),
.B1(n_620),
.B2(n_555),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_863),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_867),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_811),
.A2(n_545),
.B(n_620),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_887),
.B(n_837),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_869),
.B(n_666),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_846),
.B(n_696),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_878),
.Y(n_973)
);

NOR2x1p5_ASAP7_75t_L g974 ( 
.A(n_874),
.B(n_666),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_806),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_805),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_853),
.B(n_876),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_809),
.B(n_810),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_822),
.B(n_668),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_809),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_810),
.Y(n_981)
);

CKINVDCx6p67_ASAP7_75t_R g982 ( 
.A(n_889),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_SL g983 ( 
.A1(n_811),
.A2(n_501),
.B1(n_503),
.B2(n_492),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_889),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_879),
.B(n_668),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_880),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_812),
.B(n_680),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_886),
.A2(n_506),
.B(n_515),
.C(n_514),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_885),
.B(n_680),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_892),
.A2(n_684),
.B1(n_692),
.B2(n_683),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_978),
.A2(n_815),
.B(n_858),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_903),
.Y(n_992)
);

OR2x6_ASAP7_75t_SL g993 ( 
.A(n_894),
.B(n_327),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_939),
.A2(n_520),
.B(n_524),
.C(n_517),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_913),
.A2(n_815),
.B(n_858),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_923),
.A2(n_329),
.B(n_328),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_911),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_934),
.B(n_683),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_944),
.B(n_683),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_929),
.A2(n_540),
.B(n_529),
.C(n_491),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_933),
.B(n_684),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_924),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_962),
.B(n_684),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_910),
.B(n_692),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_969),
.A2(n_385),
.B(n_485),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_928),
.A2(n_980),
.B1(n_981),
.B2(n_976),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_924),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_SL g1009 ( 
.A(n_947),
.B(n_331),
.C(n_330),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_965),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_928),
.A2(n_518),
.B(n_523),
.C(n_497),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_964),
.A2(n_335),
.B(n_334),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_987),
.A2(n_533),
.B(n_608),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_945),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_920),
.A2(n_608),
.B(n_615),
.C(n_609),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_958),
.A2(n_949),
.B(n_984),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_933),
.B(n_692),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_956),
.A2(n_609),
.B(n_615),
.C(n_602),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_942),
.B(n_560),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_957),
.A2(n_628),
.B(n_594),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_897),
.B(n_926),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_973),
.A2(n_54),
.B(n_51),
.C(n_52),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_908),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_900),
.A2(n_902),
.B1(n_906),
.B2(n_905),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_932),
.B(n_922),
.C(n_898),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_917),
.B(n_594),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_907),
.B(n_337),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_899),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_922),
.A2(n_339),
.B(n_347),
.C(n_338),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_915),
.B(n_348),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_896),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_918),
.B(n_352),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_975),
.B(n_356),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_SL g1034 ( 
.A(n_931),
.B(n_358),
.C(n_357),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_948),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_919),
.A2(n_366),
.B1(n_368),
.B2(n_360),
.Y(n_1036)
);

AO21x1_ASAP7_75t_L g1037 ( 
.A1(n_954),
.A2(n_568),
.B(n_557),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_896),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_926),
.B(n_921),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_961),
.A2(n_375),
.B(n_372),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_924),
.Y(n_1041)
);

INVx3_ASAP7_75t_SL g1042 ( 
.A(n_896),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_917),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_940),
.B(n_381),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_925),
.B(n_768),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_917),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_970),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_946),
.A2(n_634),
.B1(n_466),
.B2(n_465),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_935),
.B(n_936),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_968),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_977),
.B(n_386),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_952),
.B(n_768),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_983),
.B(n_390),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_971),
.A2(n_568),
.B(n_557),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_970),
.Y(n_1055)
);

OAI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_904),
.A2(n_456),
.B1(n_394),
.B2(n_539),
.C(n_536),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_960),
.A2(n_912),
.B(n_901),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_989),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_972),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_901),
.A2(n_401),
.B(n_392),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_972),
.B(n_403),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_930),
.B(n_404),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_982),
.B(n_912),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_L g1064 ( 
.A(n_974),
.B(n_405),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_970),
.B(n_634),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_950),
.B(n_411),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_988),
.A2(n_51),
.B(n_52),
.C(n_54),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_914),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_914),
.B(n_413),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_991),
.A2(n_966),
.B(n_955),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_995),
.A2(n_937),
.B1(n_943),
.B2(n_959),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1006),
.A2(n_966),
.B(n_979),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1005),
.A2(n_955),
.B(n_951),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1047),
.B(n_937),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_1006),
.A2(n_967),
.B(n_963),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_1050),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1016),
.A2(n_941),
.B(n_943),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1020),
.A2(n_895),
.B(n_909),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1010),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_997),
.Y(n_1080)
);

BUFx2_ASAP7_75t_SL g1081 ( 
.A(n_1023),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1007),
.Y(n_1082)
);

INVx8_ASAP7_75t_L g1083 ( 
.A(n_1026),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1042),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_1031),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1039),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_1038),
.B(n_916),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1049),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_SL g1089 ( 
.A1(n_1024),
.A2(n_990),
.B(n_953),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1043),
.B(n_986),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1013),
.A2(n_986),
.B(n_985),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_1026),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_1002),
.B(n_968),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1035),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_1037),
.A2(n_416),
.B(n_414),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1063),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1014),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1024),
.Y(n_1098)
);

AO21x2_ASAP7_75t_L g1099 ( 
.A1(n_1001),
.A2(n_938),
.B(n_968),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_1017),
.A2(n_568),
.B(n_557),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1046),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_993),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_1028),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1054),
.A2(n_70),
.B(n_71),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1021),
.B(n_927),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_992),
.Y(n_1107)
);

BUFx2_ASAP7_75t_SL g1108 ( 
.A(n_1059),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1026),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_1055),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1050),
.Y(n_1111)
);

CKINVDCx6p67_ASAP7_75t_R g1112 ( 
.A(n_1065),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1002),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1057),
.A2(n_72),
.B(n_76),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1008),
.Y(n_1115)
);

AOI22x1_ASAP7_75t_L g1116 ( 
.A1(n_996),
.A2(n_482),
.B1(n_421),
.B2(n_424),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1025),
.B(n_634),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_1065),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1029),
.A2(n_425),
.B(n_418),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_999),
.A2(n_77),
.B(n_78),
.Y(n_1120)
);

BUFx2_ASAP7_75t_R g1121 ( 
.A(n_1053),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_1003),
.A2(n_600),
.B(n_576),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1004),
.A2(n_79),
.B(n_80),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1018),
.A2(n_428),
.B(n_427),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_998),
.B(n_430),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1058),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1019),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1011),
.A2(n_438),
.B(n_431),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1030),
.B(n_439),
.Y(n_1129)
);

BUFx4_ASAP7_75t_SL g1130 ( 
.A(n_1044),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1015),
.A2(n_600),
.B(n_576),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1068),
.Y(n_1133)
);

INVx6_ASAP7_75t_SL g1134 ( 
.A(n_1064),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1094),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1083),
.B(n_1045),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1071),
.A2(n_1068),
.B(n_1051),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1097),
.Y(n_1138)
);

OAI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1129),
.A2(n_1034),
.B(n_1032),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1079),
.Y(n_1140)
);

BUFx8_ASAP7_75t_L g1141 ( 
.A(n_1103),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1126),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1076),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1089),
.A2(n_1048),
.B1(n_1061),
.B2(n_1062),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1105),
.A2(n_1032),
.B1(n_1009),
.B2(n_1036),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1106),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1070),
.A2(n_1066),
.B(n_1012),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1102),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1107),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1092),
.B(n_1041),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1086),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1086),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1085),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1127),
.A2(n_1036),
.B1(n_1033),
.B2(n_1056),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1073),
.A2(n_994),
.B(n_1069),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1098),
.B(n_1000),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1088),
.A2(n_1027),
.B1(n_1022),
.B2(n_1060),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1080),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1129),
.A2(n_1040),
.B1(n_500),
.B2(n_499),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1082),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1072),
.A2(n_1067),
.B1(n_601),
.B2(n_600),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1096),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1072),
.A2(n_601),
.B1(n_576),
.B2(n_530),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1074),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1119),
.A2(n_601),
.B1(n_528),
.B2(n_527),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1092),
.B(n_82),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1099),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1074),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1119),
.A2(n_522),
.B1(n_519),
.B2(n_513),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1125),
.A2(n_1118),
.B1(n_1084),
.B2(n_1112),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1134),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1075),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1109),
.A2(n_512),
.B1(n_510),
.B2(n_508),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1078),
.A2(n_444),
.B(n_441),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1110),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1113),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1113),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1117),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1077),
.A2(n_502),
.B(n_498),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_1083),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1115),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1077),
.A2(n_83),
.B(n_88),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1130),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1084),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1106),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1128),
.A2(n_496),
.B(n_487),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1115),
.Y(n_1189)
);

OAI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_1128),
.A2(n_486),
.B(n_479),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1122),
.A2(n_471),
.B(n_470),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1114),
.A2(n_93),
.B(n_95),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1188),
.B(n_1101),
.C(n_1090),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_R g1194 ( 
.A(n_1185),
.B(n_1173),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1135),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1162),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1177),
.B(n_1087),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1177),
.B(n_1108),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1182),
.Y(n_1199)
);

INVx8_ASAP7_75t_L g1200 ( 
.A(n_1154),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1184),
.A2(n_1137),
.B(n_1192),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_R g1202 ( 
.A(n_1185),
.B(n_1131),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1138),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1171),
.A2(n_1124),
.B(n_1095),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1160),
.B(n_1121),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_R g1206 ( 
.A(n_1168),
.B(n_1111),
.Y(n_1206)
);

XNOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1148),
.B(n_1081),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1169),
.A2(n_1132),
.A3(n_1100),
.B(n_1091),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1144),
.A2(n_1134),
.B1(n_1124),
.B2(n_1116),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_1148),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1152),
.B(n_1111),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1142),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1140),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1174),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1153),
.B(n_1106),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1182),
.B(n_1133),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1166),
.B(n_1113),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1150),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1145),
.B(n_1133),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1143),
.Y(n_1220)
);

XOR2x2_ASAP7_75t_SL g1221 ( 
.A(n_1175),
.B(n_1093),
.Y(n_1221)
);

INVxp33_ASAP7_75t_L g1222 ( 
.A(n_1164),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1182),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1141),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_R g1225 ( 
.A(n_1168),
.B(n_1123),
.Y(n_1225)
);

AO32x2_ASAP7_75t_L g1226 ( 
.A1(n_1186),
.A2(n_1132),
.A3(n_1100),
.B1(n_1120),
.B2(n_1104),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1171),
.A2(n_1093),
.B(n_468),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1170),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1157),
.A2(n_99),
.A3(n_101),
.B(n_107),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1144),
.A2(n_461),
.B1(n_453),
.B2(n_450),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1145),
.B(n_446),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1183),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1157),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1178),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1172),
.B(n_1149),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1179),
.Y(n_1236)
);

AND2x6_ASAP7_75t_L g1237 ( 
.A(n_1180),
.B(n_115),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1189),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1141),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1188),
.A2(n_1139),
.B(n_1190),
.C(n_1155),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1159),
.B(n_116),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1167),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1159),
.B(n_141),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1233),
.Y(n_1244)
);

OAI221xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1240),
.A2(n_1165),
.B1(n_1163),
.B2(n_1158),
.C(n_1161),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1196),
.B(n_1181),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1212),
.B(n_1218),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1214),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1214),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1232),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1231),
.A2(n_1165),
.B(n_1163),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1238),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_1206),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1201),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1198),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1210),
.B(n_1182),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1215),
.B(n_1211),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1195),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1219),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1203),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1229),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1228),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1197),
.B(n_1191),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1236),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1205),
.B(n_1147),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1235),
.B(n_1147),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1213),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1204),
.A2(n_1230),
.B1(n_1193),
.B2(n_1209),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1234),
.B(n_1146),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1187),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1220),
.B(n_1187),
.Y(n_1272)
);

OR2x4_ASAP7_75t_L g1273 ( 
.A(n_1199),
.B(n_1176),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1199),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1217),
.B(n_1156),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1208),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1223),
.B(n_1151),
.Y(n_1277)
);

AND2x4_ASAP7_75t_SL g1278 ( 
.A(n_1223),
.B(n_1151),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1223),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1241),
.B(n_1158),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1216),
.B(n_1136),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1208),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1216),
.B(n_1136),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1226),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1237),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1226),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1237),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1221),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1243),
.B(n_144),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1266),
.B(n_1222),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1264),
.B(n_1207),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1252),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1248),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1257),
.B(n_1224),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1266),
.B(n_1239),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1247),
.B(n_1200),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1262),
.B(n_1200),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1265),
.B(n_1242),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1255),
.B(n_1227),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1265),
.B(n_1225),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1249),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1250),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1254),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1249),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1245),
.B(n_1194),
.C(n_1202),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1244),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1246),
.B(n_146),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1258),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1280),
.B(n_157),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1259),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1260),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1267),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1267),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1275),
.B(n_179),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1311),
.B(n_1263),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1293),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1291),
.B(n_1275),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1301),
.B(n_1284),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1296),
.B(n_1256),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1303),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1304),
.B(n_1285),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1306),
.B(n_1268),
.C(n_1251),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1307),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1296),
.B(n_1253),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1304),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1299),
.B(n_1254),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1294),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1304),
.B(n_1288),
.Y(n_1329)
);

OAI211xp5_ASAP7_75t_L g1330 ( 
.A1(n_1323),
.A2(n_1289),
.B(n_1310),
.C(n_1292),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1327),
.B(n_1286),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1316),
.B(n_1300),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1319),
.B(n_1294),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1318),
.B(n_1295),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1327),
.B(n_1297),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1325),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1317),
.Y(n_1337)
);

NAND4xp25_ASAP7_75t_L g1338 ( 
.A(n_1321),
.B(n_1298),
.C(n_1315),
.D(n_1308),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1330),
.A2(n_1290),
.B(n_1261),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1336),
.B(n_1320),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1337),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1334),
.A2(n_1329),
.B1(n_1322),
.B2(n_1281),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1332),
.B(n_1322),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1338),
.A2(n_1326),
.B(n_1287),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1335),
.A2(n_1326),
.B(n_1331),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1341),
.B(n_1333),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1340),
.Y(n_1347)
);

INVxp33_ASAP7_75t_SL g1348 ( 
.A(n_1342),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1339),
.A2(n_1269),
.B1(n_1324),
.B2(n_1328),
.Y(n_1349)
);

AOI21xp33_ASAP7_75t_L g1350 ( 
.A1(n_1339),
.A2(n_1272),
.B(n_1271),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1343),
.Y(n_1351)
);

AOI322xp5_ASAP7_75t_L g1352 ( 
.A1(n_1344),
.A2(n_1314),
.A3(n_1313),
.B1(n_1302),
.B2(n_1305),
.C1(n_1312),
.C2(n_1309),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1345),
.B(n_1279),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1347),
.B(n_1279),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1351),
.B(n_1302),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1353),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1355),
.A2(n_1352),
.B(n_1349),
.C(n_1346),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1356),
.Y(n_1359)
);

AOI22x1_ASAP7_75t_L g1360 ( 
.A1(n_1357),
.A2(n_1270),
.B1(n_1274),
.B2(n_1277),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1354),
.B(n_1273),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1360),
.Y(n_1362)
);

NAND4xp25_ASAP7_75t_L g1363 ( 
.A(n_1358),
.B(n_1283),
.C(n_1281),
.D(n_1277),
.Y(n_1363)
);

NAND4xp25_ASAP7_75t_L g1364 ( 
.A(n_1361),
.B(n_1283),
.C(n_1277),
.D(n_1273),
.Y(n_1364)
);

OAI211xp5_ASAP7_75t_L g1365 ( 
.A1(n_1359),
.A2(n_1282),
.B(n_1276),
.C(n_1278),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1363),
.B(n_184),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1362),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1364),
.B(n_185),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1365),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1367),
.B(n_1368),
.C(n_1366),
.Y(n_1370)
);

AOI211x1_ASAP7_75t_L g1371 ( 
.A1(n_1369),
.A2(n_187),
.B(n_191),
.C(n_192),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1371),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1370),
.B(n_207),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1372),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1373),
.Y(n_1375)
);

XOR2xp5_ASAP7_75t_L g1376 ( 
.A(n_1372),
.B(n_225),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1376),
.B(n_230),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1374),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1375),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1378),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1379),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1377),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1380),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1382),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1384),
.B(n_1381),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1383),
.B(n_263),
.C(n_268),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1385),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1386),
.A2(n_279),
.B1(n_288),
.B2(n_289),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1389)
);

AOI211xp5_ASAP7_75t_L g1390 ( 
.A1(n_1389),
.A2(n_295),
.B(n_298),
.C(n_300),
.Y(n_1390)
);


endmodule