module real_jpeg_8058_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_11, n_14, n_344, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_11;
input n_14;
input n_344;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_3),
.B(n_31),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_2),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_64),
.B1(n_67),
.B2(n_89),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_89),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_47),
.B(n_59),
.C(n_86),
.D(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_45),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_3),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_107),
.B(n_110),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_30),
.B(n_41),
.C(n_142),
.D(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_34),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_123),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_8),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_22),
.B1(n_64),
.B2(n_67),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_10),
.A2(n_22),
.B1(n_46),
.B2(n_47),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_33),
.B1(n_64),
.B2(n_67),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_54),
.B1(n_64),
.B2(n_67),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_54),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_64),
.B1(n_67),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_14),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_106),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_106),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_106),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_154),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_154),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_154),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_16),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_16),
.A2(n_64),
.B1(n_67),
.B2(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_101),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_16),
.A2(n_23),
.B1(n_24),
.B2(n_101),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_337),
.B(n_340),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_75),
.B(n_336),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_20),
.B(n_35),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_20),
.B(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_20),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_32),
.B2(n_34),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_21),
.A2(n_25),
.B1(n_34),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_23),
.A2(n_27),
.B(n_123),
.C(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_25),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_25),
.B(n_205),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_339)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_26),
.A2(n_29),
.B1(n_213),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_26),
.A2(n_204),
.B(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_286),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_29),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_29),
.A2(n_214),
.B(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_34),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_70),
.C(n_72),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_36),
.A2(n_37),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_57),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_38),
.A2(n_39),
.B1(n_57),
.B2(n_311),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_40),
.A2(n_49),
.B1(n_163),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_40),
.A2(n_199),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_45),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_41),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_41),
.A2(n_45),
.B1(n_239),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_41),
.A2(n_45),
.B1(n_258),
.B2(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_42),
.B(n_47),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_44),
.A2(n_46),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_49),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_49),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_49),
.A2(n_164),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_51),
.A2(n_52),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_57),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_57),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_58),
.A2(n_68),
.B1(n_100),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_58),
.A2(n_140),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_58),
.A2(n_68),
.B1(n_196),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_58),
.A2(n_68),
.B1(n_224),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_58),
.A2(n_68),
.B1(n_233),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_59),
.A2(n_63),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_67),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_64),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_67),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_68),
.A2(n_102),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_70),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_329),
.B(n_335),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_302),
.A3(n_322),
.B1(n_327),
.B2(n_328),
.C(n_344),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_250),
.A3(n_290),
.B1(n_296),
.B2(n_301),
.C(n_345),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_207),
.C(n_246),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_178),
.B(n_206),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_157),
.B(n_177),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_134),
.B(n_156),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_112),
.B(n_133),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_84),
.B(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_87),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_99),
.C(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_107),
.A2(n_125),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_107),
.A2(n_125),
.B1(n_189),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_107),
.A2(n_125),
.B1(n_222),
.B2(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_107),
.A2(n_125),
.B(n_231),
.Y(n_263)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_108),
.A2(n_109),
.B1(n_153),
.B2(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B(n_132),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_118),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_127),
.B(n_131),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_126),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_147),
.B2(n_155),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_146),
.C(n_155),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_143),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_147),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_171),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_173),
.C(n_175),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_170),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_167),
.C(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_180),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_182),
.B(n_192),
.C(n_193),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_187),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_208),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_226),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_209),
.B(n_226),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.C(n_225),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_225),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_223),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_244),
.B2(n_245),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_234),
.C(n_245),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_232),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_240),
.C(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_248),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_268),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_251),
.B(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_261),
.C(n_267),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_252),
.A2(n_253),
.B1(n_261),
.B2(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_261),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_263),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_281),
.B(n_285),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_288),
.B2(n_289),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_279),
.B2(n_280),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_280),
.C(n_289),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_278),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_276),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_304),
.B1(n_313),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_287),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_283),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.C(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_317),
.C(n_321),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_339),
.B(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);


endmodule