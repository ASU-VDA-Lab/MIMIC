module fake_ariane_641_n_2004 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2004);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2004;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_274;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_97),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

CKINVDCx11_ASAP7_75t_R g205 ( 
.A(n_4),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_84),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_77),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_196),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_144),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_72),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_30),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_20),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_149),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_29),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_8),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_9),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_13),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_14),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_61),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_161),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_52),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_16),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_51),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_174),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_49),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_74),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_156),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_66),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_95),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_67),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_53),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_119),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_152),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_19),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_107),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_70),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_92),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_39),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_96),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_75),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_135),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_98),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_64),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_121),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_37),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_88),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_106),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_182),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_6),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_79),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_71),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_100),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_41),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_115),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_172),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_93),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_142),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_164),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_35),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_101),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_55),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_76),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_192),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_94),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_5),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_55),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_7),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_127),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_134),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_25),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_30),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_110),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_68),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_180),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_36),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_11),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_86),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_2),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_45),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_78),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_81),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_89),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_22),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_82),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_102),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_1),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_122),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_21),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_38),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_150),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_50),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_7),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_137),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_40),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_116),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_56),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_14),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_15),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_22),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_42),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_28),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_64),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_91),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_40),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_53),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_125),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_108),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_57),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_154),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_188),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_175),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_56),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_28),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_62),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_85),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_145),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_0),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_9),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_157),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_68),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_39),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_52),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_27),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_118),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_132),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

BUFx10_ASAP7_75t_L g370 ( 
.A(n_126),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_29),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_46),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_104),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_136),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_195),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_167),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_160),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_185),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_44),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_1),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_103),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_173),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_186),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_0),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_57),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_49),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_65),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_32),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_123),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_67),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_37),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_70),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_163),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_105),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_2),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_45),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_158),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_257),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_312),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_205),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_257),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_278),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_203),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_312),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_312),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_296),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_363),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_283),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_223),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_224),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_307),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_322),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_335),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_335),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_342),
.Y(n_438)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_243),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_246),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_342),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_233),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_215),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_289),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_233),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_219),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_342),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_233),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_323),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_225),
.Y(n_452)
);

BUFx2_ASAP7_75t_SL g453 ( 
.A(n_370),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_236),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_220),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_370),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_320),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_264),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_265),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_370),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_269),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_217),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_272),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_275),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_344),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_297),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_330),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_302),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_309),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_383),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_316),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_324),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_327),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_383),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_333),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_372),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_341),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_213),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_343),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_199),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_359),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_360),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_213),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_380),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_199),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_201),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_201),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_204),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_344),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_217),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_344),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_344),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_216),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_216),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_221),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_254),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_396),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_236),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_254),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_311),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_454),
.B(n_281),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_403),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_436),
.B(n_290),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_262),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_281),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_262),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_432),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_457),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_431),
.B(n_328),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_415),
.A2(n_229),
.B(n_214),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_469),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_467),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_467),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_479),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_399),
.B(n_273),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_419),
.A2(n_229),
.B(n_214),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_503),
.B(n_317),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_406),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_431),
.A2(n_354),
.B1(n_387),
.B2(n_319),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_502),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_407),
.B(n_273),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_410),
.B(n_315),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_419),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_453),
.B(n_456),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_408),
.A2(n_222),
.B1(n_227),
.B2(n_221),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_453),
.B(n_315),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_423),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_424),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_425),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_456),
.B(n_366),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_427),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_434),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_445),
.B(n_366),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_497),
.B(n_311),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_429),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_429),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_497),
.B(n_386),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_433),
.B(n_325),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_435),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

NOR2x1_ASAP7_75t_L g579 ( 
.A(n_438),
.B(n_252),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_451),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_483),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_208),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_452),
.B(n_208),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_499),
.B(n_204),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_442),
.B(n_197),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_498),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_442),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_512),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_559),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_512),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_574),
.Y(n_596)
);

AOI21x1_ASAP7_75t_L g597 ( 
.A1(n_506),
.A2(n_495),
.B(n_492),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_555),
.B(n_458),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_513),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_557),
.B(n_563),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_543),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_546),
.A2(n_440),
.B1(n_439),
.B2(n_405),
.Y(n_604)
);

AND3x2_ASAP7_75t_L g605 ( 
.A(n_515),
.B(n_440),
.C(n_486),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_513),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_557),
.B(n_455),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_543),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_521),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_443),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_563),
.B(n_443),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_563),
.B(n_520),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_555),
.B(n_409),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_554),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_555),
.B(n_483),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_586),
.B(n_447),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_533),
.B(n_508),
.C(n_506),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_586),
.B(n_447),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_450),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_560),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_560),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_546),
.B(n_421),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_509),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_546),
.B(n_421),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_521),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_546),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_580),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_524),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_510),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_509),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

AND3x2_ASAP7_75t_L g640 ( 
.A(n_515),
.B(n_500),
.C(n_292),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_569),
.Y(n_641)
);

AND2x2_ASAP7_75t_SL g642 ( 
.A(n_533),
.B(n_317),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_584),
.B(n_585),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_510),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_579),
.B(n_325),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_559),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_517),
.B(n_488),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_576),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_564),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_521),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_517),
.B(n_489),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_521),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_521),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_561),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_561),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_508),
.B(n_490),
.C(n_489),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_584),
.A2(n_481),
.B1(n_505),
.B2(n_450),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_570),
.B(n_490),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_520),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_426),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_576),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_576),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_576),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_577),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_566),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_576),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_517),
.B(n_491),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_590),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_561),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_517),
.B(n_491),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_519),
.B(n_426),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_561),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_547),
.B(n_461),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_590),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_561),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_584),
.A2(n_461),
.B1(n_473),
.B2(n_465),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_528),
.B(n_465),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_523),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_584),
.B(n_473),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_528),
.B(n_477),
.Y(n_693)
);

BUFx10_ASAP7_75t_L g694 ( 
.A(n_528),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_428),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_523),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_559),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_577),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_591),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_581),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_523),
.Y(n_702)
);

AO21x2_ASAP7_75t_L g703 ( 
.A1(n_534),
.A2(n_545),
.B(n_514),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_591),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_528),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_511),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_511),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_514),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_584),
.B(n_477),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_518),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_518),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_539),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_522),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_589),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_568),
.B(n_463),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_539),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_585),
.B(n_412),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_510),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_585),
.B(n_417),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_525),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_568),
.B(n_494),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_559),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_539),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_539),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_581),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_585),
.B(n_206),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_526),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_559),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_552),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_559),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_526),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_527),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_585),
.B(n_206),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_510),
.B(n_460),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_547),
.B(n_211),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_547),
.B(n_211),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_532),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_548),
.A2(n_227),
.B1(n_232),
.B2(n_222),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_559),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_668),
.B(n_548),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_617),
.B(n_589),
.Y(n_744)
);

O2A1O1Ixp5_ASAP7_75t_L g745 ( 
.A1(n_652),
.A2(n_657),
.B(n_659),
.C(n_656),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_698),
.B(n_552),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_642),
.B(n_552),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_598),
.B(n_529),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_633),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_633),
.B(n_529),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_641),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_614),
.B(n_529),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_642),
.A2(n_556),
.B1(n_579),
.B2(n_529),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_611),
.B(n_556),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_529),
.Y(n_755)
);

NOR3xp33_ASAP7_75t_L g756 ( 
.A(n_665),
.B(n_303),
.C(n_232),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_669),
.B(n_552),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_655),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_642),
.B(n_552),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_598),
.A2(n_535),
.B1(n_541),
.B2(n_527),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_681),
.B(n_553),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_698),
.B(n_721),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_655),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_648),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_613),
.B(n_532),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_683),
.B(n_553),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_698),
.B(n_553),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_623),
.A2(n_541),
.B(n_535),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_628),
.B(n_536),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_666),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_666),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_630),
.B(n_536),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_598),
.A2(n_355),
.B1(n_356),
.B2(n_303),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_670),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_595),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_595),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_698),
.B(n_553),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_667),
.B(n_553),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_698),
.B(n_558),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_670),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_595),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_598),
.A2(n_567),
.B1(n_568),
.B2(n_544),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_651),
.B(n_675),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_598),
.B(n_562),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_619),
.B(n_542),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_644),
.B(n_562),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_698),
.B(n_565),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_621),
.B(n_565),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_721),
.B(n_328),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_624),
.B(n_542),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_625),
.B(n_550),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_706),
.A2(n_545),
.B(n_534),
.C(n_572),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_678),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_678),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_626),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_661),
.B(n_549),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_626),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_741),
.A2(n_567),
.B1(n_544),
.B2(n_572),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_737),
.B(n_550),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_721),
.B(n_507),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_661),
.B(n_549),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_607),
.B(n_550),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_637),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_715),
.B(n_567),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_684),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_715),
.A2(n_722),
.B1(n_692),
.B2(n_648),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_699),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_684),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_700),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_706),
.B(n_551),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_722),
.A2(n_398),
.B1(n_210),
.B2(n_255),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_700),
.Y(n_817)
);

OAI21xp33_ASAP7_75t_L g818 ( 
.A1(n_688),
.A2(n_356),
.B(n_355),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_704),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_648),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_721),
.B(n_507),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_635),
.B(n_551),
.Y(n_822)
);

NOR2x1p5_ASAP7_75t_L g823 ( 
.A(n_701),
.B(n_404),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_707),
.B(n_551),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_707),
.B(n_567),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_721),
.B(n_507),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_635),
.B(n_572),
.Y(n_827)
);

BUFx8_ASAP7_75t_SL g828 ( 
.A(n_674),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_362),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_593),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_721),
.B(n_507),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_708),
.B(n_567),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_708),
.B(n_544),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_599),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_710),
.B(n_544),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_710),
.B(n_544),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_711),
.B(n_713),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_653),
.B(n_462),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_623),
.A2(n_365),
.B1(n_371),
.B2(n_362),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_592),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_713),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_723),
.B(n_507),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_723),
.B(n_742),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_645),
.B(n_592),
.Y(n_844)
);

INVx3_ASAP7_75t_R g845 ( 
.A(n_714),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_648),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_L g847 ( 
.A(n_723),
.B(n_328),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_599),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_720),
.B(n_592),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_723),
.B(n_507),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_723),
.B(n_507),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_720),
.B(n_592),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_600),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_600),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_729),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_696),
.B(n_464),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_606),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_729),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_606),
.Y(n_859)
);

BUFx8_ASAP7_75t_L g860 ( 
.A(n_714),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_730),
.B(n_531),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_616),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_365),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_730),
.B(n_531),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_727),
.A2(n_740),
.B1(n_664),
.B2(n_604),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_734),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_668),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_734),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_735),
.A2(n_388),
.B1(n_392),
.B2(n_371),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_645),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_662),
.B(n_466),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_735),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_636),
.B(n_531),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_636),
.B(n_531),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_638),
.B(n_531),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_615),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_723),
.B(n_328),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_616),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_742),
.B(n_507),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_638),
.B(n_537),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_602),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_602),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_603),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_689),
.B(n_691),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_SL g885 ( 
.A(n_693),
.B(n_393),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_615),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_603),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_741),
.A2(n_537),
.B1(n_588),
.B2(n_575),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_SL g889 ( 
.A(n_649),
.B(n_393),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_742),
.B(n_328),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_689),
.B(n_537),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_654),
.B(n_677),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_680),
.B(n_235),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_691),
.B(n_537),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_634),
.B(n_468),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_696),
.B(n_238),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_695),
.B(n_537),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_687),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_615),
.B(n_470),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_615),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_605),
.B(n_472),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_742),
.B(n_534),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_754),
.A2(n_646),
.B1(n_608),
.B2(n_612),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_867),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_748),
.B(n_717),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_827),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_828),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_766),
.A2(n_687),
.B1(n_705),
.B2(n_694),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_807),
.B(n_687),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_876),
.B(n_742),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_758),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_794),
.A2(n_694),
.B1(n_705),
.B2(n_719),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_777),
.Y(n_914)
);

AND2x6_ASAP7_75t_SL g915 ( 
.A(n_744),
.B(n_474),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_749),
.B(n_694),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_838),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_811),
.B(n_728),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_748),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_795),
.B(n_694),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_763),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_764),
.B(n_643),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_764),
.B(n_643),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_856),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_796),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_748),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_902),
.A2(n_697),
.B(n_695),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_791),
.B(n_705),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_765),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_778),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_778),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_828),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_771),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_860),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_820),
.B(n_643),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_796),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_784),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_784),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_796),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_809),
.B(n_645),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_752),
.B(n_705),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_796),
.B(n_718),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_755),
.B(n_757),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_809),
.B(n_718),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_761),
.B(n_718),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_892),
.A2(n_736),
.B1(n_739),
.B2(n_738),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_753),
.B(n_610),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_899),
.B(n_610),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_772),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_856),
.B(n_612),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_809),
.B(n_640),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_856),
.A2(n_646),
.B1(n_618),
.B2(n_627),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_770),
.A2(n_242),
.B1(n_245),
.B2(n_241),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_886),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_820),
.B(n_643),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_846),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_793),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_822),
.B(n_697),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_776),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_815),
.A2(n_618),
.B(n_627),
.C(n_620),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_783),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_786),
.B(n_629),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_846),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_871),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_774),
.A2(n_646),
.B1(n_620),
.B2(n_650),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_782),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_896),
.A2(n_646),
.B1(n_671),
.B2(n_650),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_783),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_750),
.B(n_702),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_804),
.B(n_702),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_793),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_886),
.Y(n_973)
);

INVxp33_ASAP7_75t_L g974 ( 
.A(n_812),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_860),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_800),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_760),
.A2(n_716),
.B1(n_724),
.B2(n_712),
.Y(n_977)
);

AO22x2_ASAP7_75t_L g978 ( 
.A1(n_743),
.A2(n_501),
.B1(n_504),
.B2(n_499),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_798),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_860),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_785),
.B(n_716),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_823),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_799),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_895),
.B(n_475),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_901),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_801),
.B(n_724),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_787),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_824),
.B(n_725),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_876),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_900),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_726),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_900),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_898),
.B(n_643),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_788),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_865),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_783),
.B(n_643),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_808),
.B(n_679),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_806),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_810),
.B(n_732),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_808),
.B(n_679),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_813),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_845),
.A2(n_816),
.B1(n_829),
.B2(n_863),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_818),
.A2(n_251),
.B(n_248),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_800),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_814),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

NOR2x2_ASAP7_75t_L g1007 ( 
.A(n_775),
.B(n_671),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_819),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_893),
.A2(n_646),
.B1(n_673),
.B2(n_672),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_808),
.B(n_679),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_802),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_780),
.B(n_767),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_802),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_870),
.B(n_679),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_870),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_889),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_803),
.A2(n_480),
.B1(n_476),
.B2(n_487),
.C(n_478),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_889),
.A2(n_646),
.B1(n_673),
.B2(n_672),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_870),
.B(n_679),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_844),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_837),
.B(n_679),
.Y(n_1022)
);

INVx5_ASAP7_75t_L g1023 ( 
.A(n_881),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_855),
.B(n_858),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_866),
.B(n_732),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_868),
.Y(n_1026)
);

AO22x1_ASAP7_75t_L g1027 ( 
.A1(n_756),
.A2(n_839),
.B1(n_869),
.B2(n_872),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_789),
.B(n_629),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_882),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_830),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_830),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_888),
.B(n_482),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_R g1033 ( 
.A(n_885),
.B(n_746),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_882),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_825),
.B(n_632),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_832),
.B(n_484),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_745),
.A2(n_656),
.B(n_652),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_833),
.B(n_639),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_835),
.B(n_639),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_836),
.B(n_646),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_747),
.B(n_594),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_746),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_747),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_883),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_887),
.B(n_676),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_759),
.B(n_596),
.Y(n_1046)
);

BUFx8_ASAP7_75t_L g1047 ( 
.A(n_834),
.Y(n_1047)
);

BUFx12f_ASAP7_75t_L g1048 ( 
.A(n_885),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_873),
.Y(n_1049)
);

NOR2x1p5_ASAP7_75t_L g1050 ( 
.A(n_861),
.B(n_485),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_759),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_779),
.B(n_276),
.C(n_253),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_834),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_805),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_848),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_768),
.B(n_884),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_805),
.B(n_501),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_821),
.B(n_504),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_848),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_821),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_769),
.B(n_742),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_853),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_874),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_853),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_864),
.B(n_685),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_854),
.B(n_609),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_857),
.B(n_285),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_762),
.B(n_594),
.Y(n_1068)
);

BUFx2_ASAP7_75t_R g1069 ( 
.A(n_826),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_857),
.B(n_609),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_762),
.B(n_594),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_859),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_826),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_990),
.B(n_792),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_994),
.B(n_875),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_1047),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1042),
.A2(n_943),
.B(n_1012),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_908),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_SL g1079 ( 
.A(n_913),
.B(n_294),
.C(n_287),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_928),
.A2(n_840),
.B1(n_852),
.B2(n_849),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1042),
.A2(n_880),
.B1(n_894),
.B2(n_891),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_903),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_917),
.B(n_859),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_905),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_920),
.A2(n_897),
.B1(n_768),
.B2(n_790),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_917),
.B(n_862),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_998),
.B(n_831),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1002),
.B(n_831),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_926),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1043),
.A2(n_797),
.B(n_790),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_926),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_965),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_924),
.A2(n_843),
.B1(n_850),
.B2(n_842),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1012),
.A2(n_902),
.B(n_843),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_910),
.A2(n_781),
.B1(n_609),
.B2(n_631),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1061),
.A2(n_781),
.B(n_797),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_987),
.B(n_862),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_965),
.B(n_878),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_1005),
.A2(n_305),
.B(n_295),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_922),
.A2(n_923),
.B(n_956),
.C(n_935),
.Y(n_1100)
);

NOR2x1_ASAP7_75t_L g1101 ( 
.A(n_980),
.B(n_842),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_984),
.B(n_306),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_934),
.B(n_850),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_924),
.B(n_851),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_975),
.B(n_851),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_907),
.B(n_310),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_915),
.B(n_879),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1032),
.A2(n_588),
.B1(n_575),
.B2(n_573),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_907),
.B(n_879),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_941),
.A2(n_622),
.B1(n_631),
.B2(n_682),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1036),
.B(n_622),
.Y(n_1111)
);

AO32x2_ASAP7_75t_L g1112 ( 
.A1(n_977),
.A2(n_647),
.A3(n_594),
.B1(n_703),
.B2(n_792),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_957),
.B(n_622),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1047),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1061),
.A2(n_877),
.B(n_847),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_995),
.B(n_954),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_952),
.B(n_313),
.Y(n_1117)
);

NOR2xp67_ASAP7_75t_R g1118 ( 
.A(n_989),
.B(n_647),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_631),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_974),
.B(n_647),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_959),
.B(n_682),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_992),
.B(n_647),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_912),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_909),
.B(n_682),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_961),
.A2(n_890),
.B(n_877),
.C(n_847),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_921),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_919),
.B(n_731),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_906),
.B(n_731),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_929),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_906),
.B(n_731),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_927),
.A2(n_1037),
.B(n_1022),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_986),
.B(n_731),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_1051),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_986),
.B(n_733),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_945),
.A2(n_890),
.B(n_659),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_951),
.B(n_733),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1030),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_927),
.A2(n_545),
.B(n_657),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_961),
.A2(n_575),
.B(n_573),
.C(n_663),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_963),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_963),
.B(n_659),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_906),
.B(n_733),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1031),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_952),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_963),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_918),
.A2(n_573),
.B(n_663),
.C(n_660),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_939),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_932),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_916),
.A2(n_663),
.B(n_660),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_955),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_946),
.A2(n_660),
.B(n_686),
.C(n_685),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1059),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_948),
.B(n_733),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_940),
.B(n_686),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_978),
.B(n_332),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1018),
.A2(n_347),
.B1(n_350),
.B2(n_346),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_978),
.B(n_1067),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_922),
.A2(n_337),
.B(n_202),
.C(n_207),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_978),
.B(n_338),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1028),
.A2(n_703),
.B(n_209),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_940),
.B(n_212),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_971),
.A2(n_997),
.B(n_996),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1024),
.A2(n_397),
.B(n_340),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_985),
.B(n_703),
.Y(n_1164)
);

AOI21x1_ASAP7_75t_L g1165 ( 
.A1(n_923),
.A2(n_956),
.B(n_935),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_996),
.A2(n_226),
.B(n_200),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_997),
.A2(n_597),
.B(n_530),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1064),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1000),
.A2(n_1015),
.B(n_1010),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1003),
.A2(n_260),
.B(n_299),
.C(n_298),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_944),
.B(n_212),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1000),
.A2(n_230),
.B(n_228),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_944),
.B(n_218),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_904),
.A2(n_382),
.B1(n_353),
.B2(n_218),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_973),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_904),
.A2(n_384),
.B1(n_361),
.B2(n_368),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_939),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1010),
.A2(n_258),
.B(n_231),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_933),
.A2(n_368),
.B1(n_369),
.B2(n_373),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_982),
.Y(n_1180)
);

INVxp33_ASAP7_75t_SL g1181 ( 
.A(n_1033),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_949),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1029),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_925),
.B(n_277),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_1048),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_911),
.B(n_925),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1017),
.B(n_349),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1069),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1051),
.B(n_374),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_950),
.B(n_300),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_960),
.A2(n_395),
.B1(n_300),
.B2(n_301),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1021),
.B(n_516),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1034),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_967),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1018),
.B(n_379),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1021),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1023),
.B(n_301),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1050),
.A2(n_369),
.B1(n_373),
.B2(n_375),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_SL g1199 ( 
.A(n_1057),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1069),
.B(n_353),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1015),
.A2(n_304),
.B(n_282),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1027),
.A2(n_377),
.B1(n_382),
.B2(n_361),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_939),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1023),
.B(n_375),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_979),
.A2(n_378),
.B1(n_395),
.B2(n_384),
.Y(n_1205)
);

OAI22x1_ASAP7_75t_L g1206 ( 
.A1(n_983),
.A2(n_1006),
.B1(n_1008),
.B2(n_1001),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1033),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1014),
.B(n_377),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1026),
.B(n_378),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_939),
.Y(n_1210)
);

BUFx4f_ASAP7_75t_L g1211 ( 
.A(n_1021),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1044),
.B(n_516),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1053),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1054),
.B(n_198),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1020),
.A2(n_357),
.B(n_367),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1060),
.B(n_234),
.Y(n_1216)
);

AO22x1_ASAP7_75t_L g1217 ( 
.A1(n_1023),
.A2(n_331),
.B1(n_376),
.B2(n_390),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_988),
.A2(n_394),
.B(n_495),
.C(n_492),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1007),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1062),
.B(n_516),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1055),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1082),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1160),
.A2(n_993),
.B(n_1020),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_1039),
.B(n_1068),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1131),
.A2(n_1071),
.B(n_1068),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1088),
.A2(n_966),
.B(n_1025),
.C(n_1041),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1102),
.B(n_1057),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1213),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1077),
.A2(n_1056),
.B(n_1041),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1096),
.A2(n_1071),
.B(n_1045),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1115),
.A2(n_1070),
.B(n_1066),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1115),
.A2(n_942),
.B(n_999),
.Y(n_1232)
);

AOI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1094),
.A2(n_1049),
.B1(n_1063),
.B2(n_1016),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1097),
.B(n_947),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1181),
.A2(n_1025),
.B(n_1056),
.C(n_1052),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1116),
.B(n_1058),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1113),
.A2(n_1040),
.B(n_970),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1156),
.A2(n_981),
.B1(n_968),
.B2(n_953),
.Y(n_1238)
);

CKINVDCx9p33_ASAP7_75t_R g1239 ( 
.A(n_1122),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1081),
.A2(n_1065),
.B(n_964),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1150),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1080),
.A2(n_1065),
.B(n_964),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1078),
.Y(n_1243)
);

NOR2x1_ASAP7_75t_SL g1244 ( 
.A(n_1192),
.B(n_957),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1160),
.A2(n_1125),
.B(n_1135),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1202),
.A2(n_1023),
.B1(n_1009),
.B2(n_1019),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1092),
.B(n_1058),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1135),
.A2(n_930),
.B(n_914),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1167),
.A2(n_937),
.B(n_931),
.Y(n_1249)
);

INVx8_ASAP7_75t_L g1250 ( 
.A(n_1175),
.Y(n_1250)
);

AOI221xp5_ASAP7_75t_L g1251 ( 
.A1(n_1156),
.A2(n_1038),
.B1(n_1035),
.B2(n_953),
.C(n_1073),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1075),
.B(n_969),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1125),
.A2(n_964),
.B(n_957),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1221),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1132),
.A2(n_957),
.B(n_969),
.Y(n_1255)
);

BUFx4f_ASAP7_75t_L g1256 ( 
.A(n_1076),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1221),
.B(n_1016),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1134),
.A2(n_962),
.B(n_991),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1162),
.A2(n_938),
.A3(n_972),
.B(n_976),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1162),
.A2(n_962),
.B(n_991),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1098),
.B(n_1035),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1123),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1126),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1129),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1100),
.A2(n_962),
.B(n_1038),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1144),
.B(n_1072),
.Y(n_1266)
);

NAND3x1_ASAP7_75t_L g1267 ( 
.A(n_1200),
.B(n_496),
.C(n_4),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1183),
.B(n_958),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1153),
.A2(n_962),
.B(n_936),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1155),
.B(n_1106),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1169),
.A2(n_1004),
.B(n_1011),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1193),
.B(n_1013),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1207),
.A2(n_1021),
.B1(n_1046),
.B2(n_540),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1182),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1133),
.B(n_1046),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1219),
.B(n_530),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1169),
.A2(n_538),
.B(n_540),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1149),
.A2(n_538),
.B(n_540),
.Y(n_1279)
);

NOR2x1_ASAP7_75t_R g1280 ( 
.A(n_1114),
.B(n_237),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1211),
.B(n_538),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_328),
.A3(n_578),
.B(n_571),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1149),
.A2(n_325),
.B(n_358),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1157),
.B(n_571),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1188),
.B(n_571),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1206),
.A2(n_328),
.A3(n_578),
.B(n_571),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1117),
.B(n_3),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1165),
.A2(n_578),
.B(n_571),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1211),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1180),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1084),
.B(n_11),
.Y(n_1291)
);

OAI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1163),
.A2(n_263),
.B(n_261),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1194),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1199),
.B(n_325),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1148),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1089),
.B(n_239),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1090),
.A2(n_574),
.B(n_240),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1146),
.A2(n_574),
.B(n_244),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1136),
.A2(n_325),
.B(n_358),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1085),
.A2(n_351),
.B(n_358),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1185),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1079),
.A2(n_12),
.B(n_13),
.Y(n_1302)
);

AO22x2_ASAP7_75t_L g1303 ( 
.A1(n_1159),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1138),
.A2(n_578),
.B(n_328),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1138),
.A2(n_578),
.B(n_153),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1107),
.B(n_247),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1101),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1124),
.A2(n_1111),
.B(n_1204),
.C(n_1197),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1209),
.B(n_17),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_SL g1310 ( 
.A(n_1089),
.B(n_596),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1170),
.A2(n_574),
.A3(n_358),
.B(n_351),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1109),
.B(n_23),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1137),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1146),
.A2(n_351),
.B(n_358),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1139),
.A2(n_151),
.B(n_90),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1190),
.B(n_23),
.Y(n_1317)
);

NAND3x1_ASAP7_75t_L g1318 ( 
.A(n_1187),
.B(n_1087),
.C(n_1189),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1166),
.A2(n_1178),
.B(n_1172),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1198),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1189),
.B(n_24),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1143),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1141),
.B(n_1179),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1074),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1152),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1141),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1191),
.B(n_26),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1110),
.A2(n_178),
.B(n_80),
.Y(n_1328)
);

OAI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1161),
.A2(n_336),
.B1(n_266),
.B2(n_259),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1095),
.A2(n_351),
.B(n_352),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1168),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1128),
.B(n_27),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1205),
.B(n_31),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1220),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1196),
.B(n_73),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1118),
.A2(n_286),
.B(n_348),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1166),
.A2(n_574),
.A3(n_596),
.B(n_147),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1130),
.B(n_31),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1103),
.B(n_596),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1142),
.B(n_32),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1091),
.B(n_284),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1121),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1079),
.A2(n_280),
.B(n_345),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1199),
.A2(n_288),
.B1(n_250),
.B2(n_334),
.Y(n_1345)
);

BUFx8_ASAP7_75t_L g1346 ( 
.A(n_1177),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1164),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1091),
.B(n_279),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1201),
.A2(n_574),
.A3(n_596),
.B(n_130),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1215),
.A2(n_291),
.B(n_256),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1147),
.A2(n_114),
.B(n_109),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1112),
.A2(n_574),
.A3(n_596),
.B(n_138),
.Y(n_1352)
);

OAI22x1_ASAP7_75t_L g1353 ( 
.A1(n_1171),
.A2(n_270),
.B1(n_268),
.B2(n_267),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1093),
.A2(n_574),
.B(n_326),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1127),
.A2(n_321),
.B(n_314),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1104),
.B(n_33),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1212),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1203),
.A2(n_1184),
.B(n_1218),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1119),
.A2(n_308),
.B(n_293),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1119),
.A2(n_274),
.B(n_271),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1218),
.A2(n_34),
.B(n_35),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1112),
.A2(n_574),
.A3(n_187),
.B(n_194),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1208),
.A2(n_34),
.B1(n_36),
.B2(n_42),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1196),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1173),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1365)
);

NOR4xp25_ASAP7_75t_L g1366 ( 
.A(n_1174),
.B(n_43),
.C(n_47),
.D(n_50),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1154),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1176),
.A2(n_249),
.B(n_58),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1196),
.B(n_47),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1259),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1366),
.A2(n_1368),
.B1(n_1303),
.B2(n_1302),
.C(n_1320),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1347),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1346),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1302),
.A2(n_1216),
.B(n_1214),
.C(n_1099),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1222),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1254),
.B(n_1120),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1259),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1304),
.A2(n_1283),
.B(n_1305),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1346),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1241),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1229),
.A2(n_1108),
.B(n_1112),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1229),
.A2(n_1224),
.B(n_1230),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1226),
.A2(n_1158),
.B(n_1105),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1288),
.A2(n_1112),
.B(n_1186),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1228),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1300),
.A2(n_1242),
.B(n_1240),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1225),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1233),
.A2(n_1192),
.B(n_1210),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1231),
.A2(n_1232),
.B(n_1223),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1343),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1315),
.A2(n_1299),
.B(n_1298),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1248),
.A2(n_1210),
.B(n_1177),
.Y(n_1392)
);

AO32x2_ASAP7_75t_L g1393 ( 
.A1(n_1363),
.A2(n_1217),
.A3(n_1177),
.B1(n_60),
.B2(n_61),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_SL g1394 ( 
.A(n_1366),
.B(n_1321),
.C(n_1313),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1364),
.B(n_193),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1246),
.B(n_58),
.Y(n_1396)
);

AOI22x1_ASAP7_75t_L g1397 ( 
.A1(n_1329),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1321),
.B(n_63),
.Y(n_1398)
);

AOI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1253),
.A2(n_113),
.B(n_184),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1270),
.B(n_69),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1249),
.A2(n_69),
.B(n_1271),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1324),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1262),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1318),
.A2(n_1313),
.B(n_1297),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1320),
.A2(n_1363),
.B(n_1368),
.C(n_1356),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1256),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1298),
.A2(n_1237),
.B(n_1297),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_SL g1408 ( 
.A1(n_1252),
.A2(n_1333),
.B(n_1339),
.C(n_1341),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1227),
.B(n_1247),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1303),
.A2(n_1236),
.B1(n_1309),
.B2(n_1238),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1238),
.A2(n_1327),
.B1(n_1334),
.B2(n_1317),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1252),
.A2(n_1333),
.B1(n_1341),
.B2(n_1339),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1263),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1264),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1306),
.A2(n_1260),
.B(n_1354),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1279),
.A2(n_1278),
.B(n_1316),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1255),
.A2(n_1269),
.B(n_1258),
.Y(n_1417)
);

AOI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1292),
.A2(n_1350),
.B(n_1234),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1354),
.A2(n_1344),
.B(n_1330),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1287),
.B(n_1277),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1282),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1235),
.A2(n_1308),
.B(n_1328),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1364),
.B(n_1331),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1275),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1284),
.A2(n_1319),
.B(n_1358),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_L g1427 ( 
.A(n_1243),
.B(n_1295),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1294),
.A2(n_1261),
.B1(n_1312),
.B2(n_1257),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1351),
.A2(n_1284),
.B(n_1276),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1293),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1257),
.A2(n_1256),
.B1(n_1228),
.B2(n_1323),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_SL g1432 ( 
.A(n_1294),
.B(n_1301),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1365),
.A2(n_1361),
.B(n_1369),
.C(n_1291),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1243),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1335),
.B(n_1312),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1272),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1289),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1314),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1250),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1325),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1268),
.A2(n_1273),
.B(n_1357),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1332),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1326),
.B(n_1244),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1266),
.B(n_1285),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1345),
.A2(n_1267),
.B1(n_1251),
.B2(n_1348),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1353),
.A2(n_1355),
.B1(n_1296),
.B2(n_1342),
.C(n_1272),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1307),
.B(n_1250),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1336),
.A2(n_1367),
.B(n_1310),
.C(n_1337),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1290),
.A2(n_1350),
.B1(n_1239),
.B2(n_1241),
.Y(n_1449)
);

BUFx8_ASAP7_75t_SL g1450 ( 
.A(n_1280),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1340),
.A2(n_1360),
.B1(n_1359),
.B2(n_1281),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1322),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1340),
.B(n_1362),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1282),
.A2(n_1286),
.B(n_1352),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1340),
.A2(n_1362),
.B1(n_1352),
.B2(n_1338),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1362),
.A2(n_1352),
.B1(n_1338),
.B2(n_1349),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1286),
.B(n_1338),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1282),
.A2(n_1349),
.B(n_1311),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1349),
.A2(n_1304),
.B(n_1283),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1311),
.A2(n_754),
.B1(n_1366),
.B2(n_741),
.C(n_556),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1311),
.A2(n_1304),
.B(n_1283),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1326),
.B(n_1364),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1304),
.A2(n_1283),
.B(n_1305),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1283),
.B(n_1305),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1226),
.B(n_1077),
.Y(n_1466)
);

AOI21xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1250),
.A2(n_675),
.B(n_651),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1302),
.A2(n_744),
.B(n_754),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_770),
.B1(n_774),
.B2(n_1002),
.Y(n_1469)
);

INVx6_ASAP7_75t_L g1470 ( 
.A(n_1346),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1229),
.A2(n_1077),
.B(n_1113),
.Y(n_1471)
);

AO32x2_ASAP7_75t_L g1472 ( 
.A1(n_1363),
.A2(n_1320),
.A3(n_1238),
.B1(n_1274),
.B2(n_865),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1222),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1222),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1222),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1245),
.A2(n_1160),
.B(n_1315),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1254),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1226),
.A2(n_754),
.B(n_1077),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1245),
.A2(n_1304),
.B(n_1229),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1222),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1226),
.A2(n_754),
.B(n_1077),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1254),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1222),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1274),
.B(n_1258),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1366),
.A2(n_754),
.B1(n_741),
.B2(n_556),
.C(n_744),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1274),
.B(n_1258),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

AO21x1_ASAP7_75t_L g1489 ( 
.A1(n_1302),
.A2(n_1321),
.B(n_1313),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1245),
.A2(n_1160),
.B(n_1315),
.Y(n_1490)
);

AOI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1283),
.A2(n_1300),
.B(n_1245),
.Y(n_1491)
);

AOI222xp33_ASAP7_75t_L g1492 ( 
.A1(n_1309),
.A2(n_865),
.B1(n_754),
.B2(n_1195),
.C1(n_1002),
.C2(n_556),
.Y(n_1492)
);

XOR2xp5_ASAP7_75t_L g1493 ( 
.A(n_1324),
.B(n_674),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1245),
.A2(n_1283),
.B(n_1305),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1347),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1274),
.B(n_1258),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1347),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1259),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1347),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1254),
.B(n_1347),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1326),
.B(n_1364),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1346),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1245),
.A2(n_1283),
.B(n_1305),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1245),
.A2(n_1283),
.B(n_1305),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1313),
.A2(n_1202),
.B1(n_754),
.B2(n_1156),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1226),
.A2(n_754),
.B(n_1077),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1222),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1245),
.A2(n_1283),
.B(n_1305),
.Y(n_1510)
);

AOI22x1_ASAP7_75t_L g1511 ( 
.A1(n_1329),
.A2(n_900),
.B1(n_876),
.B2(n_583),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1302),
.A2(n_754),
.B1(n_744),
.B2(n_664),
.C(n_1002),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1256),
.Y(n_1514)
);

AOI21x1_ASAP7_75t_SL g1515 ( 
.A1(n_1376),
.A2(n_1468),
.B(n_1394),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1372),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1471),
.A2(n_1481),
.B(n_1478),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1513),
.A2(n_1469),
.B1(n_1374),
.B2(n_1486),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1444),
.B(n_1421),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1380),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1374),
.A2(n_1405),
.B(n_1508),
.C(n_1371),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1405),
.A2(n_1396),
.B(n_1507),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1465),
.B(n_1482),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1471),
.A2(n_1466),
.B(n_1386),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1404),
.A2(n_1394),
.B(n_1396),
.C(n_1408),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1435),
.B(n_1499),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1411),
.A2(n_1398),
.B1(n_1410),
.B2(n_1460),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1385),
.Y(n_1528)
);

OA22x2_ASAP7_75t_L g1529 ( 
.A1(n_1431),
.A2(n_1415),
.B1(n_1412),
.B2(n_1445),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1501),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1499),
.B(n_1436),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1504),
.Y(n_1532)
);

OA22x2_ASAP7_75t_L g1533 ( 
.A1(n_1449),
.A2(n_1497),
.B1(n_1512),
.B2(n_1495),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1411),
.A2(n_1398),
.B1(n_1410),
.B2(n_1397),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1409),
.B(n_1501),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1433),
.A2(n_1383),
.B(n_1420),
.C(n_1446),
.Y(n_1536)
);

BUFx2_ASAP7_75t_SL g1537 ( 
.A(n_1380),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1477),
.A2(n_1483),
.B1(n_1466),
.B2(n_1470),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1375),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1483),
.B(n_1502),
.Y(n_1541)
);

AOI221x1_ASAP7_75t_SL g1542 ( 
.A1(n_1492),
.A2(n_1489),
.B1(n_1427),
.B2(n_1430),
.C(n_1509),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_1439),
.B(n_1373),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_L g1544 ( 
.A(n_1439),
.B(n_1373),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1390),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1470),
.A2(n_1511),
.B1(n_1433),
.B2(n_1379),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1458),
.A2(n_1389),
.B(n_1386),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1390),
.B(n_1403),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1488),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1400),
.B(n_1425),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1454),
.A2(n_1417),
.B(n_1510),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1470),
.A2(n_1434),
.B1(n_1406),
.B2(n_1451),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1434),
.A2(n_1406),
.B1(n_1514),
.B2(n_1428),
.Y(n_1554)
);

AOI21x1_ASAP7_75t_SL g1555 ( 
.A1(n_1422),
.A2(n_1503),
.B(n_1462),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1473),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1480),
.B(n_1484),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1408),
.B(n_1438),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_L g1560 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1472),
.B(n_1393),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1472),
.B(n_1393),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1448),
.A2(n_1395),
.B(n_1447),
.Y(n_1563)
);

OA22x2_ASAP7_75t_L g1564 ( 
.A1(n_1472),
.A2(n_1447),
.B1(n_1485),
.B2(n_1498),
.Y(n_1564)
);

O2A1O1Ixp5_ASAP7_75t_L g1565 ( 
.A1(n_1423),
.A2(n_1417),
.B(n_1418),
.C(n_1491),
.Y(n_1565)
);

NOR2xp67_ASAP7_75t_L g1566 ( 
.A(n_1437),
.B(n_1488),
.Y(n_1566)
);

OA22x2_ASAP7_75t_L g1567 ( 
.A1(n_1472),
.A2(n_1487),
.B1(n_1498),
.B2(n_1485),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1493),
.A2(n_1423),
.B1(n_1498),
.B2(n_1487),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1485),
.A2(n_1487),
.B1(n_1419),
.B2(n_1455),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1407),
.A2(n_1448),
.B(n_1432),
.C(n_1391),
.Y(n_1570)
);

OA22x2_ASAP7_75t_L g1571 ( 
.A1(n_1419),
.A2(n_1443),
.B1(n_1442),
.B2(n_1440),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1441),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1419),
.A2(n_1455),
.B1(n_1381),
.B2(n_1456),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1453),
.B(n_1429),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1395),
.A2(n_1381),
.B(n_1393),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1393),
.B(n_1488),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1407),
.A2(n_1391),
.B(n_1381),
.C(n_1490),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1452),
.B(n_1441),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1402),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1456),
.A2(n_1424),
.B1(n_1402),
.B2(n_1453),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_SL g1581 ( 
.A(n_1426),
.B(n_1457),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1494),
.A2(n_1510),
.B(n_1506),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1476),
.A2(n_1490),
.B(n_1387),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1476),
.A2(n_1479),
.B(n_1382),
.Y(n_1584)
);

O2A1O1Ixp5_ASAP7_75t_L g1585 ( 
.A1(n_1399),
.A2(n_1370),
.B(n_1377),
.C(n_1500),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1505),
.A2(n_1401),
.B(n_1461),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1450),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1416),
.A2(n_1377),
.B(n_1500),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1392),
.B(n_1459),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1416),
.B(n_1378),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1374),
.A2(n_1481),
.B(n_1478),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1468),
.A2(n_1513),
.B1(n_1469),
.B2(n_1374),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1374),
.A2(n_1481),
.B(n_1478),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1499),
.B(n_1444),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1507),
.C(n_1374),
.Y(n_1597)
);

AOI21x1_ASAP7_75t_SL g1598 ( 
.A1(n_1376),
.A2(n_1313),
.B(n_1321),
.Y(n_1598)
);

NOR2xp67_ASAP7_75t_L g1599 ( 
.A(n_1439),
.B(n_1373),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1507),
.C(n_1374),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1372),
.B(n_1496),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1469),
.C(n_1486),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1507),
.C(n_1374),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1435),
.B(n_1499),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1385),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1493),
.B(n_651),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1499),
.B(n_1444),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1468),
.A2(n_1513),
.B1(n_1469),
.B2(n_1374),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1458),
.A2(n_1389),
.B(n_1386),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1385),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1471),
.A2(n_1481),
.B(n_1478),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1372),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1468),
.A2(n_1513),
.B1(n_1469),
.B2(n_1374),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1499),
.B(n_1444),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1458),
.A2(n_1389),
.B(n_1386),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1504),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1372),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1499),
.B(n_1444),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1507),
.C(n_1374),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1468),
.A2(n_1513),
.B1(n_1469),
.B2(n_1374),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1471),
.A2(n_1481),
.B(n_1478),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1372),
.B(n_1496),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1435),
.B(n_1499),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1444),
.B(n_1421),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1530),
.B(n_1601),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1540),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1567),
.B(n_1535),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1574),
.B(n_1576),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1537),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1549),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1557),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1558),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1518),
.A2(n_1527),
.B1(n_1594),
.B2(n_1613),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1584),
.A2(n_1583),
.B(n_1577),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1556),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1622),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1559),
.Y(n_1644)
);

OA21x2_ASAP7_75t_L g1645 ( 
.A1(n_1584),
.A2(n_1565),
.B(n_1583),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1624),
.B(n_1561),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1516),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1548),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1562),
.B(n_1564),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1574),
.B(n_1589),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1579),
.Y(n_1651)
);

BUFx12f_ASAP7_75t_L g1652 ( 
.A(n_1520),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1565),
.A2(n_1524),
.B(n_1621),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1571),
.B(n_1575),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1577),
.A2(n_1621),
.B(n_1517),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1571),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1545),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1591),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1526),
.B(n_1604),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1597),
.A2(n_1600),
.B(n_1603),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1608),
.A2(n_1620),
.B1(n_1534),
.B2(n_1529),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1564),
.B(n_1617),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1517),
.A2(n_1611),
.B(n_1588),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1612),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1532),
.B(n_1539),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1612),
.B(n_1551),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1592),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1590),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1585),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1523),
.B(n_1573),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1610),
.B(n_1616),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1623),
.Y(n_1672)
);

BUFx2_ASAP7_75t_SL g1673 ( 
.A(n_1560),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1552),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1531),
.B(n_1528),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1593),
.B(n_1595),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1541),
.B(n_1605),
.Y(n_1677)
);

AO21x1_ASAP7_75t_SL g1678 ( 
.A1(n_1515),
.A2(n_1522),
.B(n_1521),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1570),
.A2(n_1536),
.B(n_1581),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1569),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1533),
.B(n_1568),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1602),
.A2(n_1619),
.B1(n_1603),
.B2(n_1600),
.C(n_1597),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1538),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1619),
.A2(n_1525),
.B(n_1563),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1580),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1554),
.B(n_1550),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1672),
.B(n_1542),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1669),
.A2(n_1553),
.B(n_1566),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1646),
.B(n_1533),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1646),
.B(n_1552),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1627),
.B(n_1547),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1627),
.B(n_1547),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1632),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1667),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1654),
.B(n_1650),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1628),
.B(n_1615),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1626),
.B(n_1615),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1626),
.B(n_1586),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1664),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1632),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1642),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1659),
.B(n_1586),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1676),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1642),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1630),
.B(n_1529),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1675),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1631),
.B(n_1582),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1652),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1640),
.A2(n_1546),
.B(n_1515),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1647),
.Y(n_1715)
);

OAI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1660),
.A2(n_1543),
.B(n_1544),
.C(n_1599),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1643),
.B(n_1582),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1650),
.B(n_1634),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1616),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1625),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1625),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1555),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1644),
.B(n_1598),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1666),
.B(n_1555),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1687),
.A2(n_1678),
.B1(n_1681),
.B2(n_1685),
.Y(n_1725)
);

OAI211xp5_ASAP7_75t_L g1726 ( 
.A1(n_1712),
.A2(n_1682),
.B(n_1660),
.C(n_1640),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1687),
.A2(n_1678),
.B1(n_1681),
.B2(n_1676),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_L g1728 ( 
.A(n_1712),
.B(n_1661),
.C(n_1683),
.Y(n_1728)
);

OAI211xp5_ASAP7_75t_L g1729 ( 
.A1(n_1723),
.A2(n_1661),
.B(n_1653),
.C(n_1645),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1692),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1658),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1695),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1706),
.B(n_1676),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

CKINVDCx16_ASAP7_75t_R g1735 ( 
.A(n_1708),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1691),
.B(n_1658),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1723),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1708),
.A2(n_1679),
.B1(n_1649),
.B2(n_1680),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1719),
.A2(n_1654),
.B1(n_1662),
.B2(n_1680),
.C(n_1656),
.Y(n_1739)
);

OAI321xp33_ASAP7_75t_L g1740 ( 
.A1(n_1719),
.A2(n_1654),
.A3(n_1649),
.B1(n_1662),
.B2(n_1706),
.C(n_1714),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1720),
.B(n_1648),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1689),
.A2(n_1654),
.B1(n_1656),
.B2(n_1679),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1691),
.B(n_1668),
.Y(n_1743)
);

AND4x1_ASAP7_75t_L g1744 ( 
.A(n_1689),
.B(n_1651),
.C(n_1665),
.D(n_1671),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1719),
.A2(n_1654),
.B1(n_1644),
.B2(n_1670),
.C(n_1633),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1693),
.B(n_1668),
.Y(n_1746)
);

BUFx10_ASAP7_75t_L g1747 ( 
.A(n_1711),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1693),
.B(n_1668),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1718),
.B(n_1634),
.Y(n_1749)
);

OAI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1706),
.A2(n_1686),
.B1(n_1670),
.B2(n_1633),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1705),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1720),
.B(n_1648),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1688),
.A2(n_1673),
.B1(n_1635),
.B2(n_1686),
.C(n_1653),
.Y(n_1753)
);

AO21x1_ASAP7_75t_SL g1754 ( 
.A1(n_1705),
.A2(n_1698),
.B(n_1701),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1694),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1694),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1703),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

OAI33xp33_ASAP7_75t_L g1759 ( 
.A1(n_1701),
.A2(n_1677),
.A3(n_1657),
.B1(n_1637),
.B2(n_1638),
.B3(n_1639),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1713),
.A2(n_1641),
.B(n_1655),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1703),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1697),
.B(n_1663),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1721),
.B(n_1657),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1737),
.B(n_1698),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1754),
.B(n_1690),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1726),
.B(n_1636),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1755),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1737),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1761),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1755),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1754),
.B(n_1690),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1730),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1728),
.B(n_1706),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1761),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1761),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1756),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1726),
.B(n_1716),
.C(n_1715),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_SL g1780 ( 
.A(n_1728),
.B(n_1724),
.C(n_1722),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1757),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1751),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1730),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1761),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1758),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1729),
.B(n_1724),
.C(n_1722),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1758),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1757),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1749),
.B(n_1718),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1762),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1763),
.B(n_1697),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1734),
.Y(n_1792)
);

INVx8_ASAP7_75t_L g1793 ( 
.A(n_1749),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1762),
.Y(n_1794)
);

AO21x1_ASAP7_75t_L g1795 ( 
.A1(n_1751),
.A2(n_1721),
.B(n_1717),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1729),
.B(n_1653),
.C(n_1702),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1763),
.B(n_1699),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1760),
.Y(n_1798)
);

OR2x6_ASAP7_75t_L g1799 ( 
.A(n_1749),
.B(n_1696),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1732),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1735),
.B(n_1706),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1786),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1767),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1789),
.B(n_1749),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1767),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1780),
.B(n_1741),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1786),
.B(n_1673),
.Y(n_1807)
);

INVx3_ASAP7_75t_SL g1808 ( 
.A(n_1793),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1789),
.B(n_1735),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1789),
.B(n_1699),
.Y(n_1810)
);

NOR3xp33_ASAP7_75t_L g1811 ( 
.A(n_1796),
.B(n_1753),
.C(n_1759),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1789),
.B(n_1700),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1768),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1769),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1768),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1789),
.B(n_1700),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1779),
.B(n_1727),
.Y(n_1817)
);

AND2x2_ASAP7_75t_SL g1818 ( 
.A(n_1779),
.B(n_1744),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1769),
.B(n_1725),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1766),
.B(n_1772),
.Y(n_1820)
);

NOR2xp67_ASAP7_75t_SL g1821 ( 
.A(n_1796),
.B(n_1652),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1799),
.B(n_1766),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1765),
.B(n_1741),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1766),
.B(n_1736),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1752),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1752),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1772),
.B(n_1743),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1791),
.B(n_1704),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1791),
.B(n_1797),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1797),
.B(n_1746),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1799),
.B(n_1663),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1707),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1793),
.B(n_1746),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1793),
.B(n_1748),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1771),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1771),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1765),
.B(n_1764),
.Y(n_1839)
);

AOI322xp5_ASAP7_75t_L g1840 ( 
.A1(n_1774),
.A2(n_1738),
.A3(n_1750),
.B1(n_1742),
.B2(n_1801),
.C1(n_1635),
.C2(n_1759),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1793),
.B(n_1748),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1793),
.B(n_1731),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1765),
.B(n_1764),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1799),
.B(n_1663),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1777),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1777),
.B(n_1778),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1809),
.B(n_1793),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1808),
.B(n_1809),
.Y(n_1848)
);

NAND2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1821),
.B(n_1587),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1819),
.B(n_1778),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1811),
.B(n_1738),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1845),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1807),
.B(n_1808),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1806),
.B(n_1781),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1818),
.B(n_1781),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1814),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1846),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1802),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1808),
.B(n_1747),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1806),
.B(n_1788),
.Y(n_1861)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1862 ( 
.A1(n_1817),
.A2(n_1795),
.B(n_1753),
.C(n_1774),
.D(n_1801),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1818),
.A2(n_1745),
.B1(n_1793),
.B2(n_1739),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1830),
.B(n_1788),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1846),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1813),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1839),
.B(n_1790),
.Y(n_1867)
);

NAND2x1p5_ASAP7_75t_L g1868 ( 
.A(n_1807),
.B(n_1744),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1813),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1815),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1818),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1803),
.A2(n_1745),
.B1(n_1739),
.B2(n_1799),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1840),
.A2(n_1740),
.B(n_1795),
.C(n_1733),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1815),
.Y(n_1874)
);

CKINVDCx16_ASAP7_75t_R g1875 ( 
.A(n_1822),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1837),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1837),
.Y(n_1877)
);

OAI21xp33_ASAP7_75t_L g1878 ( 
.A1(n_1840),
.A2(n_1783),
.B(n_1773),
.Y(n_1878)
);

NAND2x1_ASAP7_75t_L g1879 ( 
.A(n_1822),
.B(n_1800),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1805),
.B(n_1790),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1822),
.A2(n_1799),
.B1(n_1750),
.B2(n_1709),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1822),
.B(n_1820),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1804),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1820),
.B(n_1747),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1823),
.B(n_1794),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1882),
.B(n_1835),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1847),
.B(n_1835),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1866),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1850),
.Y(n_1889)
);

AOI222xp33_ASAP7_75t_L g1890 ( 
.A1(n_1859),
.A2(n_1850),
.B1(n_1852),
.B2(n_1871),
.C1(n_1878),
.C2(n_1873),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1871),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1868),
.Y(n_1892)
);

CKINVDCx16_ASAP7_75t_R g1893 ( 
.A(n_1875),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1869),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1859),
.B(n_1838),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1848),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1870),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1856),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1874),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1855),
.B(n_1823),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1861),
.B(n_1825),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1847),
.B(n_1836),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1857),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1883),
.B(n_1804),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1851),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1858),
.B(n_1831),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1867),
.B(n_1827),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1884),
.B(n_1836),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1864),
.B(n_1839),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1860),
.B(n_1841),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1883),
.B(n_1841),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1865),
.B(n_1831),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1853),
.B(n_1880),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1893),
.B(n_1854),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1889),
.B(n_1876),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1904),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1905),
.B(n_1885),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1889),
.B(n_1843),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1893),
.B(n_1832),
.Y(n_1919)
);

O2A1O1Ixp33_ASAP7_75t_SL g1920 ( 
.A1(n_1896),
.A2(n_1873),
.B(n_1879),
.C(n_1862),
.Y(n_1920)
);

AOI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1890),
.A2(n_1877),
.B(n_1821),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1891),
.B(n_1832),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_SL g1923 ( 
.A1(n_1891),
.A2(n_1854),
.B(n_1838),
.C(n_1800),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1891),
.B(n_1824),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1890),
.A2(n_1868),
.B1(n_1863),
.B2(n_1872),
.C(n_1849),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1896),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1903),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1888),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1887),
.B(n_1747),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1887),
.B(n_1747),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1909),
.B(n_1843),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1892),
.A2(n_1849),
.B1(n_1795),
.B2(n_1881),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1904),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1898),
.B(n_1824),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1892),
.Y(n_1935)
);

AOI31xp33_ASAP7_75t_L g1936 ( 
.A1(n_1892),
.A2(n_1842),
.A3(n_1826),
.B(n_1828),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1926),
.B(n_1900),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1914),
.B(n_1913),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1916),
.B(n_1902),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_R g1940 ( 
.A(n_1929),
.B(n_1910),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1916),
.B(n_1900),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1933),
.B(n_1902),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1919),
.B(n_1909),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1915),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1931),
.B(n_1911),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1922),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1918),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1930),
.B(n_1911),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1924),
.B(n_1908),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1927),
.B(n_1895),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1934),
.B(n_1908),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1938),
.B(n_1925),
.Y(n_1952)
);

AO21x1_ASAP7_75t_L g1953 ( 
.A1(n_1950),
.A2(n_1921),
.B(n_1915),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1938),
.B(n_1939),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1944),
.A2(n_1921),
.B1(n_1920),
.B2(n_1935),
.C(n_1932),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1886),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1944),
.A2(n_1923),
.B(n_1895),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1942),
.Y(n_1958)
);

AOI211xp5_ASAP7_75t_L g1959 ( 
.A1(n_1950),
.A2(n_1917),
.B(n_1886),
.C(n_1901),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1945),
.B(n_1910),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1947),
.A2(n_1904),
.B1(n_1901),
.B2(n_1912),
.Y(n_1961)
);

OAI211xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1937),
.A2(n_1928),
.B(n_1899),
.C(n_1888),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1947),
.B(n_1949),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1963),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1954),
.Y(n_1965)
);

AOI221x1_ASAP7_75t_L g1966 ( 
.A1(n_1962),
.A2(n_1941),
.B1(n_1946),
.B2(n_1943),
.C(n_1899),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1953),
.A2(n_1951),
.B1(n_1948),
.B2(n_1904),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1958),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1956),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1960),
.B(n_1936),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1964),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1965),
.B(n_1952),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1965),
.B(n_1959),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1969),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1967),
.B(n_1961),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1968),
.B(n_1957),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1970),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1966),
.B(n_1955),
.Y(n_1978)
);

AOI332xp33_ASAP7_75t_L g1979 ( 
.A1(n_1971),
.A2(n_1897),
.A3(n_1894),
.B1(n_1940),
.B2(n_1906),
.B3(n_1907),
.C1(n_1776),
.C2(n_1775),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1973),
.B(n_1907),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1978),
.A2(n_1897),
.B1(n_1894),
.B2(n_1844),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1972),
.B(n_1842),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1976),
.A2(n_1834),
.B(n_1829),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1974),
.Y(n_1984)
);

NOR3x2_ASAP7_75t_L g1985 ( 
.A(n_1980),
.B(n_1977),
.C(n_1984),
.Y(n_1985)
);

OAI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1981),
.A2(n_1975),
.B1(n_1784),
.B2(n_1770),
.C(n_1776),
.Y(n_1986)
);

NOR3xp33_ASAP7_75t_L g1987 ( 
.A(n_1983),
.B(n_1844),
.C(n_1833),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1982),
.A2(n_1776),
.B1(n_1770),
.B2(n_1775),
.C(n_1784),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1986),
.A2(n_1979),
.B1(n_1826),
.B2(n_1828),
.Y(n_1989)
);

NOR2x1_ASAP7_75t_L g1990 ( 
.A(n_1985),
.B(n_1800),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1989),
.A2(n_1987),
.B1(n_1988),
.B2(n_1810),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1990),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1992),
.B(n_1785),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1991),
.B(n_1785),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1994),
.B(n_1993),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1993),
.A2(n_1844),
.B(n_1833),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1995),
.Y(n_1997)
);

AO22x2_ASAP7_75t_L g1998 ( 
.A1(n_1996),
.A2(n_1844),
.B1(n_1833),
.B2(n_1770),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1998),
.B1(n_1810),
.B2(n_1816),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1775),
.B1(n_1784),
.B2(n_1833),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1816),
.B(n_1812),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_1812),
.B1(n_1785),
.B2(n_1787),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_2002),
.A2(n_1773),
.B1(n_1783),
.B2(n_1792),
.Y(n_2003)
);

AOI211xp5_ASAP7_75t_L g2004 ( 
.A1(n_2003),
.A2(n_1792),
.B(n_1798),
.C(n_1787),
.Y(n_2004)
);


endmodule