module real_aes_6855_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g501 ( .A(n_1), .Y(n_501) );
INVx1_ASAP7_75t_L g208 ( .A(n_2), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_3), .A2(n_37), .B1(n_169), .B2(n_531), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_4), .A2(n_150), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_5), .B(n_143), .Y(n_514) );
AND2x6_ASAP7_75t_L g155 ( .A(n_6), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_7), .A2(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_8), .B(n_38), .Y(n_467) );
INVx1_ASAP7_75t_L g183 ( .A(n_9), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_10), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g148 ( .A(n_11), .Y(n_148) );
INVx1_ASAP7_75t_L g495 ( .A(n_12), .Y(n_495) );
INVx1_ASAP7_75t_L g264 ( .A(n_13), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_14), .B(n_191), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_15), .B(n_144), .Y(n_572) );
AO32x2_ASAP7_75t_L g544 ( .A1(n_16), .A2(n_143), .A3(n_188), .B1(n_523), .B2(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_17), .A2(n_62), .B1(n_132), .B2(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_17), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_18), .B(n_169), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_19), .B(n_164), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_20), .B(n_144), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_21), .A2(n_50), .B1(n_169), .B2(n_531), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_22), .B(n_150), .Y(n_220) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_23), .A2(n_79), .B1(n_169), .B2(n_191), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_24), .B(n_169), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_25), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_26), .A2(n_262), .B(n_263), .C(n_265), .Y(n_261) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_27), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_28), .B(n_185), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_29), .B(n_181), .Y(n_210) );
INVx1_ASAP7_75t_L g197 ( .A(n_30), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_31), .A2(n_32), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_31), .Y(n_127) );
INVxp67_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_32), .B(n_185), .Y(n_561) );
INVx2_ASAP7_75t_L g153 ( .A(n_33), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_34), .B(n_169), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_35), .B(n_185), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_36), .A2(n_155), .B(n_159), .C(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_38), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g195 ( .A(n_39), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_40), .A2(n_475), .B1(n_478), .B2(n_479), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_40), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_41), .B(n_181), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_42), .B(n_169), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_43), .A2(n_90), .B1(n_227), .B2(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_44), .B(n_169), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_45), .B(n_169), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_46), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_47), .A2(n_69), .B1(n_476), .B2(n_477), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_47), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_48), .B(n_500), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_49), .B(n_150), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_51), .A2(n_60), .B1(n_169), .B2(n_191), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_52), .A2(n_159), .B1(n_191), .B2(n_193), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_53), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_54), .B(n_169), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_55), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_56), .B(n_169), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_57), .A2(n_168), .B(n_180), .C(n_182), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_58), .Y(n_240) );
INVx1_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
INVx1_ASAP7_75t_L g156 ( .A(n_61), .Y(n_156) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_63), .B(n_169), .Y(n_502) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_66), .A2(n_143), .A3(n_244), .B1(n_523), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g521 ( .A(n_67), .Y(n_521) );
INVx1_ASAP7_75t_L g556 ( .A(n_68), .Y(n_556) );
INVx1_ASAP7_75t_L g476 ( .A(n_69), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_SL g163 ( .A1(n_70), .A2(n_164), .B(n_165), .C(n_168), .Y(n_163) );
INVxp67_ASAP7_75t_L g166 ( .A(n_71), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_72), .B(n_191), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_73), .A2(n_473), .B1(n_474), .B2(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_73), .Y(n_473) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_75), .B(n_463), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_76), .A2(n_465), .B1(n_471), .B2(n_775), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_77), .Y(n_201) );
INVx1_ASAP7_75t_L g233 ( .A(n_78), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_80), .A2(n_155), .B(n_159), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_81), .B(n_531), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_82), .B(n_191), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_83), .A2(n_105), .B1(n_118), .B2(n_780), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_84), .B(n_209), .Y(n_223) );
INVx2_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_86), .B(n_164), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_87), .B(n_191), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_88), .A2(n_155), .B(n_159), .C(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g114 ( .A(n_89), .Y(n_114) );
OR2x2_ASAP7_75t_L g464 ( .A(n_89), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_91), .A2(n_103), .B1(n_191), .B2(n_192), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_92), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_93), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_94), .A2(n_155), .B(n_159), .C(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_95), .Y(n_254) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_97), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_98), .B(n_209), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_99), .B(n_191), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_100), .B(n_143), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_101), .B(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_102), .A2(n_150), .B(n_157), .Y(n_149) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx4f_ASAP7_75t_SL g780 ( .A(n_106), .Y(n_780) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g466 ( .A(n_113), .B(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_SL g481 ( .A1(n_114), .A2(n_134), .B1(n_482), .B2(n_774), .Y(n_481) );
INVx2_ASAP7_75t_L g774 ( .A(n_114), .Y(n_774) );
NOR2x2_ASAP7_75t_L g777 ( .A(n_114), .B(n_465), .Y(n_777) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_469), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g779 ( .A(n_122), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_461), .B(n_468), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_128), .B1(n_129), .B2(n_460), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_125), .Y(n_460) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B1(n_134), .B2(n_459), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g459 ( .A(n_134), .Y(n_459) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND4x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_377), .C(n_424), .D(n_444), .Y(n_135) );
NOR3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_307), .C(n_332), .Y(n_136) );
OAI211xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_215), .B(n_267), .C(n_297), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_186), .Y(n_139) );
INVx3_ASAP7_75t_SL g349 ( .A(n_140), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_140), .B(n_280), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_140), .B(n_202), .Y(n_430) );
AND2x2_ASAP7_75t_L g453 ( .A(n_140), .B(n_319), .Y(n_453) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_174), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g271 ( .A(n_142), .B(n_175), .Y(n_271) );
INVx3_ASAP7_75t_L g284 ( .A(n_142), .Y(n_284) );
AND2x2_ASAP7_75t_L g289 ( .A(n_142), .B(n_174), .Y(n_289) );
OR2x2_ASAP7_75t_L g340 ( .A(n_142), .B(n_281), .Y(n_340) );
BUFx2_ASAP7_75t_L g360 ( .A(n_142), .Y(n_360) );
AND2x2_ASAP7_75t_L g370 ( .A(n_142), .B(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g376 ( .A(n_142), .B(n_187), .Y(n_376) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_149), .B(n_171), .Y(n_142) );
INVx4_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_143), .A2(n_507), .B(n_514), .Y(n_506) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_145), .B(n_146), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx2_ASAP7_75t_L g258 ( .A(n_150), .Y(n_258) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_151), .B(n_155), .Y(n_199) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g500 ( .A(n_152), .Y(n_500) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
INVx1_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx1_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
INVx1_ASAP7_75t_L g164 ( .A(n_154), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
INVx4_ASAP7_75t_SL g170 ( .A(n_155), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_155), .A2(n_494), .B(n_498), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_511), .Y(n_507) );
BUFx3_ASAP7_75t_L g523 ( .A(n_155), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_155), .A2(n_536), .B(n_540), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_155), .A2(n_555), .B(n_558), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_162), .B(n_163), .C(n_170), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_170), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_158), .A2(n_170), .B(n_260), .C(n_261), .Y(n_259) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
BUFx3_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g531 ( .A(n_160), .Y(n_531) );
INVx1_ASAP7_75t_L g539 ( .A(n_164), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_167), .B(n_183), .Y(n_182) );
INVx5_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g529 ( .A1(n_167), .A2(n_181), .B1(n_530), .B2(n_532), .Y(n_529) );
O2A1O1Ixp5_ASAP7_75t_SL g555 ( .A1(n_168), .A2(n_209), .B(n_556), .C(n_557), .Y(n_555) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_169), .Y(n_251) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_170), .A2(n_190), .B1(n_198), .B2(n_199), .Y(n_189) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_172), .A2(n_176), .B(n_184), .Y(n_175) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_173), .B(n_230), .Y(n_229) );
AO21x1_ASAP7_75t_L g567 ( .A1(n_173), .A2(n_568), .B(n_571), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_173), .B(n_523), .C(n_568), .Y(n_586) );
INVx1_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_175), .B(n_281), .Y(n_295) );
INVx2_ASAP7_75t_L g305 ( .A(n_175), .Y(n_305) );
AND2x2_ASAP7_75t_L g318 ( .A(n_175), .B(n_284), .Y(n_318) );
OR2x2_ASAP7_75t_L g329 ( .A(n_175), .B(n_281), .Y(n_329) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_175), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g387 ( .A(n_175), .Y(n_387) );
AND2x2_ASAP7_75t_L g433 ( .A(n_175), .B(n_187), .Y(n_433) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_180), .A2(n_499), .B(n_521), .C(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_180), .A2(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g250 ( .A(n_181), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_181), .A2(n_503), .B1(n_546), .B2(n_547), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_181), .A2(n_503), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g214 ( .A(n_185), .Y(n_214) );
INVx2_ASAP7_75t_L g244 ( .A(n_185), .Y(n_244) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_185), .A2(n_257), .B(n_266), .Y(n_256) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_185), .A2(n_535), .B(n_543), .Y(n_534) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_185), .A2(n_554), .B(n_561), .Y(n_553) );
INVx3_ASAP7_75t_SL g306 ( .A(n_186), .Y(n_306) );
OR2x2_ASAP7_75t_L g359 ( .A(n_186), .B(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_202), .Y(n_186) );
INVx3_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
AND2x2_ASAP7_75t_L g348 ( .A(n_187), .B(n_203), .Y(n_348) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_187), .Y(n_416) );
AOI33xp33_ASAP7_75t_L g420 ( .A1(n_187), .A2(n_349), .A3(n_356), .B1(n_365), .B2(n_421), .B3(n_422), .Y(n_420) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_200), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_188), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_188), .A2(n_204), .B(n_212), .Y(n_203) );
INVx2_ASAP7_75t_L g228 ( .A(n_188), .Y(n_228) );
INVx2_ASAP7_75t_L g211 ( .A(n_191), .Y(n_211) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_195), .B1(n_196), .B2(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g196 ( .A(n_194), .Y(n_196) );
INVx4_ASAP7_75t_L g262 ( .A(n_194), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_199), .A2(n_205), .B(n_206), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_199), .A2(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_202), .B(n_284), .Y(n_283) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_202), .B(n_344), .C(n_346), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_202), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_202), .B(n_376), .Y(n_379) );
AND2x2_ASAP7_75t_L g432 ( .A(n_202), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
OR2x2_ASAP7_75t_L g382 ( .A(n_203), .B(n_281), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .C(n_211), .Y(n_207) );
INVx2_ASAP7_75t_L g503 ( .A(n_209), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_209), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_209), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_211), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_214), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_214), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_241), .Y(n_215) );
AOI32xp33_ASAP7_75t_L g333 ( .A1(n_216), .A2(n_334), .A3(n_336), .B1(n_338), .B2(n_341), .Y(n_333) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_216), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g436 ( .A(n_216), .Y(n_436) );
INVx4_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g368 ( .A(n_217), .B(n_352), .Y(n_368) );
AND2x2_ASAP7_75t_L g388 ( .A(n_217), .B(n_314), .Y(n_388) );
AND2x2_ASAP7_75t_L g456 ( .A(n_217), .B(n_374), .Y(n_456) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx3_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_275), .Y(n_291) );
OR2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_274), .Y(n_296) );
INVx1_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
AND2x2_ASAP7_75t_L g311 ( .A(n_218), .B(n_285), .Y(n_311) );
AND2x2_ASAP7_75t_L g313 ( .A(n_218), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_218), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g366 ( .A(n_218), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_218), .B(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_228), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_225), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_228), .A2(n_493), .B(n_504), .Y(n_492) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_228), .A2(n_516), .B(n_524), .Y(n_515) );
INVx2_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
AND2x2_ASAP7_75t_L g321 ( .A(n_231), .B(n_242), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_231), .B(n_256), .Y(n_331) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
INVx2_ASAP7_75t_L g451 ( .A(n_241), .Y(n_451) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_255), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_242), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g292 ( .A(n_242), .Y(n_292) );
AND2x2_ASAP7_75t_L g336 ( .A(n_242), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g352 ( .A(n_242), .B(n_315), .Y(n_352) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_243), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g365 ( .A(n_243), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_243), .B(n_275), .Y(n_397) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_253), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_252), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_251), .Y(n_247) );
AND2x2_ASAP7_75t_L g276 ( .A(n_255), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_255), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g374 ( .A(n_255), .Y(n_374) );
INVx1_ASAP7_75t_L g407 ( .A(n_255), .Y(n_407) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g285 ( .A(n_256), .B(n_275), .Y(n_285) );
INVx1_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_262), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g497 ( .A(n_262), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_262), .A2(n_559), .B(n_560), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B1(n_278), .B2(n_285), .C(n_286), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_269), .B(n_289), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_269), .B(n_352), .Y(n_429) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_271), .B(n_319), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_271), .B(n_280), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_271), .B(n_294), .Y(n_423) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g345 ( .A(n_275), .Y(n_345) );
AND2x2_ASAP7_75t_L g320 ( .A(n_276), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g398 ( .A(n_276), .Y(n_398) );
AND2x2_ASAP7_75t_L g330 ( .A(n_277), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_277), .B(n_300), .Y(n_346) );
AND2x2_ASAP7_75t_L g410 ( .A(n_277), .B(n_336), .Y(n_410) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_288), .Y(n_319) );
AND2x2_ASAP7_75t_L g415 ( .A(n_282), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_284), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_285), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_285), .B(n_292), .Y(n_380) );
AND2x2_ASAP7_75t_L g400 ( .A(n_285), .B(n_300), .Y(n_400) );
AND2x2_ASAP7_75t_L g421 ( .A(n_285), .B(n_365), .Y(n_421) );
OAI32xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .A3(n_292), .B1(n_293), .B2(n_296), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_SL g294 ( .A(n_288), .Y(n_294) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_288), .B(n_318), .Y(n_335) );
OR2x2_ASAP7_75t_L g339 ( .A(n_288), .B(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_288), .B(n_387), .Y(n_440) );
INVx1_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
OAI221xp5_ASAP7_75t_SL g426 ( .A1(n_290), .A2(n_381), .B1(n_427), .B2(n_430), .C(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_291), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g341 ( .A(n_291), .B(n_314), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_291), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_291), .B(n_352), .Y(n_419) );
INVxp67_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g425 ( .A(n_294), .B(n_412), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_294), .B(n_375), .Y(n_448) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_296), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g441 ( .A(n_296), .B(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_301), .B(n_304), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_299), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g394 ( .A(n_303), .B(n_314), .Y(n_394) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g412 ( .A(n_305), .B(n_370), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_305), .B(n_369), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_306), .B(n_318), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_312), .C(n_322), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_308), .A2(n_343), .B1(n_347), .B2(n_350), .C(n_353), .Y(n_342) );
AOI31xp33_ASAP7_75t_L g437 ( .A1(n_308), .A2(n_438), .A3(n_439), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B1(n_318), .B2(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g438 ( .A(n_318), .Y(n_438) );
INVx1_ASAP7_75t_L g401 ( .A(n_319), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g444 ( .A1(n_321), .A2(n_445), .B(n_447), .C(n_449), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_326), .B2(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_327), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_329), .A2(n_363), .B1(n_382), .B2(n_418), .C(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g413 ( .A(n_330), .Y(n_413) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
NAND3xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_342), .C(n_357), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_334), .A2(n_384), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_336), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g443 ( .A(n_337), .Y(n_443) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g381 ( .A(n_344), .B(n_364), .Y(n_381) );
INVx1_ASAP7_75t_L g356 ( .A(n_345), .Y(n_356) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g354 ( .A(n_348), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_348), .B(n_386), .Y(n_385) );
NOR4xp25_ASAP7_75t_L g353 ( .A(n_349), .B(n_354), .C(n_355), .D(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B1(n_368), .B2(n_369), .C1(n_371), .C2(n_375), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g455 ( .A(n_359), .Y(n_455) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_371), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_376), .A2(n_432), .B(n_434), .Y(n_431) );
NOR4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_389), .C(n_402), .D(n_417), .Y(n_377) );
OAI221xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_380), .B1(n_381), .B2(n_382), .C(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_386), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B1(n_395), .B2(n_396), .C1(n_399), .C2(n_401), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_394), .A2(n_425), .B(n_426), .C(n_437), .Y(n_424) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
OAI222xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_408), .B1(n_409), .B2(n_411), .C1(n_413), .C2(n_414), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_419), .A2(n_422), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_452), .B(n_454), .C(n_457), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_468), .A2(n_470), .B(n_778), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_474), .Y(n_480) );
INVx1_ASAP7_75t_L g478 ( .A(n_475), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_484), .B(n_740), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_644), .C(n_728), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_587), .C(n_609), .D(n_625), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_525), .B1(n_548), .B2(n_566), .C(n_573), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_505), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_489), .B(n_566), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_489), .B(n_627), .C(n_640), .D(n_642), .Y(n_639) );
INVxp67_ASAP7_75t_L g756 ( .A(n_489), .Y(n_756) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g638 ( .A(n_490), .B(n_576), .Y(n_638) );
AND2x2_ASAP7_75t_L g662 ( .A(n_490), .B(n_505), .Y(n_662) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g629 ( .A(n_491), .B(n_565), .Y(n_629) );
AND2x2_ASAP7_75t_L g669 ( .A(n_491), .B(n_650), .Y(n_669) );
AND2x2_ASAP7_75t_L g686 ( .A(n_491), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_491), .B(n_506), .Y(n_710) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g593 ( .A(n_492), .B(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_492), .B(n_515), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_501), .B(n_502), .C(n_503), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_503), .A2(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g596 ( .A(n_505), .B(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_505), .A2(n_646), .B1(n_649), .B2(n_651), .C(n_655), .Y(n_645) );
AND2x2_ASAP7_75t_L g704 ( .A(n_505), .B(n_669), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_505), .B(n_686), .Y(n_738) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx3_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
AND2x2_ASAP7_75t_L g613 ( .A(n_506), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g667 ( .A(n_506), .B(n_582), .Y(n_667) );
AND2x2_ASAP7_75t_L g725 ( .A(n_506), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g582 ( .A(n_515), .Y(n_582) );
INVx1_ASAP7_75t_L g637 ( .A(n_515), .Y(n_637) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_515), .Y(n_643) );
AND2x2_ASAP7_75t_L g688 ( .A(n_515), .B(n_565), .Y(n_688) );
OR2x2_ASAP7_75t_L g727 ( .A(n_515), .B(n_567), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_520), .B(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_525), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_533), .Y(n_525) );
AND2x2_ASAP7_75t_L g723 ( .A(n_526), .B(n_720), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_526), .B(n_705), .Y(n_755) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g654 ( .A(n_527), .B(n_578), .Y(n_654) );
AND2x2_ASAP7_75t_L g703 ( .A(n_527), .B(n_551), .Y(n_703) );
INVx1_ASAP7_75t_L g749 ( .A(n_527), .Y(n_749) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_528), .Y(n_563) );
AND2x2_ASAP7_75t_L g604 ( .A(n_528), .B(n_578), .Y(n_604) );
INVx1_ASAP7_75t_L g621 ( .A(n_528), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_528), .B(n_544), .Y(n_627) );
AND2x2_ASAP7_75t_L g695 ( .A(n_533), .B(n_603), .Y(n_695) );
INVx2_ASAP7_75t_L g760 ( .A(n_533), .Y(n_760) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_544), .Y(n_533) );
AND2x2_ASAP7_75t_L g577 ( .A(n_534), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_552), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_534), .B(n_551), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_534), .Y(n_624) );
INVx1_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_534), .Y(n_653) );
INVx2_ASAP7_75t_L g721 ( .A(n_534), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
BUFx2_ASAP7_75t_L g675 ( .A(n_544), .Y(n_675) );
AND2x2_ASAP7_75t_L g720 ( .A(n_544), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_550), .B(n_657), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_550), .A2(n_719), .B(n_733), .Y(n_743) );
AND2x2_ASAP7_75t_L g768 ( .A(n_550), .B(n_654), .Y(n_768) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g690 ( .A(n_552), .Y(n_690) );
AND2x2_ASAP7_75t_L g719 ( .A(n_552), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
INVx2_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g576 ( .A(n_563), .Y(n_576) );
OR2x2_ASAP7_75t_L g589 ( .A(n_563), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g657 ( .A(n_563), .B(n_653), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_563), .B(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g758 ( .A(n_563), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_563), .B(n_695), .Y(n_770) );
AND2x2_ASAP7_75t_L g649 ( .A(n_564), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g672 ( .A(n_564), .B(n_566), .Y(n_672) );
INVx2_ASAP7_75t_L g584 ( .A(n_565), .Y(n_584) );
AND2x2_ASAP7_75t_L g612 ( .A(n_565), .B(n_585), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_565), .B(n_637), .Y(n_693) );
AND2x2_ASAP7_75t_L g607 ( .A(n_566), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g754 ( .A(n_566), .Y(n_754) );
AND2x2_ASAP7_75t_L g766 ( .A(n_566), .B(n_629), .Y(n_766) );
AND2x2_ASAP7_75t_L g592 ( .A(n_567), .B(n_582), .Y(n_592) );
INVx1_ASAP7_75t_L g687 ( .A(n_567), .Y(n_687) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_576), .B(n_623), .Y(n_632) );
OR2x2_ASAP7_75t_L g764 ( .A(n_576), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g681 ( .A(n_577), .B(n_622), .Y(n_681) );
AND2x2_ASAP7_75t_L g689 ( .A(n_577), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g748 ( .A(n_577), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g772 ( .A(n_577), .B(n_619), .Y(n_772) );
NOR2xp67_ASAP7_75t_L g730 ( .A(n_578), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g759 ( .A(n_578), .B(n_622), .Y(n_759) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g611 ( .A(n_581), .B(n_612), .Y(n_611) );
INVxp67_ASAP7_75t_L g773 ( .A(n_581), .Y(n_773) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g608 ( .A(n_584), .Y(n_608) );
AND2x2_ASAP7_75t_L g659 ( .A(n_584), .B(n_592), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_584), .B(n_727), .Y(n_753) );
INVx2_ASAP7_75t_L g598 ( .A(n_585), .Y(n_598) );
INVx3_ASAP7_75t_L g650 ( .A(n_585), .Y(n_650) );
OR2x2_ASAP7_75t_L g678 ( .A(n_585), .B(n_679), .Y(n_678) );
AOI311xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .A3(n_593), .B(n_594), .C(n_605), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_588), .A2(n_626), .B(n_628), .C(n_630), .Y(n_625) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g610 ( .A(n_590), .Y(n_610) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g628 ( .A(n_592), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_592), .B(n_608), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_592), .B(n_593), .Y(n_761) );
AND2x2_ASAP7_75t_L g683 ( .A(n_593), .B(n_597), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B(n_600), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g741 ( .A(n_597), .B(n_629), .Y(n_741) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_598), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g635 ( .A(n_598), .Y(n_635) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g626 ( .A(n_602), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g671 ( .A(n_604), .Y(n_671) );
AND2x4_ASAP7_75t_L g733 ( .A(n_604), .B(n_702), .Y(n_733) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_607), .A2(n_673), .B1(n_685), .B2(n_689), .C1(n_691), .C2(n_695), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_613), .C(n_616), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_610), .B(n_654), .Y(n_677) );
INVx1_ASAP7_75t_L g699 ( .A(n_612), .Y(n_699) );
INVx1_ASAP7_75t_L g633 ( .A(n_614), .Y(n_633) );
OR2x2_ASAP7_75t_L g698 ( .A(n_615), .B(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .B(n_623), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_617), .B(n_635), .C(n_636), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_617), .A2(n_654), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_621), .Y(n_674) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_622), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_622), .Y(n_747) );
INVx2_ASAP7_75t_L g705 ( .A(n_623), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_627), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g679 ( .A(n_629), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_634), .B2(n_638), .C(n_639), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_633), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g767 ( .A(n_633), .Y(n_767) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g648 ( .A(n_640), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_640), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g706 ( .A(n_640), .B(n_654), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_640), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g739 ( .A(n_640), .B(n_674), .Y(n_739) );
BUFx3_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_684), .D(n_696), .E(n_711), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI32xp33_ASAP7_75t_L g736 ( .A1(n_648), .A2(n_675), .A3(n_691), .B1(n_737), .B2(n_739), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_650), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g660 ( .A(n_654), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_670), .B1(n_672), .B2(n_673), .C(n_676), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g735 ( .A(n_667), .B(n_686), .Y(n_735) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_672), .A2(n_733), .B1(n_751), .B2(n_756), .C(n_757), .Y(n_750) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx2_ASAP7_75t_L g716 ( .A(n_675), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g694 ( .A(n_686), .Y(n_694) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_707), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_705), .A2(n_752), .B1(n_754), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .B(n_724), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g765 ( .A(n_720), .Y(n_765) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B(n_734), .C(n_736), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B(n_744), .C(n_769), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_741), .Y(n_745) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_750), .C(n_762), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_761), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
endmodule