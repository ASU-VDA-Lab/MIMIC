module fake_netlist_5_1141_n_2812 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2812);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2812;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1556;
wire n_1384;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2320;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2424;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2650;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2415;
wire n_2309;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_2429;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2282;
wire n_2002;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2377;
wire n_2080;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2437;
wire n_2219;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_293),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_156),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_314),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_17),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_271),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_351),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_131),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_597),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_256),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_239),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_443),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_587),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_388),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_19),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_264),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_510),
.Y(n_644)
);

CKINVDCx11_ASAP7_75t_R g645 ( 
.A(n_386),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_475),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_540),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_326),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_535),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_144),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_184),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_179),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_51),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_194),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_530),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_341),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_171),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_457),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_75),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_44),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_389),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_138),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_16),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_315),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_483),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_20),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_0),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_508),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_104),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_284),
.Y(n_670)
);

CKINVDCx14_ASAP7_75t_R g671 ( 
.A(n_471),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_134),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_22),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_278),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_73),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_617),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_218),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_167),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_91),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_413),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_295),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_207),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_148),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_513),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_581),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_599),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_301),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_422),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_61),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_37),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_433),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_434),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_425),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_85),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_502),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_262),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_570),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_353),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_621),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_102),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_579),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_249),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_379),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_367),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_22),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_345),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_489),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_534),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_492),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_319),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_148),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_30),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_17),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_578),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_178),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_410),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_166),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_528),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_519),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_211),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_214),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_188),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_596),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_503),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_411),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_20),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_382),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_624),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_133),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_448),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_569),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_218),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_39),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_583),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_628),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_533),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_377),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_565),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_456),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_585),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_240),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_612),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_142),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_524),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_232),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_568),
.Y(n_747)
);

INVxp67_ASAP7_75t_SL g748 ( 
.A(n_417),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_623),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_38),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_48),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_121),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_130),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_555),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_396),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_6),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_276),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_611),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_29),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_511),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_222),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_546),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_313),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_608),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_539),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_381),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_273),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_431),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_257),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_473),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_324),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_566),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_110),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_592),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_43),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_531),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_472),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_453),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_111),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_625),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_337),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_512),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_543),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_277),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_133),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_419),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_549),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_372),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_454),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_298),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_547),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_141),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_577),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_603),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_591),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_620),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_16),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_446),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_232),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_165),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_409),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_598),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_62),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_275),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_605),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_256),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_480),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_576),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_516),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_553),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_308),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_572),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_334),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_290),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_506),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_461),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_338),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_373),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_0),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_525),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_188),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_111),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_47),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_273),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_344),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_541),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_287),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_152),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_436),
.Y(n_830)
);

BUFx10_ASAP7_75t_L g831 ( 
.A(n_451),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_140),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_122),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_501),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_486),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_126),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_168),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_468),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_222),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_498),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_61),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_416),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_536),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_622),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_92),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_550),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_469),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_349),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_199),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_521),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_606),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_557),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_602),
.Y(n_853)
);

BUFx2_ASAP7_75t_SL g854 ( 
.A(n_101),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_230),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_99),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_488),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_354),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_556),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_269),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_183),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_269),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_66),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_496),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_3),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_33),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_5),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_167),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_44),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_144),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_415),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_286),
.Y(n_872)
);

CKINVDCx16_ASAP7_75t_R g873 ( 
.A(n_470),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_507),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_62),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_614),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_346),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_98),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_37),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_4),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_593),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_178),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_113),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_522),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_532),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_192),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_277),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_610),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_327),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_445),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_262),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_590),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_112),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_493),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_106),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_23),
.Y(n_896)
);

BUFx10_ASAP7_75t_L g897 ( 
.A(n_259),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_80),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_358),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_395),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_267),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_398),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_467),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_616),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_542),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_527),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_615),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_212),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_125),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_40),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_517),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_271),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_584),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_103),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_123),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_300),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_336),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_211),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_518),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_272),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_561),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_52),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_383),
.Y(n_923)
);

CKINVDCx16_ASAP7_75t_R g924 ( 
.A(n_123),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_203),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_221),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_134),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_28),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_82),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_138),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_57),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_427),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_497),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_404),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_288),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_247),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_267),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_552),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_574),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_481),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_255),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_81),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_428),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_328),
.Y(n_944)
);

INVxp33_ASAP7_75t_SL g945 ( 
.A(n_523),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_438),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_122),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_177),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_48),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_23),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_586),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_217),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_50),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_85),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_12),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_435),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_258),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_14),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_90),
.Y(n_959)
);

CKINVDCx11_ASAP7_75t_R g960 ( 
.A(n_279),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_226),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_186),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_202),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_613),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_66),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_187),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_94),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_175),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_32),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_505),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_50),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_156),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_573),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_476),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_495),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_399),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_594),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_46),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_261),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_30),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_7),
.Y(n_981)
);

CKINVDCx16_ASAP7_75t_R g982 ( 
.A(n_504),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_207),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_478),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_494),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_357),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_537),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_68),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_51),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_560),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_479),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_289),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_281),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_87),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_112),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_105),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_184),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_432),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_265),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_551),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_7),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_169),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_544),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_216),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_253),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_176),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_490),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_95),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_323),
.Y(n_1009)
);

BUFx8_ASAP7_75t_SL g1010 ( 
.A(n_515),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_335),
.Y(n_1011)
);

CKINVDCx16_ASAP7_75t_R g1012 ( 
.A(n_238),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_209),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_514),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_439),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_140),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_609),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_229),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_580),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_408),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_67),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_365),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_165),
.Y(n_1023)
);

CKINVDCx16_ASAP7_75t_R g1024 ( 
.A(n_310),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_113),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_589),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_249),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_582),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_78),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_230),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_474),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_39),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_216),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_105),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_491),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_418),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_191),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_499),
.Y(n_1038)
);

CKINVDCx14_ASAP7_75t_R g1039 ( 
.A(n_618),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_359),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_588),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_321),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_374),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_529),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_200),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_11),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_129),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_526),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_509),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_302),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_562),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_482),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_563),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_487),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_202),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_601),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_32),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_559),
.Y(n_1058)
);

BUFx8_ASAP7_75t_SL g1059 ( 
.A(n_225),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_333),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_567),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_274),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_604),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_558),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_265),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_213),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_545),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_538),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_463),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_155),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_206),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_392),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_153),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_131),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_24),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_21),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_33),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_564),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_121),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_548),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_170),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_520),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_600),
.Y(n_1083)
);

BUFx5_ASAP7_75t_L g1084 ( 
.A(n_75),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_179),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_316),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_268),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_440),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_84),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_57),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_35),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_58),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_330),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_294),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_191),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_485),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_215),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_500),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_378),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_59),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_152),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_607),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_129),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_362),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_331),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_190),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_477),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_166),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_291),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_96),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_484),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_401),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_299),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_215),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_571),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_12),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_221),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_554),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_575),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_11),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_430),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_126),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_173),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_852),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_652),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_652),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_960),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_652),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_689),
.B(n_1),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_852),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_730),
.B(n_1),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_852),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_652),
.B(n_2),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_652),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_652),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_839),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_839),
.Y(n_1137)
);

BUFx12f_ASAP7_75t_L g1138 ( 
.A(n_960),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_696),
.B(n_785),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_652),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1084),
.B(n_2),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_839),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1084),
.B(n_3),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_839),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_875),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_858),
.B(n_4),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1033),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_858),
.B(n_5),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1033),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1033),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1059),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_766),
.B(n_6),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_889),
.B(n_8),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1018),
.B(n_8),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_709),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1084),
.Y(n_1156)
);

INVx6_ASAP7_75t_L g1157 ( 
.A(n_740),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1084),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1084),
.B(n_9),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1084),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1084),
.B(n_9),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_852),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1033),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1077),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_709),
.B(n_10),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_723),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_723),
.B(n_10),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_820),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_864),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1122),
.B(n_657),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_695),
.B(n_13),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1077),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_864),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_945),
.B(n_13),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1082),
.B(n_14),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_656),
.B(n_15),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1077),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1059),
.Y(n_1179)
);

BUFx12f_ASAP7_75t_L g1180 ( 
.A(n_820),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_657),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_864),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_667),
.B(n_15),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_864),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_658),
.B(n_18),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_656),
.B(n_18),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_667),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_902),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_737),
.B(n_19),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_688),
.B(n_742),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_705),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_688),
.B(n_21),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_705),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_866),
.B(n_24),
.Y(n_1194)
);

INVx5_ASAP7_75t_L g1195 ( 
.A(n_902),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_866),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_949),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_949),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_737),
.B(n_25),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1045),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1045),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_902),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_675),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_742),
.B(n_25),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_902),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_820),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_806),
.B(n_26),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_975),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_975),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_675),
.B(n_711),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_975),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_763),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_975),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_924),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_897),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_847),
.B(n_26),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_897),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_651),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_763),
.B(n_876),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_876),
.B(n_27),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_897),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1001),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_1001),
.Y(n_1223)
);

BUFx8_ASAP7_75t_L g1224 ( 
.A(n_711),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_836),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_636),
.B(n_27),
.Y(n_1226)
);

AND2x6_ASAP7_75t_L g1227 ( 
.A(n_986),
.B(n_280),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_847),
.B(n_28),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1001),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_629),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_646),
.B(n_29),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_986),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_906),
.B(n_31),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_836),
.B(n_31),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_986),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_906),
.B(n_34),
.Y(n_1236)
);

AND2x6_ASAP7_75t_L g1237 ( 
.A(n_986),
.B(n_282),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_1020),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_874),
.B(n_34),
.Y(n_1239)
);

BUFx8_ASAP7_75t_L g1240 ( 
.A(n_909),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_909),
.B(n_35),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_947),
.B(n_36),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_893),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_648),
.B(n_36),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1087),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_661),
.B(n_38),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_653),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_947),
.B(n_40),
.Y(n_1248)
);

INVx5_ASAP7_75t_L g1249 ( 
.A(n_1020),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1020),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1020),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1051),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1051),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1012),
.B(n_41),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_668),
.B(n_41),
.Y(n_1255)
);

CKINVDCx16_ASAP7_75t_R g1256 ( 
.A(n_1090),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_671),
.B(n_42),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1087),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1120),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_978),
.B(n_42),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_663),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_978),
.B(n_43),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1040),
.B(n_45),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_666),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_999),
.B(n_45),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_687),
.B(n_46),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_999),
.Y(n_1267)
);

AND2x6_ASAP7_75t_L g1268 ( 
.A(n_1051),
.B(n_283),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1051),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1113),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1087),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1113),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_681),
.B(n_47),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_671),
.B(n_49),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_669),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_1010),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1085),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_684),
.B(n_693),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_682),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1039),
.B(n_49),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1085),
.B(n_52),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_699),
.B(n_53),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_740),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1113),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1039),
.B(n_53),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_683),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_812),
.B(n_54),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_740),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_936),
.B(n_54),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1113),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_744),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_965),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_971),
.B(n_55),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1123),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1285),
.A2(n_734),
.B1(n_873),
.B2(n_761),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1230),
.B(n_714),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1136),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1257),
.A2(n_982),
.B1(n_1069),
.B2(n_1024),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1256),
.A2(n_860),
.B1(n_868),
.B2(n_638),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1170),
.B(n_903),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1136),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1170),
.B(n_744),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1137),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1163),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1283),
.B(n_744),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1214),
.B(n_1215),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1139),
.B(n_872),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1177),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1285),
.A2(n_835),
.B1(n_859),
.B2(n_680),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1137),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1145),
.A2(n_1092),
.B1(n_632),
.B2(n_721),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1152),
.A2(n_835),
.B1(n_859),
.B2(n_680),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1153),
.A2(n_1274),
.B1(n_1280),
.B2(n_1174),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1146),
.A2(n_698),
.B1(n_716),
.B2(n_686),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1148),
.A2(n_736),
.B1(n_813),
.B2(n_724),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1145),
.A2(n_750),
.B1(n_829),
.B2(n_720),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1142),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1288),
.B(n_792),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1142),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1266),
.A2(n_933),
.B1(n_970),
.B2(n_913),
.Y(n_1320)
);

AO22x2_ASAP7_75t_L g1321 ( 
.A1(n_1129),
.A2(n_1114),
.B1(n_968),
.B2(n_854),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1155),
.B(n_792),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1144),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1144),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1243),
.A2(n_878),
.B1(n_901),
.B2(n_870),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1254),
.A2(n_1032),
.B1(n_633),
.B2(n_635),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1147),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1166),
.B(n_792),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1147),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1127),
.B(n_712),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1212),
.B(n_831),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1287),
.A2(n_1072),
.B1(n_1088),
.B2(n_1031),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_R g1333 ( 
.A1(n_1168),
.A2(n_1025),
.B1(n_1023),
.B2(n_1004),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1157),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1197),
.B(n_831),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1181),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1197),
.B(n_831),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1217),
.B(n_840),
.Y(n_1338)
);

AO22x2_ASAP7_75t_L g1339 ( 
.A1(n_1129),
.A2(n_1154),
.B1(n_1131),
.B2(n_1289),
.Y(n_1339)
);

AO22x2_ASAP7_75t_L g1340 ( 
.A1(n_1154),
.A2(n_746),
.B1(n_751),
.B2(n_717),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1138),
.B(n_754),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1149),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1149),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1221),
.B(n_1055),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1222),
.B(n_630),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1157),
.A2(n_642),
.B1(n_643),
.B2(n_637),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_SL g1347 ( 
.A(n_1291),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1219),
.B(n_840),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1171),
.B(n_984),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1150),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1150),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1175),
.A2(n_654),
.B1(n_659),
.B2(n_650),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1181),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1164),
.Y(n_1355)
);

AO22x2_ASAP7_75t_L g1356 ( 
.A1(n_1289),
.A2(n_774),
.B1(n_776),
.B2(n_757),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1190),
.A2(n_662),
.B1(n_672),
.B2(n_660),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1139),
.A2(n_1094),
.B1(n_673),
.B2(n_677),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1243),
.A2(n_674),
.B1(n_679),
.B2(n_678),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1185),
.B(n_1086),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1229),
.B(n_690),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1133),
.A2(n_700),
.B1(n_702),
.B2(n_694),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1292),
.A2(n_1259),
.B1(n_1271),
.B2(n_1245),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1293),
.A2(n_713),
.B1(n_722),
.B2(n_715),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1191),
.B(n_1187),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1176),
.A2(n_726),
.B1(n_732),
.B2(n_729),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1164),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1172),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1207),
.A2(n_860),
.B1(n_868),
.B2(n_638),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1293),
.A2(n_733),
.B1(n_753),
.B2(n_743),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1187),
.B(n_758),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1239),
.A2(n_762),
.B1(n_768),
.B2(n_760),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1263),
.A2(n_798),
.B1(n_800),
.B2(n_770),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1193),
.B(n_840),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1180),
.A2(n_805),
.B1(n_807),
.B2(n_801),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1141),
.A2(n_824),
.B1(n_825),
.B2(n_823),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1172),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1206),
.A2(n_1258),
.B1(n_1223),
.B2(n_1179),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1178),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1143),
.A2(n_833),
.B1(n_837),
.B2(n_832),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1178),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1224),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1186),
.A2(n_845),
.B1(n_855),
.B2(n_849),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1193),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1196),
.B(n_1198),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1165),
.A2(n_786),
.B1(n_804),
.B2(n_780),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1192),
.A2(n_862),
.B1(n_863),
.B2(n_861),
.Y(n_1387)
);

XOR2xp5_ASAP7_75t_L g1388 ( 
.A(n_1151),
.B(n_741),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1196),
.B(n_991),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1167),
.A2(n_1189),
.B1(n_1220),
.B2(n_1199),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1198),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1200),
.B(n_991),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1183),
.A2(n_841),
.B1(n_856),
.B2(n_822),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1200),
.B(n_867),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1278),
.B(n_748),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1204),
.A2(n_912),
.B1(n_922),
.B2(n_793),
.Y(n_1396)
);

INVxp33_ASAP7_75t_L g1397 ( 
.A(n_1276),
.Y(n_1397)
);

AOI22x1_ASAP7_75t_SL g1398 ( 
.A1(n_1286),
.A2(n_972),
.B1(n_1047),
.B2(n_958),
.Y(n_1398)
);

AO22x2_ASAP7_75t_L g1399 ( 
.A1(n_1194),
.A2(n_882),
.B1(n_891),
.B2(n_869),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1205),
.Y(n_1400)
);

AO22x2_ASAP7_75t_L g1401 ( 
.A1(n_1234),
.A2(n_898),
.B1(n_908),
.B2(n_896),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1226),
.B(n_725),
.Y(n_1402)
);

OA22x2_ASAP7_75t_L g1403 ( 
.A1(n_1247),
.A2(n_918),
.B1(n_920),
.B2(n_910),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1205),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1201),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1231),
.A2(n_865),
.B1(n_880),
.B2(n_879),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_1234),
.A2(n_928),
.B1(n_941),
.B2(n_927),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1209),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1201),
.B(n_991),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1244),
.B(n_731),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1159),
.A2(n_886),
.B1(n_887),
.B2(n_883),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_SL g1412 ( 
.A(n_1246),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1209),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_895),
.B1(n_915),
.B2(n_914),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1216),
.A2(n_1057),
.B1(n_926),
.B2(n_929),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1240),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1273),
.A2(n_925),
.B1(n_931),
.B2(n_930),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1228),
.A2(n_942),
.B1(n_948),
.B2(n_937),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1211),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1210),
.B(n_645),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1210),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1218),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1282),
.A2(n_950),
.B1(n_953),
.B2(n_952),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1130),
.B(n_645),
.Y(n_1424)
);

AO22x2_ASAP7_75t_L g1425 ( 
.A1(n_1241),
.A2(n_959),
.B1(n_962),
.B2(n_957),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1211),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1233),
.B(n_752),
.Y(n_1427)
);

INVx8_ASAP7_75t_L g1428 ( 
.A(n_1227),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1161),
.A2(n_955),
.B1(n_961),
.B2(n_954),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1130),
.B(n_631),
.Y(n_1430)
);

AO22x2_ASAP7_75t_L g1431 ( 
.A1(n_1241),
.A2(n_969),
.B1(n_981),
.B2(n_963),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1236),
.B(n_755),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1261),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1242),
.A2(n_967),
.B1(n_979),
.B2(n_966),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1124),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_R g1436 ( 
.A1(n_1286),
.A2(n_989),
.B1(n_996),
.B2(n_988),
.Y(n_1436)
);

AO22x2_ASAP7_75t_L g1437 ( 
.A1(n_1242),
.A2(n_1029),
.B1(n_1030),
.B2(n_1006),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1248),
.A2(n_1081),
.B1(n_1091),
.B2(n_1062),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1248),
.A2(n_983),
.B1(n_994),
.B2(n_980),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1260),
.A2(n_997),
.B1(n_1002),
.B2(n_995),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1232),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1162),
.B(n_634),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1162),
.B(n_1173),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1232),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1260),
.A2(n_1008),
.B1(n_1013),
.B2(n_1005),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1169),
.B(n_639),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1169),
.B(n_640),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1262),
.A2(n_1021),
.B1(n_1027),
.B2(n_1016),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1235),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1173),
.B(n_641),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1235),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1262),
.A2(n_1037),
.B1(n_1046),
.B2(n_1034),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_R g1453 ( 
.A1(n_1294),
.A2(n_1117),
.B1(n_1106),
.B2(n_764),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1265),
.A2(n_1066),
.B1(n_1070),
.B2(n_1065),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1251),
.Y(n_1455)
);

AND2x2_ASAP7_75t_SL g1456 ( 
.A(n_1265),
.B(n_759),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1264),
.B(n_767),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1251),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1252),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1294),
.A2(n_1073),
.B1(n_1074),
.B2(n_1071),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1281),
.A2(n_1076),
.B1(n_1079),
.B2(n_1075),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1252),
.Y(n_1462)
);

AO22x2_ASAP7_75t_L g1463 ( 
.A1(n_1281),
.A2(n_773),
.B1(n_777),
.B2(n_771),
.Y(n_1463)
);

AO22x2_ASAP7_75t_L g1464 ( 
.A1(n_1275),
.A2(n_782),
.B1(n_783),
.B2(n_779),
.Y(n_1464)
);

OA22x2_ASAP7_75t_L g1465 ( 
.A1(n_1279),
.A2(n_1095),
.B1(n_1097),
.B2(n_1089),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1227),
.A2(n_1101),
.B1(n_1103),
.B2(n_1100),
.Y(n_1466)
);

AO22x2_ASAP7_75t_L g1467 ( 
.A1(n_1203),
.A2(n_788),
.B1(n_790),
.B2(n_787),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1253),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1182),
.B(n_644),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1253),
.Y(n_1470)
);

BUFx10_ASAP7_75t_L g1471 ( 
.A(n_1203),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1132),
.B(n_1202),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1227),
.A2(n_1110),
.B1(n_1116),
.B2(n_1108),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1182),
.B(n_647),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1237),
.A2(n_655),
.B1(n_664),
.B2(n_649),
.Y(n_1475)
);

AO22x2_ASAP7_75t_L g1476 ( 
.A1(n_1225),
.A2(n_803),
.B1(n_808),
.B2(n_799),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1184),
.B(n_665),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1184),
.B(n_670),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1277),
.A2(n_857),
.B1(n_892),
.B2(n_819),
.Y(n_1479)
);

AOI22x1_ASAP7_75t_L g1480 ( 
.A1(n_1225),
.A2(n_685),
.B1(n_691),
.B2(n_676),
.Y(n_1480)
);

AO22x2_ASAP7_75t_L g1481 ( 
.A1(n_1267),
.A2(n_817),
.B1(n_826),
.B2(n_811),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1188),
.B(n_692),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1267),
.A2(n_853),
.B1(n_907),
.B2(n_834),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1135),
.B(n_911),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1269),
.Y(n_1485)
);

AND2x2_ASAP7_75t_SL g1486 ( 
.A(n_1208),
.B(n_939),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1188),
.B(n_1195),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1156),
.B(n_946),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1269),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1270),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1270),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1284),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1284),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1158),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1125),
.A2(n_701),
.B1(n_703),
.B2(n_697),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1126),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1237),
.A2(n_706),
.B1(n_707),
.B2(n_704),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1134),
.Y(n_1498)
);

AO22x2_ASAP7_75t_L g1499 ( 
.A1(n_1125),
.A2(n_956),
.B1(n_985),
.B2(n_951),
.Y(n_1499)
);

AO22x2_ASAP7_75t_L g1500 ( 
.A1(n_1128),
.A2(n_1007),
.B1(n_1011),
.B2(n_1000),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1128),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1160),
.A2(n_1035),
.B1(n_1042),
.B2(n_1022),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1195),
.B(n_708),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1237),
.A2(n_718),
.B1(n_719),
.B2(n_710),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1140),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1213),
.Y(n_1506)
);

AND2x2_ASAP7_75t_SL g1507 ( 
.A(n_1160),
.B(n_1048),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1213),
.A2(n_1061),
.B1(n_1080),
.B2(n_1050),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1238),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1238),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1249),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1268),
.A2(n_728),
.B1(n_735),
.B2(n_727),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1268),
.A2(n_739),
.B1(n_745),
.B2(n_738),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1249),
.B(n_747),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_SL g1515 ( 
.A(n_1268),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1250),
.A2(n_1102),
.B1(n_1105),
.B2(n_1096),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1250),
.A2(n_756),
.B1(n_765),
.B2(n_749),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1272),
.Y(n_1518)
);

AO22x2_ASAP7_75t_L g1519 ( 
.A1(n_1272),
.A2(n_1109),
.B1(n_58),
.B2(n_55),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1290),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1290),
.A2(n_772),
.B1(n_775),
.B2(n_769),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1256),
.A2(n_781),
.B1(n_784),
.B2(n_778),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1157),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1163),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1163),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1170),
.B(n_789),
.Y(n_1526)
);

AO22x2_ASAP7_75t_L g1527 ( 
.A1(n_1129),
.A2(n_60),
.B1(n_56),
.B2(n_59),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1163),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1136),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1256),
.A2(n_794),
.B1(n_795),
.B2(n_791),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_R g1531 ( 
.A1(n_1168),
.A2(n_63),
.B1(n_56),
.B2(n_60),
.Y(n_1531)
);

CKINVDCx6p67_ASAP7_75t_R g1532 ( 
.A(n_1127),
.Y(n_1532)
);

AO22x2_ASAP7_75t_L g1533 ( 
.A1(n_1129),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1285),
.B(n_796),
.Y(n_1534)
);

INVx5_ASAP7_75t_L g1535 ( 
.A(n_1157),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1163),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1170),
.B(n_797),
.Y(n_1537)
);

AO22x2_ASAP7_75t_L g1538 ( 
.A1(n_1129),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1285),
.A2(n_809),
.B1(n_810),
.B2(n_802),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1163),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1214),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1170),
.B(n_814),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1170),
.B(n_815),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1136),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1257),
.A2(n_818),
.B1(n_821),
.B2(n_816),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1136),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1256),
.A2(n_828),
.B1(n_830),
.B2(n_827),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1136),
.Y(n_1548)
);

AO22x2_ASAP7_75t_L g1549 ( 
.A1(n_1129),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1163),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1230),
.B(n_838),
.Y(n_1551)
);

AO22x2_ASAP7_75t_L g1552 ( 
.A1(n_1129),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1129),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1285),
.A2(n_843),
.B1(n_844),
.B2(n_842),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1163),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1256),
.A2(n_848),
.B1(n_850),
.B2(n_846),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1163),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1285),
.A2(n_871),
.B1(n_877),
.B2(n_851),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1256),
.A2(n_884),
.B1(n_885),
.B2(n_881),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1163),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1285),
.A2(n_890),
.B1(n_894),
.B2(n_888),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1257),
.A2(n_900),
.B1(n_904),
.B2(n_899),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1170),
.B(n_905),
.Y(n_1563)
);

INVxp33_ASAP7_75t_L g1564 ( 
.A(n_1214),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1163),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1256),
.A2(n_917),
.B1(n_919),
.B2(n_916),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1285),
.A2(n_923),
.B1(n_932),
.B2(n_921),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1163),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1157),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1230),
.B(n_1121),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1170),
.B(n_934),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1256),
.A2(n_938),
.B1(n_940),
.B2(n_935),
.Y(n_1572)
);

NAND3x1_ASAP7_75t_L g1573 ( 
.A(n_1146),
.B(n_72),
.C(n_74),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1285),
.B(n_943),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1170),
.B(n_944),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1256),
.A2(n_973),
.B1(n_974),
.B2(n_964),
.Y(n_1576)
);

AO22x2_ASAP7_75t_L g1577 ( 
.A1(n_1129),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1170),
.B(n_976),
.Y(n_1578)
);

BUFx10_ASAP7_75t_L g1579 ( 
.A(n_1157),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1285),
.A2(n_987),
.B1(n_990),
.B2(n_977),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1127),
.B(n_1010),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1285),
.A2(n_993),
.B1(n_998),
.B2(n_992),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1163),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1230),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1254),
.A2(n_1009),
.B1(n_1014),
.B2(n_1003),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1230),
.B(n_1015),
.Y(n_1586)
);

XOR2xp5_ASAP7_75t_L g1587 ( 
.A(n_1256),
.B(n_1017),
.Y(n_1587)
);

AO22x2_ASAP7_75t_L g1588 ( 
.A1(n_1129),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1136),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1256),
.A2(n_1026),
.B1(n_1028),
.B2(n_1019),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1163),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1254),
.A2(n_1038),
.B1(n_1041),
.B2(n_1036),
.Y(n_1592)
);

AOI22x1_ASAP7_75t_SL g1593 ( 
.A1(n_1283),
.A2(n_1044),
.B1(n_1049),
.B2(n_1043),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1136),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1254),
.A2(n_1053),
.B1(n_1054),
.B2(n_1052),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1136),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1256),
.A2(n_1058),
.B1(n_1060),
.B2(n_1056),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1285),
.A2(n_1064),
.B1(n_1067),
.B2(n_1063),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1163),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1136),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1136),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1256),
.A2(n_1078),
.B1(n_1083),
.B2(n_1068),
.Y(n_1602)
);

OAI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1256),
.A2(n_1098),
.B1(n_1099),
.B2(n_1093),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1170),
.B(n_1104),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1157),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1163),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1285),
.A2(n_1111),
.B1(n_1112),
.B2(n_1107),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1163),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1256),
.A2(n_1118),
.B1(n_1119),
.B2(n_1115),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1285),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_R g1611 ( 
.A1(n_1168),
.A2(n_83),
.B1(n_79),
.B2(n_82),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1170),
.B(n_285),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1163),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1163),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1157),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1136),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1256),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1254),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1170),
.B(n_292),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1256),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1129),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_R g1622 ( 
.A1(n_1168),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1230),
.B(n_93),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1170),
.B(n_296),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1170),
.B(n_297),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1163),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1285),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1256),
.A2(n_100),
.B1(n_97),
.B2(n_99),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1400),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1385),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1360),
.B(n_100),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1320),
.Y(n_1632)
);

AND2x6_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_303),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1365),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1507),
.B(n_304),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1408),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1501),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1344),
.B(n_101),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1494),
.Y(n_1639)
);

AND2x6_ASAP7_75t_L g1640 ( 
.A(n_1619),
.B(n_305),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1332),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1421),
.B(n_306),
.Y(n_1642)
);

XOR2x2_ASAP7_75t_L g1643 ( 
.A(n_1299),
.B(n_102),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1413),
.Y(n_1644)
);

INVxp33_ASAP7_75t_SL g1645 ( 
.A(n_1587),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1349),
.B(n_103),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1419),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1451),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1496),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1458),
.Y(n_1650)
);

XOR2xp5_ASAP7_75t_L g1651 ( 
.A(n_1388),
.B(n_307),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1498),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1300),
.B(n_104),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1505),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1584),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1374),
.B(n_309),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1422),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1389),
.B(n_311),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1314),
.Y(n_1659)
);

INVxp33_ASAP7_75t_SL g1660 ( 
.A(n_1530),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1404),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1433),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1459),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1462),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1470),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1435),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1485),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1489),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1426),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1441),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1335),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1296),
.B(n_106),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1444),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1551),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1570),
.B(n_1586),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1449),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1347),
.B(n_107),
.Y(n_1677)
);

XOR2xp5_ASAP7_75t_L g1678 ( 
.A(n_1315),
.B(n_312),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1455),
.Y(n_1679)
);

CKINVDCx16_ASAP7_75t_R g1680 ( 
.A(n_1309),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1468),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1472),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1306),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1298),
.B(n_107),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1420),
.B(n_108),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1490),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1532),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1492),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1493),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1310),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1313),
.B(n_108),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1317),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1579),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1354),
.B(n_317),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1305),
.B(n_109),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1319),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1337),
.B(n_109),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1323),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1345),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1329),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1350),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1404),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1318),
.B(n_110),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1351),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1392),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1491),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1302),
.B(n_114),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1491),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1427),
.B(n_114),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1355),
.Y(n_1710)
);

AOI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1379),
.A2(n_320),
.B(n_318),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1368),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1432),
.B(n_115),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1307),
.B(n_115),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1361),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1354),
.B(n_1486),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1304),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1471),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1308),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1522),
.B(n_116),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1297),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1301),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1535),
.B(n_627),
.Y(n_1723)
);

INVxp33_ASAP7_75t_L g1724 ( 
.A(n_1564),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1295),
.B(n_116),
.Y(n_1725)
);

XOR2xp5_ASAP7_75t_L g1726 ( 
.A(n_1397),
.B(n_322),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1303),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1324),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1342),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1343),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1535),
.B(n_1334),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1377),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1371),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1581),
.B(n_117),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1327),
.Y(n_1735)
);

NAND2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1336),
.B(n_325),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1556),
.B(n_117),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1409),
.B(n_329),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1524),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1529),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1525),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1509),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1544),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1593),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1546),
.Y(n_1745)
);

NOR2xp67_ASAP7_75t_L g1746 ( 
.A(n_1523),
.B(n_332),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1548),
.Y(n_1747)
);

INVx4_ASAP7_75t_L g1748 ( 
.A(n_1509),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1589),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1594),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1596),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1348),
.B(n_118),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1600),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1601),
.Y(n_1754)
);

INVxp33_ASAP7_75t_L g1755 ( 
.A(n_1359),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1526),
.B(n_1537),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1616),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1528),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1536),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1540),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1550),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1555),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1547),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1557),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1560),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1565),
.Y(n_1766)
);

XOR2xp5_ASAP7_75t_L g1767 ( 
.A(n_1312),
.B(n_339),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1390),
.A2(n_342),
.B(n_340),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1322),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1354),
.B(n_343),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1568),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1511),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1402),
.B(n_347),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1583),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1591),
.Y(n_1775)
);

XNOR2xp5_ASAP7_75t_L g1776 ( 
.A(n_1396),
.B(n_118),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1599),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1606),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1572),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_SL g1780 ( 
.A(n_1416),
.B(n_119),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1541),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1456),
.B(n_348),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1430),
.B(n_1442),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1608),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1613),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1614),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1328),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1585),
.B(n_119),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1626),
.Y(n_1789)
);

XNOR2xp5_ASAP7_75t_L g1790 ( 
.A(n_1369),
.B(n_120),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1384),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1353),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1381),
.Y(n_1793)
);

XOR2xp5_ASAP7_75t_L g1794 ( 
.A(n_1398),
.B(n_350),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1391),
.Y(n_1795)
);

INVx8_ASAP7_75t_L g1796 ( 
.A(n_1581),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1559),
.B(n_120),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1405),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1446),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1506),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1602),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1624),
.A2(n_355),
.B(n_352),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1542),
.B(n_124),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1566),
.B(n_1576),
.Y(n_1804)
);

XNOR2xp5_ASAP7_75t_L g1805 ( 
.A(n_1378),
.B(n_124),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1327),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1367),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1367),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1543),
.B(n_1563),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1403),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1394),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1358),
.Y(n_1812)
);

XNOR2xp5_ASAP7_75t_L g1813 ( 
.A(n_1375),
.B(n_125),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1394),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1590),
.B(n_127),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1539),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1390),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1495),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1518),
.Y(n_1819)
);

XNOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1415),
.B(n_127),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1410),
.B(n_356),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1331),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1554),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1464),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1443),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1464),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1625),
.A2(n_361),
.B(n_360),
.Y(n_1827)
);

XOR2x2_ASAP7_75t_L g1828 ( 
.A(n_1573),
.B(n_1418),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1395),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1597),
.B(n_128),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1571),
.B(n_128),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1484),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1575),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1484),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1447),
.B(n_363),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1487),
.Y(n_1836)
);

XNOR2xp5_ASAP7_75t_L g1837 ( 
.A(n_1527),
.B(n_130),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1488),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1450),
.B(n_364),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1488),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1578),
.B(n_132),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1558),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1457),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1520),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1457),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1604),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1561),
.Y(n_1847)
);

INVxp33_ASAP7_75t_L g1848 ( 
.A(n_1372),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1603),
.B(n_132),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1469),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1510),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1474),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1477),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1478),
.Y(n_1854)
);

XNOR2xp5_ASAP7_75t_L g1855 ( 
.A(n_1527),
.B(n_1533),
.Y(n_1855)
);

OR2x6_ASAP7_75t_L g1856 ( 
.A(n_1533),
.B(n_1538),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1482),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1503),
.B(n_366),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1514),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1499),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1499),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1609),
.B(n_135),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1500),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1500),
.Y(n_1864)
);

XOR2xp5_ASAP7_75t_L g1865 ( 
.A(n_1465),
.B(n_368),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1338),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1569),
.B(n_135),
.Y(n_1867)
);

XNOR2xp5_ASAP7_75t_L g1868 ( 
.A(n_1538),
.B(n_136),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1467),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1467),
.Y(n_1870)
);

INVx4_ASAP7_75t_SL g1871 ( 
.A(n_1515),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1567),
.B(n_136),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1580),
.B(n_137),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1582),
.Y(n_1874)
);

NAND2xp33_ASAP7_75t_R g1875 ( 
.A(n_1623),
.B(n_137),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1476),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1476),
.Y(n_1877)
);

CKINVDCx20_ASAP7_75t_R g1878 ( 
.A(n_1598),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1481),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1534),
.B(n_369),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1481),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1386),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1424),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1605),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1386),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1339),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1339),
.Y(n_1887)
);

INVxp67_ASAP7_75t_SL g1888 ( 
.A(n_1574),
.Y(n_1888)
);

AND2x2_ASAP7_75t_SL g1889 ( 
.A(n_1610),
.B(n_139),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1615),
.B(n_139),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1321),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1592),
.B(n_1595),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1401),
.Y(n_1893)
);

INVxp33_ASAP7_75t_L g1894 ( 
.A(n_1373),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1434),
.B(n_141),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1401),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1407),
.Y(n_1897)
);

CKINVDCx16_ASAP7_75t_R g1898 ( 
.A(n_1412),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1407),
.Y(n_1899)
);

NAND2xp33_ASAP7_75t_SL g1900 ( 
.A(n_1483),
.B(n_1620),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1439),
.B(n_142),
.Y(n_1901)
);

INVx4_ASAP7_75t_SL g1902 ( 
.A(n_1628),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1425),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1364),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1425),
.Y(n_1905)
);

INVxp67_ASAP7_75t_SL g1906 ( 
.A(n_1480),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1431),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1431),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1437),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1437),
.Y(n_1910)
);

XNOR2x2_ASAP7_75t_L g1911 ( 
.A(n_1549),
.B(n_143),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1607),
.B(n_143),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1438),
.Y(n_1913)
);

XNOR2x2_ASAP7_75t_L g1914 ( 
.A(n_1549),
.B(n_145),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1406),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1445),
.B(n_145),
.Y(n_1916)
);

OR2x6_ASAP7_75t_L g1917 ( 
.A(n_1552),
.B(n_146),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1438),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1393),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1356),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1452),
.B(n_146),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1330),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1393),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1466),
.B(n_370),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1356),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1399),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1414),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1454),
.B(n_147),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1399),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1545),
.B(n_147),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1502),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1340),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1370),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_SL g1934 ( 
.A(n_1382),
.B(n_149),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1340),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1463),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1473),
.B(n_371),
.Y(n_1937)
);

XOR2xp5_ASAP7_75t_L g1938 ( 
.A(n_1362),
.B(n_375),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1475),
.B(n_376),
.Y(n_1939)
);

OAI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1497),
.A2(n_384),
.B(n_380),
.Y(n_1940)
);

CKINVDCx20_ASAP7_75t_R g1941 ( 
.A(n_1417),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1428),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1330),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1562),
.B(n_149),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1504),
.A2(n_387),
.B(n_385),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1463),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_SL g1947 ( 
.A(n_1341),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1321),
.Y(n_1948)
);

AND2x6_ASAP7_75t_L g1949 ( 
.A(n_1512),
.B(n_390),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1423),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1627),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1674),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1787),
.B(n_1440),
.Y(n_1953)
);

AND2x2_ASAP7_75t_SL g1954 ( 
.A(n_1889),
.B(n_1448),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1717),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1724),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1742),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1655),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1675),
.B(n_1326),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1906),
.A2(n_1513),
.B(n_1461),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1719),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1810),
.B(n_1517),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1833),
.B(n_1341),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1716),
.A2(n_1383),
.B(n_1366),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1656),
.B(n_1428),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1798),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1661),
.Y(n_1967)
);

AND2x2_ASAP7_75t_SL g1968 ( 
.A(n_1680),
.B(n_1552),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1656),
.B(n_1387),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1739),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1658),
.B(n_1521),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1741),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1661),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1658),
.B(n_1376),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1661),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1630),
.Y(n_1976)
);

INVx8_ASAP7_75t_L g1977 ( 
.A(n_1796),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1702),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1781),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1777),
.Y(n_1980)
);

INVxp67_ASAP7_75t_L g1981 ( 
.A(n_1683),
.Y(n_1981)
);

NOR2xp67_ASAP7_75t_L g1982 ( 
.A(n_1942),
.B(n_391),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1671),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1642),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1769),
.B(n_1733),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1942),
.B(n_1380),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1793),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1756),
.B(n_1809),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1634),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1738),
.B(n_1411),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1699),
.B(n_1553),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1715),
.B(n_1553),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1875),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1807),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1705),
.B(n_1577),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1884),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1738),
.B(n_1429),
.Y(n_1997)
);

BUFx5_ASAP7_75t_L g1998 ( 
.A(n_1633),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1822),
.B(n_1577),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1758),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1702),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1759),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1760),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1942),
.B(n_1588),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1631),
.B(n_1357),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1649),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1652),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1702),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1867),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1682),
.B(n_1352),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1783),
.B(n_1519),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1848),
.B(n_1363),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1761),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1706),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1637),
.B(n_1519),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1654),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1646),
.B(n_1618),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1762),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1764),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1817),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1639),
.B(n_1460),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1850),
.B(n_1508),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1846),
.B(n_1588),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1859),
.B(n_1516),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1642),
.B(n_1666),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1890),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1765),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1766),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1852),
.B(n_1479),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1706),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1771),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1657),
.B(n_393),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1697),
.B(n_1621),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1853),
.B(n_1346),
.Y(n_2034)
);

BUFx5_ASAP7_75t_L g2035 ( 
.A(n_1633),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1774),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1706),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1775),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1854),
.B(n_1311),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1694),
.A2(n_397),
.B(n_394),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1662),
.B(n_400),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1857),
.B(n_1621),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1695),
.B(n_1316),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1714),
.B(n_1333),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1703),
.B(n_1325),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1888),
.B(n_1617),
.Y(n_2046)
);

AND2x6_ASAP7_75t_L g2047 ( 
.A(n_1937),
.B(n_1531),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1778),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1784),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1785),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1786),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1883),
.B(n_150),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1789),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1629),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1799),
.B(n_150),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1636),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1644),
.Y(n_2057)
);

INVxp67_ASAP7_75t_SL g2058 ( 
.A(n_1708),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1894),
.B(n_151),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1708),
.Y(n_2060)
);

AND2x2_ASAP7_75t_SL g2061 ( 
.A(n_1691),
.B(n_1611),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1647),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1948),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_1708),
.Y(n_2064)
);

INVxp33_ASAP7_75t_L g2065 ( 
.A(n_1638),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_1693),
.Y(n_2066)
);

INVxp33_ASAP7_75t_L g2067 ( 
.A(n_1684),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1773),
.B(n_402),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1718),
.B(n_151),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1735),
.Y(n_2070)
);

OAI21xp33_ASAP7_75t_L g2071 ( 
.A1(n_1709),
.A2(n_1713),
.B(n_1916),
.Y(n_2071)
);

AND2x2_ASAP7_75t_SL g2072 ( 
.A(n_1720),
.B(n_1622),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1829),
.B(n_153),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1819),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1648),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1650),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1866),
.B(n_154),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1665),
.Y(n_2078)
);

NAND2x1p5_ASAP7_75t_L g2079 ( 
.A(n_1843),
.B(n_1773),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1663),
.Y(n_2080)
);

INVxp33_ASAP7_75t_L g2081 ( 
.A(n_1837),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1821),
.B(n_403),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1653),
.B(n_154),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1856),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1821),
.B(n_405),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1664),
.Y(n_2086)
);

AND2x6_ASAP7_75t_L g2087 ( 
.A(n_1937),
.B(n_1453),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1755),
.B(n_155),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1667),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1735),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1931),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1635),
.B(n_406),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_1851),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1782),
.B(n_1707),
.Y(n_2094)
);

OAI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1770),
.A2(n_1436),
.B(n_412),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1856),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1672),
.B(n_407),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1904),
.B(n_157),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1825),
.B(n_157),
.Y(n_2099)
);

INVx4_ASAP7_75t_L g2100 ( 
.A(n_1735),
.Y(n_2100)
);

OR2x2_ASAP7_75t_SL g2101 ( 
.A(n_1951),
.B(n_158),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1752),
.B(n_414),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1668),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1690),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1692),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1836),
.B(n_420),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1844),
.B(n_421),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1696),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1891),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1698),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1933),
.B(n_1804),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1871),
.B(n_158),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_1843),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1803),
.B(n_423),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1871),
.B(n_159),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1895),
.B(n_159),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1808),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1808),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1901),
.B(n_160),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1700),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1917),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1701),
.Y(n_2122)
);

AND2x2_ASAP7_75t_SL g2123 ( 
.A(n_1737),
.B(n_160),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1843),
.B(n_1731),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1704),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1710),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1831),
.B(n_161),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1886),
.B(n_424),
.Y(n_2128)
);

NOR2xp67_ASAP7_75t_L g2129 ( 
.A(n_1748),
.B(n_626),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1712),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1887),
.B(n_426),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1669),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1841),
.B(n_161),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1918),
.B(n_162),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1824),
.B(n_429),
.Y(n_2135)
);

INVxp67_ASAP7_75t_L g2136 ( 
.A(n_1921),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1818),
.B(n_162),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1670),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1685),
.B(n_163),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1892),
.A2(n_441),
.B1(n_442),
.B2(n_437),
.Y(n_2140)
);

BUFx4f_ASAP7_75t_L g2141 ( 
.A(n_1949),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1673),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1882),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1920),
.B(n_1925),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1725),
.B(n_163),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1676),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1808),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_1826),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1893),
.B(n_164),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1679),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1681),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1885),
.Y(n_2152)
);

INVx2_ASAP7_75t_SL g2153 ( 
.A(n_1845),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1686),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1896),
.B(n_164),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1897),
.B(n_168),
.Y(n_2156)
);

INVx4_ASAP7_75t_L g2157 ( 
.A(n_1748),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1772),
.B(n_444),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1688),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1899),
.B(n_1903),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1802),
.A2(n_449),
.B(n_447),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1689),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1806),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1721),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1827),
.B(n_450),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1811),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_1722),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1633),
.B(n_452),
.Y(n_2168)
);

AND2x2_ASAP7_75t_SL g2169 ( 
.A(n_1797),
.B(n_169),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1727),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1832),
.B(n_455),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1905),
.B(n_170),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1860),
.A2(n_459),
.B(n_458),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_1928),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_1861),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1907),
.B(n_171),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1633),
.B(n_460),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1908),
.B(n_1909),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1728),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1729),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1730),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1732),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1740),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_1863),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1640),
.B(n_462),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1743),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_1864),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1745),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1640),
.B(n_464),
.Y(n_2189)
);

AND2x6_ASAP7_75t_L g2190 ( 
.A(n_1936),
.B(n_465),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1640),
.B(n_466),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1747),
.Y(n_2192)
);

BUFx2_ASAP7_75t_L g2193 ( 
.A(n_1917),
.Y(n_2193)
);

INVx4_ASAP7_75t_L g2194 ( 
.A(n_1640),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1749),
.Y(n_2195)
);

INVx4_ASAP7_75t_L g2196 ( 
.A(n_1800),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1987),
.Y(n_2197)
);

OR2x6_ASAP7_75t_L g2198 ( 
.A(n_1977),
.B(n_1796),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_1956),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2063),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_1979),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2143),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1984),
.B(n_1869),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2179),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1988),
.B(n_1910),
.Y(n_2205)
);

CKINVDCx20_ASAP7_75t_R g2206 ( 
.A(n_1958),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1984),
.B(n_1870),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1957),
.B(n_1814),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2111),
.B(n_1632),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2071),
.B(n_1876),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_1993),
.B(n_1932),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_1975),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_1998),
.B(n_1949),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2067),
.B(n_1641),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1955),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2025),
.B(n_1877),
.Y(n_2216)
);

INVx5_ASAP7_75t_L g2217 ( 
.A(n_1977),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1966),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1985),
.B(n_1913),
.Y(n_2219)
);

NAND2xp33_ASAP7_75t_L g2220 ( 
.A(n_1998),
.B(n_1949),
.Y(n_2220)
);

INVxp67_ASAP7_75t_SL g2221 ( 
.A(n_1975),
.Y(n_2221)
);

INVxp67_ASAP7_75t_SL g2222 ( 
.A(n_1975),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2179),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2136),
.B(n_1935),
.Y(n_2224)
);

NOR2x1_ASAP7_75t_L g2225 ( 
.A(n_2157),
.B(n_1939),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2181),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2094),
.B(n_1881),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_1996),
.B(n_1919),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2181),
.Y(n_2229)
);

BUFx2_ASAP7_75t_L g2230 ( 
.A(n_2109),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2186),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1978),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2186),
.Y(n_2233)
);

BUFx4f_ASAP7_75t_L g2234 ( 
.A(n_2079),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2093),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1959),
.B(n_2017),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1953),
.B(n_1923),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1978),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_1967),
.Y(n_2239)
);

NAND2x1p5_ASAP7_75t_L g2240 ( 
.A(n_2157),
.B(n_1791),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1978),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_2166),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1983),
.B(n_1926),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_2152),
.Y(n_2244)
);

BUFx2_ASAP7_75t_L g2245 ( 
.A(n_2084),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2174),
.B(n_1929),
.Y(n_2246)
);

INVx5_ASAP7_75t_L g2247 ( 
.A(n_2008),
.Y(n_2247)
);

CKINVDCx6p67_ASAP7_75t_R g2248 ( 
.A(n_2066),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1973),
.Y(n_2249)
);

BUFx12f_ASAP7_75t_L g2250 ( 
.A(n_2121),
.Y(n_2250)
);

BUFx4f_ASAP7_75t_L g2251 ( 
.A(n_2128),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2031),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2124),
.B(n_1834),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1981),
.B(n_1872),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1969),
.B(n_1879),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2065),
.B(n_1873),
.Y(n_2256)
);

OR2x6_ASAP7_75t_L g2257 ( 
.A(n_2004),
.B(n_1734),
.Y(n_2257)
);

AND2x2_ASAP7_75t_SL g2258 ( 
.A(n_2123),
.B(n_1815),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_2153),
.B(n_1838),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1989),
.B(n_1946),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_2008),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_2113),
.B(n_2171),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2008),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1960),
.B(n_1912),
.Y(n_2264)
);

INVx4_ASAP7_75t_L g2265 ( 
.A(n_2014),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2031),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1961),
.Y(n_2267)
);

NAND2x1_ASAP7_75t_L g2268 ( 
.A(n_2194),
.B(n_1750),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2175),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2096),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2171),
.B(n_2144),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2095),
.B(n_1971),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2127),
.B(n_1930),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2036),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2133),
.B(n_1944),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2077),
.B(n_2044),
.Y(n_2276)
);

INVxp67_ASAP7_75t_L g2277 ( 
.A(n_2088),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2043),
.B(n_1840),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_1976),
.B(n_1943),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1952),
.B(n_1830),
.Y(n_2280)
);

NAND2x1p5_ASAP7_75t_L g2281 ( 
.A(n_2060),
.B(n_1751),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2036),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2001),
.B(n_1753),
.Y(n_2283)
);

BUFx2_ASAP7_75t_SL g2284 ( 
.A(n_1982),
.Y(n_2284)
);

BUFx4f_ASAP7_75t_L g2285 ( 
.A(n_2128),
.Y(n_2285)
);

BUFx5_ASAP7_75t_L g2286 ( 
.A(n_2190),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_2014),
.Y(n_2287)
);

BUFx8_ASAP7_75t_SL g2288 ( 
.A(n_2193),
.Y(n_2288)
);

INVxp67_ASAP7_75t_L g2289 ( 
.A(n_2098),
.Y(n_2289)
);

AND2x6_ASAP7_75t_L g2290 ( 
.A(n_2140),
.B(n_1849),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2009),
.B(n_1880),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2037),
.B(n_1754),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2090),
.B(n_1757),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2026),
.B(n_2091),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1964),
.B(n_1862),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2038),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2083),
.B(n_1924),
.Y(n_2297)
);

BUFx12f_ASAP7_75t_L g2298 ( 
.A(n_2101),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2038),
.Y(n_2299)
);

BUFx4f_ASAP7_75t_L g2300 ( 
.A(n_2131),
.Y(n_2300)
);

AND2x2_ASAP7_75t_SL g2301 ( 
.A(n_2169),
.B(n_1677),
.Y(n_2301)
);

BUFx12f_ASAP7_75t_L g2302 ( 
.A(n_2112),
.Y(n_2302)
);

INVx4_ASAP7_75t_L g2303 ( 
.A(n_2014),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_SL g2304 ( 
.A(n_2012),
.B(n_1687),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2048),
.Y(n_2305)
);

BUFx8_ASAP7_75t_L g2306 ( 
.A(n_1963),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_2030),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_2118),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_2055),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2048),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2160),
.B(n_1788),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2059),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1970),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2011),
.B(n_1940),
.Y(n_2314)
);

NAND2x1p5_ASAP7_75t_L g2315 ( 
.A(n_2060),
.B(n_1792),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2178),
.B(n_1855),
.Y(n_2316)
);

NOR2x1_ASAP7_75t_SL g2317 ( 
.A(n_2194),
.B(n_1835),
.Y(n_2317)
);

OR2x6_ASAP7_75t_L g2318 ( 
.A(n_2131),
.B(n_1734),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_2020),
.Y(n_2319)
);

BUFx3_ASAP7_75t_L g2320 ( 
.A(n_2030),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2030),
.Y(n_2321)
);

INVx4_ASAP7_75t_L g2322 ( 
.A(n_2070),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_1962),
.Y(n_2323)
);

AND2x6_ASAP7_75t_L g2324 ( 
.A(n_2033),
.B(n_1839),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2116),
.B(n_1945),
.Y(n_2325)
);

INVx4_ASAP7_75t_L g2326 ( 
.A(n_2070),
.Y(n_2326)
);

INVx8_ASAP7_75t_L g2327 ( 
.A(n_2070),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2142),
.B(n_1795),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2045),
.B(n_1911),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1972),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2148),
.Y(n_2331)
);

BUFx12f_ASAP7_75t_L g2332 ( 
.A(n_2115),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2089),
.Y(n_2333)
);

INVx11_ASAP7_75t_L g2334 ( 
.A(n_2087),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_2117),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2119),
.B(n_1801),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2089),
.Y(n_2337)
);

OR2x6_ASAP7_75t_L g2338 ( 
.A(n_2046),
.B(n_1768),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2151),
.B(n_1858),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2039),
.B(n_1914),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2042),
.B(n_1898),
.Y(n_2341)
);

INVx4_ASAP7_75t_L g2342 ( 
.A(n_2117),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2184),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2010),
.B(n_1767),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2061),
.B(n_1659),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2134),
.B(n_1678),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2151),
.B(n_1949),
.Y(n_2347)
);

AND2x6_ASAP7_75t_L g2348 ( 
.A(n_2168),
.B(n_1660),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_1962),
.Y(n_2349)
);

AND2x2_ASAP7_75t_SL g2350 ( 
.A(n_1954),
.B(n_1780),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2117),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_2087),
.Y(n_2352)
);

BUFx3_ASAP7_75t_L g2353 ( 
.A(n_2147),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2201),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_2218),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2230),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2204),
.Y(n_2357)
);

INVx2_ASAP7_75t_SL g2358 ( 
.A(n_2235),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2277),
.B(n_1812),
.Y(n_2359)
);

INVx2_ASAP7_75t_SL g2360 ( 
.A(n_2253),
.Y(n_2360)
);

INVx4_ASAP7_75t_L g2361 ( 
.A(n_2327),
.Y(n_2361)
);

BUFx3_ASAP7_75t_L g2362 ( 
.A(n_2217),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2212),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2248),
.Y(n_2364)
);

INVx5_ASAP7_75t_L g2365 ( 
.A(n_2198),
.Y(n_2365)
);

NAND2x1p5_ASAP7_75t_L g2366 ( 
.A(n_2247),
.B(n_2217),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2223),
.Y(n_2367)
);

INVxp67_ASAP7_75t_SL g2368 ( 
.A(n_2212),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_2232),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2199),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_2323),
.Y(n_2371)
);

OR2x6_ASAP7_75t_L g2372 ( 
.A(n_2198),
.B(n_2032),
.Y(n_2372)
);

BUFx2_ASAP7_75t_L g2373 ( 
.A(n_2245),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2226),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2252),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2276),
.B(n_2137),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2229),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_2206),
.Y(n_2378)
);

BUFx3_ASAP7_75t_L g2379 ( 
.A(n_2242),
.Y(n_2379)
);

BUFx3_ASAP7_75t_L g2380 ( 
.A(n_2270),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2256),
.B(n_2072),
.Y(n_2381)
);

INVx4_ASAP7_75t_L g2382 ( 
.A(n_2327),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_2349),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_2247),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2232),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2238),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2266),
.Y(n_2387)
);

INVxp67_ASAP7_75t_SL g2388 ( 
.A(n_2238),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_2241),
.Y(n_2389)
);

INVx3_ASAP7_75t_SL g2390 ( 
.A(n_2341),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_2329),
.B(n_2015),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2279),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2274),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_2250),
.Y(n_2394)
);

BUFx6f_ASAP7_75t_L g2395 ( 
.A(n_2241),
.Y(n_2395)
);

BUFx3_ASAP7_75t_L g2396 ( 
.A(n_2208),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2282),
.Y(n_2397)
);

BUFx12f_ASAP7_75t_L g2398 ( 
.A(n_2306),
.Y(n_2398)
);

BUFx3_ASAP7_75t_L g2399 ( 
.A(n_2302),
.Y(n_2399)
);

BUFx12f_ASAP7_75t_L g2400 ( 
.A(n_2332),
.Y(n_2400)
);

BUFx2_ASAP7_75t_SL g2401 ( 
.A(n_2286),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2259),
.Y(n_2402)
);

INVx1_ASAP7_75t_SL g2403 ( 
.A(n_2228),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2331),
.Y(n_2404)
);

INVx3_ASAP7_75t_SL g2405 ( 
.A(n_2257),
.Y(n_2405)
);

BUFx12f_ASAP7_75t_L g2406 ( 
.A(n_2257),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_2261),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2264),
.B(n_2141),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2236),
.B(n_2139),
.Y(n_2409)
);

BUFx2_ASAP7_75t_R g2410 ( 
.A(n_2288),
.Y(n_2410)
);

OR2x6_ASAP7_75t_L g2411 ( 
.A(n_2318),
.B(n_2032),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2261),
.Y(n_2412)
);

INVxp67_ASAP7_75t_SL g2413 ( 
.A(n_2263),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2296),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2312),
.B(n_1645),
.Y(n_2415)
);

BUFx4_ASAP7_75t_SL g2416 ( 
.A(n_2318),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2200),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2231),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2336),
.B(n_2023),
.Y(n_2419)
);

BUFx6f_ASAP7_75t_L g2420 ( 
.A(n_2263),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2295),
.B(n_2005),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2243),
.Y(n_2422)
);

INVx4_ASAP7_75t_L g2423 ( 
.A(n_2287),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2271),
.Y(n_2424)
);

INVx3_ASAP7_75t_SL g2425 ( 
.A(n_2352),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_2244),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_2214),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2299),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_2269),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2211),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2233),
.Y(n_2431)
);

BUFx3_ASAP7_75t_L g2432 ( 
.A(n_2202),
.Y(n_2432)
);

NAND2x1p5_ASAP7_75t_L g2433 ( 
.A(n_2265),
.B(n_2064),
.Y(n_2433)
);

BUFx4f_ASAP7_75t_L g2434 ( 
.A(n_2348),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2305),
.Y(n_2435)
);

BUFx12f_ASAP7_75t_L g2436 ( 
.A(n_2298),
.Y(n_2436)
);

BUFx5_ASAP7_75t_L g2437 ( 
.A(n_2310),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2319),
.Y(n_2438)
);

INVxp67_ASAP7_75t_SL g2439 ( 
.A(n_2287),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2262),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2307),
.Y(n_2441)
);

NAND2x1p5_ASAP7_75t_L g2442 ( 
.A(n_2303),
.B(n_2064),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_SL g2443 ( 
.A(n_2348),
.Y(n_2443)
);

INVx3_ASAP7_75t_SL g2444 ( 
.A(n_2278),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2351),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2254),
.B(n_1995),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_SL g2447 ( 
.A(n_2348),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2325),
.B(n_2187),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2333),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2307),
.Y(n_2450)
);

BUFx2_ASAP7_75t_SL g2451 ( 
.A(n_2286),
.Y(n_2451)
);

NAND2x1p5_ASAP7_75t_L g2452 ( 
.A(n_2322),
.B(n_2100),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2367),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2376),
.B(n_2346),
.Y(n_2454)
);

INVx6_ASAP7_75t_L g2455 ( 
.A(n_2365),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_SL g2456 ( 
.A1(n_2381),
.A2(n_2301),
.B1(n_2258),
.B2(n_2350),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2409),
.A2(n_2325),
.B1(n_2251),
.B2(n_2300),
.Y(n_2457)
);

OAI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2448),
.A2(n_2285),
.B1(n_2273),
.B2(n_2275),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2367),
.Y(n_2459)
);

INVx1_ASAP7_75t_SL g2460 ( 
.A(n_2356),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2419),
.A2(n_2290),
.B1(n_2087),
.B2(n_2047),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2377),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2446),
.B(n_2346),
.Y(n_2463)
);

CKINVDCx11_ASAP7_75t_R g2464 ( 
.A(n_2398),
.Y(n_2464)
);

INVx6_ASAP7_75t_L g2465 ( 
.A(n_2365),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2403),
.B(n_2316),
.Y(n_2466)
);

OAI22xp33_ASAP7_75t_SL g2467 ( 
.A1(n_2444),
.A2(n_1934),
.B1(n_2272),
.B2(n_2289),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_SL g2468 ( 
.A1(n_2359),
.A2(n_2209),
.B1(n_2087),
.B2(n_2304),
.Y(n_2468)
);

CKINVDCx11_ASAP7_75t_R g2469 ( 
.A(n_2400),
.Y(n_2469)
);

CKINVDCx11_ASAP7_75t_R g2470 ( 
.A(n_2436),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2391),
.B(n_2316),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_SL g2472 ( 
.A(n_2362),
.Y(n_2472)
);

BUFx8_ASAP7_75t_L g2473 ( 
.A(n_2443),
.Y(n_2473)
);

INVx8_ASAP7_75t_L g2474 ( 
.A(n_2365),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_SL g2475 ( 
.A1(n_2415),
.A2(n_1779),
.B1(n_1763),
.B2(n_1790),
.Y(n_2475)
);

BUFx2_ASAP7_75t_L g2476 ( 
.A(n_2356),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2377),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2418),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_SL g2479 ( 
.A1(n_2427),
.A2(n_2280),
.B1(n_2290),
.B2(n_2047),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2421),
.A2(n_2297),
.B1(n_2314),
.B2(n_2141),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2418),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2357),
.Y(n_2482)
);

OAI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2408),
.A2(n_2161),
.B(n_2165),
.Y(n_2483)
);

BUFx3_ASAP7_75t_L g2484 ( 
.A(n_2380),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2410),
.Y(n_2485)
);

OAI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2390),
.A2(n_2344),
.B1(n_2340),
.B2(n_2309),
.Y(n_2486)
);

CKINVDCx11_ASAP7_75t_R g2487 ( 
.A(n_2405),
.Y(n_2487)
);

CKINVDCx20_ASAP7_75t_R g2488 ( 
.A(n_2378),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2422),
.B(n_2237),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2440),
.A2(n_2345),
.B1(n_1823),
.B2(n_1842),
.Y(n_2490)
);

INVx8_ASAP7_75t_L g2491 ( 
.A(n_2363),
.Y(n_2491)
);

AOI22xp33_ASAP7_75t_L g2492 ( 
.A1(n_2383),
.A2(n_2290),
.B1(n_2047),
.B2(n_2145),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2375),
.Y(n_2493)
);

INVx4_ASAP7_75t_L g2494 ( 
.A(n_2361),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2374),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2431),
.Y(n_2496)
);

AOI22xp33_ASAP7_75t_L g2497 ( 
.A1(n_2383),
.A2(n_2047),
.B1(n_1828),
.B2(n_1968),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2411),
.A2(n_2220),
.B(n_2213),
.Y(n_2498)
);

BUFx4_ASAP7_75t_SL g2499 ( 
.A(n_2399),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2430),
.B(n_2227),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2449),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2424),
.A2(n_1847),
.B1(n_1874),
.B2(n_1816),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_SL g2503 ( 
.A1(n_2427),
.A2(n_1878),
.B1(n_1927),
.B2(n_1915),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2387),
.Y(n_2504)
);

INVx4_ASAP7_75t_L g2505 ( 
.A(n_2384),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2373),
.Y(n_2506)
);

OAI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2364),
.A2(n_2294),
.B1(n_1990),
.B2(n_1997),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2393),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2363),
.Y(n_2509)
);

AOI22xp33_ASAP7_75t_SL g2510 ( 
.A1(n_2371),
.A2(n_1950),
.B1(n_1941),
.B2(n_2190),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_2371),
.A2(n_1900),
.B1(n_2324),
.B2(n_2311),
.Y(n_2511)
);

CKINVDCx11_ASAP7_75t_R g2512 ( 
.A(n_2406),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2397),
.A2(n_1965),
.B1(n_2255),
.B2(n_2347),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2414),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2428),
.Y(n_2515)
);

INVx6_ASAP7_75t_L g2516 ( 
.A(n_2361),
.Y(n_2516)
);

OAI21xp5_ASAP7_75t_L g2517 ( 
.A1(n_2435),
.A2(n_2097),
.B(n_2338),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2358),
.B(n_2205),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_L g2519 ( 
.A1(n_2424),
.A2(n_2324),
.B1(n_2311),
.B2(n_1776),
.Y(n_2519)
);

INVx2_ASAP7_75t_SL g2520 ( 
.A(n_2379),
.Y(n_2520)
);

CKINVDCx11_ASAP7_75t_R g2521 ( 
.A(n_2394),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2438),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2384),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2426),
.B(n_2216),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2411),
.A2(n_2324),
.B1(n_1643),
.B2(n_2246),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2372),
.A2(n_2210),
.B1(n_2337),
.B2(n_2339),
.Y(n_2526)
);

OAI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_2372),
.A2(n_1974),
.B1(n_2207),
.B2(n_2203),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2437),
.Y(n_2528)
);

INVx6_ASAP7_75t_L g2529 ( 
.A(n_2382),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_SL g2530 ( 
.A1(n_2467),
.A2(n_2447),
.B1(n_2173),
.B2(n_2190),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_SL g2531 ( 
.A1(n_2475),
.A2(n_2190),
.B1(n_2434),
.B2(n_1744),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_SL g2532 ( 
.A1(n_2458),
.A2(n_2069),
.B1(n_2286),
.B2(n_1947),
.Y(n_2532)
);

BUFx4f_ASAP7_75t_SL g2533 ( 
.A(n_2488),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2478),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2481),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2471),
.B(n_2219),
.Y(n_2536)
);

AOI22xp33_ASAP7_75t_L g2537 ( 
.A1(n_2468),
.A2(n_1986),
.B1(n_1820),
.B2(n_2034),
.Y(n_2537)
);

AOI22xp33_ASAP7_75t_SL g2538 ( 
.A1(n_2457),
.A2(n_2035),
.B1(n_1998),
.B2(n_2404),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2482),
.Y(n_2539)
);

OAI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2456),
.A2(n_2334),
.B1(n_2234),
.B2(n_2429),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2454),
.B(n_1999),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2486),
.A2(n_2052),
.B1(n_2338),
.B2(n_1938),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2495),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2466),
.A2(n_2021),
.B1(n_2099),
.B2(n_2284),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2496),
.Y(n_2545)
);

AOI22xp33_ASAP7_75t_L g2546 ( 
.A1(n_2510),
.A2(n_1813),
.B1(n_2107),
.B2(n_2073),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2519),
.A2(n_2107),
.B1(n_2114),
.B2(n_1868),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2492),
.A2(n_2373),
.B1(n_2432),
.B2(n_2425),
.Y(n_2548)
);

AOI22xp33_ASAP7_75t_L g2549 ( 
.A1(n_2463),
.A2(n_2158),
.B1(n_2225),
.B2(n_2102),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2497),
.B(n_1991),
.Y(n_2550)
);

AOI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_2507),
.A2(n_2158),
.B1(n_2041),
.B2(n_1865),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_L g2552 ( 
.A1(n_2461),
.A2(n_2041),
.B1(n_2167),
.B2(n_2154),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_2479),
.A2(n_2167),
.B1(n_2182),
.B2(n_2154),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2494),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2525),
.A2(n_2182),
.B1(n_2092),
.B2(n_2074),
.Y(n_2555)
);

AOI22xp33_ASAP7_75t_SL g2556 ( 
.A1(n_2483),
.A2(n_2474),
.B1(n_2465),
.B2(n_2455),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_SL g2557 ( 
.A1(n_2474),
.A2(n_2035),
.B1(n_1998),
.B2(n_1922),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2503),
.A2(n_1651),
.B1(n_2360),
.B2(n_2354),
.Y(n_2558)
);

OAI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2511),
.A2(n_2417),
.B1(n_2068),
.B2(n_2085),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2501),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2500),
.A2(n_2082),
.B1(n_2224),
.B2(n_2291),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2453),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2459),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2489),
.B(n_1992),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2527),
.A2(n_2480),
.B1(n_2526),
.B2(n_2476),
.Y(n_2565)
);

AOI222xp33_ASAP7_75t_L g2566 ( 
.A1(n_2524),
.A2(n_1902),
.B1(n_1805),
.B2(n_2260),
.C1(n_2081),
.C2(n_2029),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2506),
.A2(n_2000),
.B1(n_2003),
.B2(n_2002),
.Y(n_2567)
);

AOI22xp33_ASAP7_75t_L g2568 ( 
.A1(n_2513),
.A2(n_2027),
.B1(n_2028),
.B2(n_2013),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2460),
.A2(n_2138),
.B1(n_2146),
.B2(n_2132),
.Y(n_2569)
);

OAI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2490),
.A2(n_2343),
.B1(n_2370),
.B2(n_2445),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2494),
.B(n_2368),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2522),
.A2(n_2159),
.B1(n_2170),
.B2(n_2150),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2517),
.A2(n_2192),
.B1(n_2164),
.B2(n_2180),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2502),
.A2(n_2388),
.B1(n_2439),
.B2(n_2413),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2462),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_SL g2576 ( 
.A1(n_2518),
.A2(n_1794),
.B(n_1726),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2477),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2493),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2508),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2504),
.A2(n_2183),
.B1(n_2188),
.B2(n_2162),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2514),
.B(n_2402),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2484),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2515),
.B(n_2149),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_SL g2584 ( 
.A1(n_2455),
.A2(n_1998),
.B1(n_2035),
.B2(n_2177),
.Y(n_2584)
);

INVx8_ASAP7_75t_L g2585 ( 
.A(n_2491),
.Y(n_2585)
);

INVx3_ASAP7_75t_L g2586 ( 
.A(n_2516),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2487),
.A2(n_2195),
.B1(n_2086),
.B2(n_2105),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2465),
.A2(n_2108),
.B1(n_2122),
.B2(n_2080),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2498),
.A2(n_2126),
.B1(n_2006),
.B2(n_2016),
.Y(n_2589)
);

AOI22xp33_ASAP7_75t_L g2590 ( 
.A1(n_2521),
.A2(n_2007),
.B1(n_2019),
.B2(n_2018),
.Y(n_2590)
);

INVx4_ASAP7_75t_SL g2591 ( 
.A(n_2516),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2520),
.B(n_2155),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2509),
.B(n_2156),
.Y(n_2593)
);

OAI21xp5_ASAP7_75t_SL g2594 ( 
.A1(n_2523),
.A2(n_2176),
.B(n_2172),
.Y(n_2594)
);

OAI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2529),
.A2(n_2240),
.B1(n_2135),
.B2(n_2366),
.Y(n_2595)
);

AOI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2528),
.A2(n_2049),
.B1(n_2051),
.B2(n_2050),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2512),
.A2(n_2053),
.B1(n_2125),
.B2(n_2120),
.Y(n_2597)
);

OAI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2529),
.A2(n_2239),
.B1(n_2308),
.B2(n_2249),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2509),
.Y(n_2599)
);

BUFx3_ASAP7_75t_L g2600 ( 
.A(n_2491),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2505),
.A2(n_2353),
.B1(n_2281),
.B2(n_2441),
.Y(n_2601)
);

OR2x2_ASAP7_75t_L g2602 ( 
.A(n_2509),
.B(n_2441),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2473),
.A2(n_2130),
.B1(n_2328),
.B2(n_2437),
.Y(n_2603)
);

AOI22xp33_ASAP7_75t_SL g2604 ( 
.A1(n_2473),
.A2(n_2035),
.B1(n_2189),
.B2(n_2185),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2469),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2485),
.A2(n_2058),
.B1(n_2442),
.B2(n_2433),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2470),
.B(n_2355),
.Y(n_2607)
);

OAI21xp33_ASAP7_75t_L g2608 ( 
.A1(n_2542),
.A2(n_2024),
.B(n_2022),
.Y(n_2608)
);

OAI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2546),
.A2(n_2191),
.B1(n_2394),
.B2(n_2315),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2551),
.A2(n_2452),
.B1(n_2392),
.B2(n_2423),
.Y(n_2610)
);

NAND3xp33_ASAP7_75t_L g2611 ( 
.A(n_2537),
.B(n_2106),
.C(n_2104),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_SL g2612 ( 
.A1(n_2559),
.A2(n_2540),
.B1(n_2550),
.B2(n_2548),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2547),
.A2(n_2423),
.B1(n_2407),
.B2(n_2396),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2532),
.A2(n_2566),
.B1(n_2530),
.B2(n_2541),
.Y(n_2614)
);

OAI221xp5_ASAP7_75t_SL g2615 ( 
.A1(n_2576),
.A2(n_1902),
.B1(n_2163),
.B2(n_2416),
.C(n_2104),
.Y(n_2615)
);

AOI221xp5_ASAP7_75t_L g2616 ( 
.A1(n_2561),
.A2(n_2103),
.B1(n_2293),
.B2(n_2283),
.C(n_2292),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2544),
.A2(n_2103),
.B1(n_2437),
.B2(n_2110),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2536),
.B(n_2437),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2531),
.A2(n_2407),
.B1(n_2382),
.B2(n_2221),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2603),
.A2(n_2222),
.B1(n_2386),
.B2(n_2385),
.Y(n_2620)
);

OAI21xp33_ASAP7_75t_L g2621 ( 
.A1(n_2594),
.A2(n_2062),
.B(n_2054),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2570),
.A2(n_2110),
.B1(n_2062),
.B2(n_2075),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2565),
.A2(n_2075),
.B1(n_2076),
.B2(n_2054),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2569),
.A2(n_2451),
.B1(n_2401),
.B2(n_2472),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_2602),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2549),
.A2(n_2076),
.B1(n_2035),
.B2(n_1746),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2564),
.B(n_2363),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2576),
.A2(n_2464),
.B1(n_2129),
.B2(n_1980),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2578),
.B(n_2197),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2562),
.B(n_2563),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2555),
.A2(n_1723),
.B1(n_1736),
.B2(n_2215),
.Y(n_2631)
);

INVxp67_ASAP7_75t_L g2632 ( 
.A(n_2582),
.Y(n_2632)
);

BUFx3_ASAP7_75t_L g2633 ( 
.A(n_2533),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_SL g2634 ( 
.A1(n_2574),
.A2(n_2401),
.B1(n_2451),
.B2(n_2317),
.Y(n_2634)
);

AOI22xp33_ASAP7_75t_L g2635 ( 
.A1(n_2556),
.A2(n_2313),
.B1(n_2330),
.B2(n_2267),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2534),
.Y(n_2636)
);

AOI22xp33_ASAP7_75t_L g2637 ( 
.A1(n_2552),
.A2(n_2056),
.B1(n_2078),
.B2(n_2057),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2594),
.A2(n_1994),
.B1(n_2196),
.B2(n_2100),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2558),
.A2(n_2196),
.B1(n_2268),
.B2(n_2369),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2590),
.A2(n_2587),
.B1(n_2538),
.B2(n_2597),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2553),
.A2(n_2335),
.B1(n_2320),
.B2(n_2040),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2595),
.B(n_2369),
.Y(n_2642)
);

OA21x2_ASAP7_75t_L g2643 ( 
.A1(n_2535),
.A2(n_1711),
.B(n_2326),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_SL g2644 ( 
.A1(n_2605),
.A2(n_2369),
.B1(n_2395),
.B2(n_2389),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2593),
.B(n_2389),
.Y(n_2645)
);

OAI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_2567),
.A2(n_2389),
.B1(n_2412),
.B2(n_2395),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_SL g2647 ( 
.A1(n_2605),
.A2(n_2395),
.B1(n_2420),
.B2(n_2412),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2539),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2575),
.B(n_2412),
.Y(n_2649)
);

OAI211xp5_ASAP7_75t_SL g2650 ( 
.A1(n_2572),
.A2(n_2499),
.B(n_174),
.C(n_172),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_2573),
.A2(n_2321),
.B1(n_2342),
.B2(n_2420),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2592),
.A2(n_2321),
.B1(n_2450),
.B2(n_2420),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_2583),
.B(n_2450),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2554),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2605),
.A2(n_2450),
.B1(n_174),
.B2(n_172),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2543),
.A2(n_176),
.B1(n_173),
.B2(n_175),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_2568),
.A2(n_1800),
.B1(n_181),
.B2(n_177),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2577),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2589),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2604),
.A2(n_2588),
.B1(n_2596),
.B2(n_2581),
.Y(n_2660)
);

OAI21xp33_ASAP7_75t_L g2661 ( 
.A1(n_2580),
.A2(n_180),
.B(n_182),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2625),
.B(n_2545),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2615),
.B(n_2607),
.Y(n_2663)
);

OAI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2611),
.A2(n_2557),
.B1(n_2601),
.B2(n_2606),
.Y(n_2664)
);

NOR3xp33_ASAP7_75t_L g2665 ( 
.A(n_2650),
.B(n_2598),
.C(n_2579),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2636),
.Y(n_2666)
);

OAI21xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2612),
.A2(n_2586),
.B(n_2571),
.Y(n_2667)
);

NAND3xp33_ASAP7_75t_L g2668 ( 
.A(n_2614),
.B(n_2560),
.C(n_2599),
.Y(n_2668)
);

NAND3xp33_ASAP7_75t_L g2669 ( 
.A(n_2656),
.B(n_2584),
.C(n_2571),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2621),
.A2(n_2586),
.B1(n_2554),
.B2(n_2600),
.Y(n_2670)
);

AOI221xp5_ASAP7_75t_L g2671 ( 
.A1(n_2656),
.A2(n_2585),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_2671)
);

OAI21xp33_ASAP7_75t_L g2672 ( 
.A1(n_2661),
.A2(n_183),
.B(n_185),
.Y(n_2672)
);

OAI221xp5_ASAP7_75t_L g2673 ( 
.A1(n_2608),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.C(n_193),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2658),
.B(n_2591),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2628),
.B(n_2591),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2618),
.B(n_2585),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2648),
.B(n_2630),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2627),
.B(n_189),
.Y(n_2678)
);

OAI21xp33_ASAP7_75t_L g2679 ( 
.A1(n_2655),
.A2(n_193),
.B(n_194),
.Y(n_2679)
);

NAND4xp25_ASAP7_75t_SL g2680 ( 
.A(n_2640),
.B(n_195),
.C(n_196),
.D(n_197),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2632),
.B(n_2585),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2649),
.B(n_195),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2645),
.B(n_196),
.Y(n_2683)
);

NOR3xp33_ASAP7_75t_L g2684 ( 
.A(n_2609),
.B(n_197),
.C(n_198),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2653),
.B(n_198),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2629),
.B(n_199),
.Y(n_2686)
);

OAI221xp5_ASAP7_75t_SL g2687 ( 
.A1(n_2657),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.C(n_204),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2654),
.B(n_201),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2654),
.B(n_204),
.Y(n_2689)
);

NAND3xp33_ASAP7_75t_L g2690 ( 
.A(n_2659),
.B(n_205),
.C(n_206),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2652),
.B(n_2633),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2623),
.B(n_205),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2660),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2613),
.B(n_208),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2624),
.B(n_210),
.Y(n_2695)
);

NAND3xp33_ASAP7_75t_L g2696 ( 
.A(n_2616),
.B(n_212),
.C(n_213),
.Y(n_2696)
);

OAI211xp5_ASAP7_75t_L g2697 ( 
.A1(n_2671),
.A2(n_2647),
.B(n_2644),
.C(n_2642),
.Y(n_2697)
);

AO21x2_ASAP7_75t_L g2698 ( 
.A1(n_2684),
.A2(n_2638),
.B(n_2624),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2666),
.B(n_2634),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2677),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2662),
.Y(n_2701)
);

AO21x2_ASAP7_75t_L g2702 ( 
.A1(n_2684),
.A2(n_2646),
.B(n_2639),
.Y(n_2702)
);

NAND3xp33_ASAP7_75t_L g2703 ( 
.A(n_2696),
.B(n_2635),
.C(n_2610),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_SL g2704 ( 
.A(n_2680),
.B(n_2619),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2691),
.B(n_2641),
.Y(n_2705)
);

AOI221xp5_ASAP7_75t_L g2706 ( 
.A1(n_2673),
.A2(n_2620),
.B1(n_2622),
.B2(n_2617),
.C(n_2651),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2678),
.B(n_2643),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2664),
.B(n_2626),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2676),
.B(n_2643),
.Y(n_2709)
);

BUFx2_ASAP7_75t_L g2710 ( 
.A(n_2674),
.Y(n_2710)
);

NOR3xp33_ASAP7_75t_L g2711 ( 
.A(n_2668),
.B(n_2631),
.C(n_2637),
.Y(n_2711)
);

NOR3xp33_ASAP7_75t_L g2712 ( 
.A(n_2687),
.B(n_214),
.C(n_217),
.Y(n_2712)
);

NOR3xp33_ASAP7_75t_L g2713 ( 
.A(n_2687),
.B(n_219),
.C(n_220),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_L g2714 ( 
.A1(n_2672),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2681),
.B(n_223),
.Y(n_2715)
);

INVx1_ASAP7_75t_SL g2716 ( 
.A(n_2685),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2700),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2700),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2710),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2701),
.B(n_2683),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2707),
.B(n_2695),
.Y(n_2721)
);

INVx1_ASAP7_75t_SL g2722 ( 
.A(n_2707),
.Y(n_2722)
);

NAND4xp75_ASAP7_75t_SL g2723 ( 
.A(n_2699),
.B(n_2694),
.C(n_2663),
.D(n_2689),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2709),
.B(n_2699),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2715),
.Y(n_2725)
);

NAND4xp75_ASAP7_75t_L g2726 ( 
.A(n_2708),
.B(n_2675),
.C(n_2688),
.D(n_2682),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2715),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2715),
.Y(n_2728)
);

INVx1_ASAP7_75t_SL g2729 ( 
.A(n_2720),
.Y(n_2729)
);

OA22x2_ASAP7_75t_L g2730 ( 
.A1(n_2725),
.A2(n_2728),
.B1(n_2727),
.B2(n_2667),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2717),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2718),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2724),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2722),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2724),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2719),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2721),
.Y(n_2737)
);

XNOR2xp5_ASAP7_75t_L g2738 ( 
.A(n_2723),
.B(n_2716),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2731),
.Y(n_2739)
);

XNOR2x1_ASAP7_75t_L g2740 ( 
.A(n_2738),
.B(n_2726),
.Y(n_2740)
);

XNOR2x1_ASAP7_75t_L g2741 ( 
.A(n_2730),
.B(n_2693),
.Y(n_2741)
);

OA22x2_ASAP7_75t_L g2742 ( 
.A1(n_2729),
.A2(n_2722),
.B1(n_2697),
.B2(n_2708),
.Y(n_2742)
);

OA22x2_ASAP7_75t_L g2743 ( 
.A1(n_2733),
.A2(n_2679),
.B1(n_2713),
.B2(n_2712),
.Y(n_2743)
);

XOR2x2_ASAP7_75t_L g2744 ( 
.A(n_2737),
.B(n_2703),
.Y(n_2744)
);

AO22x2_ASAP7_75t_L g2745 ( 
.A1(n_2734),
.A2(n_2705),
.B1(n_2690),
.B2(n_2711),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2739),
.Y(n_2746)
);

OAI322xp33_ASAP7_75t_L g2747 ( 
.A1(n_2743),
.A2(n_2704),
.A3(n_2735),
.B1(n_2734),
.B2(n_2692),
.C1(n_2686),
.C2(n_2732),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2745),
.Y(n_2748)
);

INVx2_ASAP7_75t_SL g2749 ( 
.A(n_2742),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2740),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2744),
.Y(n_2751)
);

NAND2x1_ASAP7_75t_SL g2752 ( 
.A(n_2748),
.B(n_2736),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2746),
.Y(n_2753)
);

OAI322xp33_ASAP7_75t_L g2754 ( 
.A1(n_2749),
.A2(n_2741),
.A3(n_2669),
.B1(n_2714),
.B2(n_227),
.C1(n_228),
.C2(n_229),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2753),
.Y(n_2755)
);

AOI221x1_ASAP7_75t_SL g2756 ( 
.A1(n_2754),
.A2(n_2751),
.B1(n_2747),
.B2(n_2750),
.C(n_2752),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2753),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2753),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2755),
.Y(n_2759)
);

NOR4xp25_ASAP7_75t_L g2760 ( 
.A(n_2757),
.B(n_2747),
.C(n_2714),
.D(n_2706),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2758),
.A2(n_2698),
.B1(n_2702),
.B2(n_2665),
.Y(n_2761)
);

NOR4xp25_ASAP7_75t_L g2762 ( 
.A(n_2756),
.B(n_2670),
.C(n_225),
.D(n_226),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2755),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2755),
.B(n_2665),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2755),
.Y(n_2765)
);

AOI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2762),
.A2(n_2698),
.B1(n_2702),
.B2(n_228),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_SL g2767 ( 
.A(n_2760),
.B(n_224),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2759),
.Y(n_2768)
);

NOR3xp33_ASAP7_75t_L g2769 ( 
.A(n_2763),
.B(n_224),
.C(n_227),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2765),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2764),
.Y(n_2771)
);

NOR2x1_ASAP7_75t_L g2772 ( 
.A(n_2761),
.B(n_231),
.Y(n_2772)
);

NAND4xp25_ASAP7_75t_L g2773 ( 
.A(n_2766),
.B(n_231),
.C(n_233),
.D(n_234),
.Y(n_2773)
);

NAND4xp25_ASAP7_75t_L g2774 ( 
.A(n_2767),
.B(n_233),
.C(n_234),
.D(n_235),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2771),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_2775)
);

AO22x2_ASAP7_75t_L g2776 ( 
.A1(n_2768),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2770),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2769),
.B(n_2772),
.Y(n_2778)
);

NOR4xp25_ASAP7_75t_L g2779 ( 
.A(n_2767),
.B(n_239),
.C(n_240),
.D(n_241),
.Y(n_2779)
);

OAI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2773),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2776),
.Y(n_2781)
);

CKINVDCx20_ASAP7_75t_R g2782 ( 
.A(n_2775),
.Y(n_2782)
);

INVx8_ASAP7_75t_L g2783 ( 
.A(n_2778),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2777),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2779),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2774),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2776),
.Y(n_2787)
);

CKINVDCx20_ASAP7_75t_R g2788 ( 
.A(n_2775),
.Y(n_2788)
);

AO22x2_ASAP7_75t_L g2789 ( 
.A1(n_2781),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_2789)
);

OAI22x1_ASAP7_75t_L g2790 ( 
.A1(n_2785),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2782),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_2791)
);

AOI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2788),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_2792)
);

INVxp67_ASAP7_75t_L g2793 ( 
.A(n_2787),
.Y(n_2793)
);

OAI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2786),
.A2(n_2783),
.B1(n_2784),
.B2(n_2780),
.Y(n_2794)
);

OAI22x1_ASAP7_75t_L g2795 ( 
.A1(n_2783),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_2795)
);

AOI22xp33_ASAP7_75t_L g2796 ( 
.A1(n_2783),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2782),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2789),
.Y(n_2798)
);

INVxp67_ASAP7_75t_SL g2799 ( 
.A(n_2795),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2789),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2790),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2797),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2793),
.Y(n_2803)
);

AOI221xp5_ASAP7_75t_L g2804 ( 
.A1(n_2799),
.A2(n_2794),
.B1(n_2796),
.B2(n_2792),
.C(n_2791),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2803),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_SL g2806 ( 
.A1(n_2801),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2802),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2806),
.Y(n_2808)
);

OAI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2808),
.A2(n_2798),
.B1(n_2800),
.B2(n_2804),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2809),
.Y(n_2810)
);

AOI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2810),
.A2(n_2807),
.B1(n_2805),
.B2(n_270),
.C(n_272),
.Y(n_2811)
);

AOI211xp5_ASAP7_75t_L g2812 ( 
.A1(n_2811),
.A2(n_266),
.B(n_268),
.C(n_270),
.Y(n_2812)
);


endmodule