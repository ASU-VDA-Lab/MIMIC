module fake_jpeg_15534_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_46),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_26),
.B1(n_21),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_51),
.B1(n_74),
.B2(n_29),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_26),
.B1(n_21),
.B2(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_66),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_34),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_39),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_42),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_68),
.C(n_61),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_87),
.C(n_31),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_104),
.B1(n_34),
.B2(n_31),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2x1_ASAP7_75t_R g119 ( 
.A(n_91),
.B(n_28),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_39),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_31),
.B(n_29),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_44),
.B1(n_60),
.B2(n_45),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_69),
.B1(n_44),
.B2(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_107),
.B1(n_115),
.B2(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_64),
.B1(n_48),
.B2(n_53),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_120),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_67),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_102),
.B(n_76),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_48),
.B1(n_59),
.B2(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_87),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_76),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_46),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_129),
.C(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_129),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_48),
.B1(n_59),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_77),
.A2(n_48),
.B1(n_47),
.B2(n_41),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_90),
.B1(n_85),
.B2(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_97),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_138),
.B(n_144),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_96),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_145),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_96),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_22),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_128),
.B1(n_131),
.B2(n_106),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_160),
.B(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_103),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_121),
.B(n_119),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_107),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_29),
.B(n_34),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_105),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_169),
.C(n_177),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_170),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_130),
.B(n_115),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_131),
.C(n_106),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_117),
.B(n_122),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_109),
.B1(n_85),
.B2(n_117),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_175),
.B1(n_182),
.B2(n_183),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_23),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_133),
.B1(n_41),
.B2(n_47),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_126),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_185),
.C(n_38),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_35),
.B(n_25),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_181),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_25),
.B(n_30),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_159),
.B1(n_154),
.B2(n_142),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_92),
.B1(n_81),
.B2(n_110),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_38),
.C(n_111),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_140),
.B1(n_141),
.B2(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_141),
.B1(n_145),
.B2(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_137),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_203),
.C(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_158),
.B1(n_161),
.B2(n_139),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_143),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_215),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_208),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_151),
.B1(n_139),
.B2(n_109),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_152),
.B1(n_134),
.B2(n_111),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_173),
.B1(n_186),
.B2(n_175),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_63),
.C(n_33),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_152),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_17),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_17),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_23),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_63),
.C(n_47),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_28),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_188),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_163),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_232),
.C(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_170),
.C(n_162),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_167),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_214),
.C(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_210),
.B1(n_188),
.B2(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_181),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_175),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_33),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_240),
.C(n_88),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_33),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_88),
.B1(n_83),
.B2(n_47),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_41),
.C(n_83),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_193),
.C(n_207),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_252),
.C(n_27),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_218),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_244),
.B(n_253),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_193),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_248),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_204),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_235),
.B(n_9),
.Y(n_269)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_254),
.B1(n_259),
.B2(n_27),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_204),
.B1(n_200),
.B2(n_12),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_30),
.B1(n_33),
.B2(n_18),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_10),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_263),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_261),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_239),
.C(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_234),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_27),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_267),
.C(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_228),
.B1(n_237),
.B2(n_221),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_219),
.C(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_272),
.Y(n_295)
);

AO221x1_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_27),
.B1(n_18),
.B2(n_9),
.C(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_248),
.C(n_249),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_7),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_281),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_7),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_296),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_290),
.C(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_11),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_293),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_241),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_15),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_18),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_14),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_273),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_308),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_275),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_307),
.C(n_312),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_269),
.B(n_268),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_0),
.B(n_1),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_276),
.C(n_266),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_276),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_279),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_282),
.C(n_272),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_292),
.B(n_298),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_309),
.B(n_4),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_303),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_322),
.B(n_323),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_304),
.B(n_2),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_3),
.B(n_4),
.Y(n_323)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_328),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_3),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_315),
.B(n_313),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_336),
.B(n_337),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_335),
.B(n_3),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_316),
.B(n_319),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_339),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_5),
.B(n_6),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_343),
.Y(n_344)
);


endmodule