module fake_jpeg_21044_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_46),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_8),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_60),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_55),
.B1(n_38),
.B2(n_39),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_70),
.B1(n_86),
.B2(n_99),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_69),
.B(n_71),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_23),
.B1(n_49),
.B2(n_40),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_23),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_22),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_48),
.B(n_40),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_31),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_38),
.B1(n_37),
.B2(n_45),
.Y(n_86)
);

OA22x2_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_31),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_33),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

AO22x2_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_48),
.B1(n_49),
.B2(n_44),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_32),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_21),
.B1(n_34),
.B2(n_25),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_25),
.B1(n_34),
.B2(n_21),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_116),
.B1(n_92),
.B2(n_91),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_108),
.A2(n_114),
.B(n_117),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_109),
.A2(n_130),
.B1(n_131),
.B2(n_12),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_42),
.C(n_43),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_129),
.C(n_36),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_31),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_44),
.B1(n_43),
.B2(n_26),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_31),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_98),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_36),
.C(n_19),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_27),
.B1(n_35),
.B2(n_26),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_18),
.B1(n_35),
.B2(n_27),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_18),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_110),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_137),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_100),
.B1(n_82),
.B2(n_74),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_139),
.B1(n_152),
.B2(n_128),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_143),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_96),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_123),
.B(n_3),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_106),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_92),
.B1(n_97),
.B2(n_84),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_20),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_26),
.B1(n_35),
.B2(n_19),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_111),
.B1(n_121),
.B2(n_128),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_105),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_105),
.B(n_124),
.C(n_103),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_0),
.B(n_2),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_162),
.B(n_173),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_127),
.B1(n_118),
.B2(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_177),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_121),
.B1(n_118),
.B2(n_111),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_168),
.B1(n_179),
.B2(n_145),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_160),
.C(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_103),
.B1(n_124),
.B2(n_30),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_123),
.B1(n_13),
.B2(n_14),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_192),
.B1(n_157),
.B2(n_147),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_20),
.B(n_3),
.Y(n_220)
);

AO21x2_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_140),
.B(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_2),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_12),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_190),
.B(n_134),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_194),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_135),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_203),
.B1(n_217),
.B2(n_177),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_200),
.B(n_174),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_160),
.B(n_156),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_220),
.B(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_151),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_200),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_147),
.B1(n_138),
.B2(n_136),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_222),
.B1(n_223),
.B2(n_180),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_154),
.B1(n_158),
.B2(n_14),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_180),
.B1(n_189),
.B2(n_29),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_36),
.C(n_30),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_219),
.C(n_4),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_20),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_172),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_182),
.B(n_171),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_187),
.C(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_36),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_176),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_226),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_231),
.B1(n_236),
.B2(n_210),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_212),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_188),
.B1(n_165),
.B2(n_187),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_188),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_243),
.C(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_165),
.B1(n_171),
.B2(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_174),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_199),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_196),
.A2(n_2),
.B1(n_4),
.B2(n_16),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_197),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_252),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_209),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_229),
.B1(n_218),
.B2(n_245),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_256),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_268),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_233),
.C(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_195),
.C(n_207),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_226),
.C(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_211),
.B1(n_193),
.B2(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_265),
.B1(n_238),
.B2(n_221),
.Y(n_284)
);

OAI22x1_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_218),
.B1(n_203),
.B2(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_213),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_220),
.C(n_206),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_232),
.B(n_214),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_205),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_264),
.B1(n_269),
.B2(n_252),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_255),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_237),
.B1(n_249),
.B2(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_290),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_241),
.C(n_205),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.C(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_246),
.C(n_5),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_4),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_259),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_297),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_251),
.B(n_253),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_296),
.Y(n_311)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_289),
.B1(n_286),
.B2(n_276),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_301),
.C(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_5),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_275),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_273),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_272),
.C(n_281),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_285),
.C(n_272),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_309),
.C(n_292),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_278),
.C(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_316),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_277),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_300),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_323),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_293),
.B(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_277),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_308),
.C(n_313),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_326),
.B(n_306),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

INVx11_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_278),
.B1(n_318),
.B2(n_294),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_332),
.Y(n_336)
);

AO21x2_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_333),
.B(n_334),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_309),
.C(n_313),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_290),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_321),
.B(n_322),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_338),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_329),
.B(n_326),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_336),
.C(n_337),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_330),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_15),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_7),
.C(n_9),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_9),
.Y(n_345)
);


endmodule