module fake_jpeg_20990_n_77 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_21),
.B(n_18),
.Y(n_26)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_9),
.Y(n_35)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_46),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_8),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_8),
.B(n_12),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_20),
.C(n_25),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_30),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_41),
.B(n_46),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_33),
.B1(n_12),
.B2(n_21),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_34),
.B1(n_14),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_14),
.B1(n_17),
.B2(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_15),
.B1(n_17),
.B2(n_16),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_39),
.C(n_28),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_45),
.B(n_38),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_53),
.Y(n_64)
);

BUFx12f_ASAP7_75t_SL g65 ( 
.A(n_58),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_54),
.B1(n_52),
.B2(n_58),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_62),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.C(n_71),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_57),
.B(n_7),
.C(n_5),
.D(n_3),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_50),
.C(n_1),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_0),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_72),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_3),
.B(n_4),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_3),
.Y(n_77)
);


endmodule