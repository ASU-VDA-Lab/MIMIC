module fake_jpeg_21073_n_174 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_29),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_31),
.B1(n_33),
.B2(n_15),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_21),
.B(n_26),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_29),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_14),
.B1(n_15),
.B2(n_25),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_26),
.B1(n_25),
.B2(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_46),
.B1(n_31),
.B2(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_71),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_20),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_34),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_18),
.B1(n_28),
.B2(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_87),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_42),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_55),
.A3(n_38),
.B1(n_54),
.B2(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_23),
.B(n_22),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_51),
.B1(n_23),
.B2(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_107),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_73),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_79),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_74),
.B1(n_69),
.B2(n_81),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_73),
.B(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_96),
.B1(n_103),
.B2(n_97),
.Y(n_132)
);

AOI21x1_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_80),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_110),
.C(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_112),
.C(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_135),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_108),
.B1(n_105),
.B2(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_137),
.B1(n_129),
.B2(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_93),
.B1(n_16),
.B2(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_139),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_113),
.A3(n_124),
.B1(n_114),
.B2(n_121),
.C(n_126),
.Y(n_140)
);

AOI31xp67_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_149),
.A3(n_8),
.B(n_13),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_116),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.C(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_111),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_148),
.A2(n_133),
.B1(n_131),
.B2(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_7),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_153),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_156),
.C(n_146),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_9),
.B(n_12),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_161),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_141),
.B(n_140),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_160),
.B(n_163),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_135),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_12),
.C(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_170),
.B(n_1),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_169),
.B(n_5),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.Y(n_174)
);


endmodule