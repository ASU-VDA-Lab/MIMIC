module fake_jpeg_26732_n_176 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_13),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_21),
.B1(n_14),
.B2(n_20),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_29),
.B(n_25),
.C(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_22),
.B1(n_16),
.B2(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_27),
.Y(n_52)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_47),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_55),
.B1(n_34),
.B2(n_40),
.Y(n_56)
);

NAND2x1_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_24),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

AOI22x1_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_29),
.B1(n_40),
.B2(n_36),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_40),
.B1(n_34),
.B2(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_27),
.C(n_23),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_19),
.B(n_18),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_66),
.C(n_60),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_48),
.B1(n_45),
.B2(n_51),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_11),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_36),
.B1(n_38),
.B2(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_72),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_35),
.B(n_12),
.C(n_13),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_49),
.B(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_80),
.B(n_84),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_43),
.B(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_89),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_42),
.B(n_19),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_85),
.B(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_92),
.B1(n_89),
.B2(n_70),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_22),
.B(n_16),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_73),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_0),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_3),
.C(n_5),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_54),
.B(n_24),
.C(n_14),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_73),
.B(n_1),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_19),
.B1(n_20),
.B2(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_0),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_91),
.B(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_65),
.C(n_7),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_79),
.C(n_81),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_91),
.B1(n_5),
.B2(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_85),
.B(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_113),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_79),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_124),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_125),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_93),
.B1(n_84),
.B2(n_92),
.C(n_87),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_109),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_91),
.B(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_91),
.C(n_5),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_105),
.C(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_104),
.B1(n_106),
.B2(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_99),
.B1(n_98),
.B2(n_97),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_129),
.B1(n_130),
.B2(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_127),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_144),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_119),
.C(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_136),
.C(n_132),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_127),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_133),
.B(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_131),
.B1(n_126),
.B2(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_157),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_140),
.B(n_117),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_147),
.B(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_146),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_161),
.C(n_103),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_157),
.B1(n_151),
.B2(n_108),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_128),
.B1(n_103),
.B2(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_102),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_110),
.B(n_162),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_100),
.C(n_9),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_166),
.B1(n_165),
.B2(n_10),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_2),
.B1(n_10),
.B2(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_2),
.Y(n_176)
);


endmodule