module fake_netlist_6_1737_n_77 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_77);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_77;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_27;
wire n_38;
wire n_61;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_5),
.B1(n_0),
.B2(n_11),
.Y(n_28)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_0),
.B(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_15),
.B1(n_2),
.B2(n_10),
.Y(n_35)
);

OA21x2_ASAP7_75t_L g36 ( 
.A1(n_16),
.A2(n_3),
.B(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_36),
.B1(n_26),
.B2(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_30),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_25),
.B(n_33),
.C(n_30),
.Y(n_46)
);

AND3x4_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_28),
.C(n_35),
.Y(n_47)
);

OAI21x1_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_29),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_24),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_39),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_46),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_56),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_52),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_26),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_58),
.B(n_63),
.C(n_60),
.Y(n_66)
);

AOI211xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_33),
.B(n_45),
.C(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_65),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_29),
.C(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_47),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_57),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_24),
.B1(n_27),
.B2(n_75),
.Y(n_76)
);

OR2x6_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_27),
.Y(n_77)
);


endmodule