module fake_jpeg_8173_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_4),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_5),
.A2(n_1),
.B(n_8),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_18),
.B1(n_11),
.B2(n_20),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_2),
.C(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.Y(n_31)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_18),
.B1(n_13),
.B2(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_35),
.B1(n_39),
.B2(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_20),
.B1(n_12),
.B2(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_57),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_36),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_42),
.C(n_49),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_51),
.B(n_47),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_65),
.B1(n_52),
.B2(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.C(n_55),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_51),
.C(n_33),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_69),
.C(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_72),
.B1(n_69),
.B2(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_68),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_48),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_R g76 ( 
.A1(n_73),
.A2(n_67),
.B(n_69),
.C(n_26),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_67),
.C(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);


endmodule