module fake_jpeg_21100_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_46),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_17),
.B1(n_16),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_74),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_34),
.B1(n_36),
.B2(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_16),
.B1(n_32),
.B2(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_16),
.B1(n_32),
.B2(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_89),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

OA22x2_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_42),
.B1(n_44),
.B2(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_102),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_37),
.B1(n_22),
.B2(n_18),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_100),
.B1(n_108),
.B2(n_113),
.Y(n_128)
);

AND2x4_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_44),
.B1(n_18),
.B2(n_27),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_104),
.C(n_55),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_23),
.B1(n_49),
.B2(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_65),
.B1(n_54),
.B2(n_73),
.Y(n_122)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_13),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_42),
.B(n_23),
.C(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

AOI22x1_ASAP7_75t_SL g110 ( 
.A1(n_52),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_33),
.B(n_1),
.C(n_2),
.Y(n_141)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_54),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_115),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_29),
.B1(n_11),
.B2(n_15),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_70),
.C(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_105),
.C(n_115),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_122),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_176)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_90),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_65),
.B1(n_70),
.B2(n_63),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_54),
.B1(n_75),
.B2(n_70),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_75),
.B1(n_65),
.B2(n_64),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_135),
.B1(n_86),
.B2(n_91),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_30),
.B1(n_28),
.B2(n_15),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_30),
.B1(n_28),
.B2(n_33),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_83),
.B(n_14),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_108),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_144),
.B(n_80),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_0),
.B(n_2),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_84),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_154),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_158),
.Y(n_194)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_79),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_164),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_92),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_92),
.B1(n_115),
.B2(n_98),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_136),
.B1(n_122),
.B2(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_115),
.C(n_85),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_154),
.C(n_155),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_170),
.B(n_178),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_82),
.B1(n_109),
.B2(n_97),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_81),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_174),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_81),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_111),
.B1(n_86),
.B2(n_91),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_93),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_145),
.B1(n_134),
.B2(n_149),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_0),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_14),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_120),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_3),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_116),
.B1(n_148),
.B2(n_151),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_132),
.B1(n_144),
.B2(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_205),
.B1(n_208),
.B2(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_195),
.B(n_199),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_130),
.B(n_141),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_128),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_206),
.B(n_6),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_130),
.B1(n_125),
.B2(n_116),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_159),
.C(n_163),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_137),
.B1(n_151),
.B2(n_116),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_117),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_178),
.B(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_178),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_117),
.B(n_123),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_168),
.B(n_170),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_147),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_225),
.B1(n_232),
.B2(n_199),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_219),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_229),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_222),
.B(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_160),
.B1(n_170),
.B2(n_168),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_174),
.B(n_152),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_159),
.B1(n_176),
.B2(n_163),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_180),
.C(n_156),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_123),
.A3(n_4),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_3),
.C(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_243),
.B1(n_196),
.B2(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_241),
.B1(n_210),
.B2(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_9),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_10),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_188),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_186),
.B1(n_201),
.B2(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_247),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_223),
.B(n_221),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_194),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_228),
.B1(n_222),
.B2(n_231),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_189),
.B1(n_213),
.B2(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_207),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_200),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_189),
.B1(n_191),
.B2(n_193),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_228),
.B1(n_223),
.B2(n_238),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_193),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_230),
.C(n_216),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_268),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_250),
.A2(n_252),
.B1(n_244),
.B2(n_231),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_248),
.A2(n_235),
.B1(n_236),
.B2(n_234),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

OAI22x1_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_197),
.B1(n_237),
.B2(n_232),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_204),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_204),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_249),
.C(n_192),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_246),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_246),
.C(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_296),
.C(n_297),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_290),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_259),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_261),
.C(n_264),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_242),
.C(n_243),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_305),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_303),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_267),
.B1(n_269),
.B2(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_268),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_300),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_271),
.B1(n_266),
.B2(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_289),
.C(n_297),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_312),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_305),
.B(n_280),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_269),
.B(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_279),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_315),
.C(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_318),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_321),
.C(n_313),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_309),
.B1(n_310),
.B2(n_295),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_316),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_318),
.B(n_217),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_217),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_192),
.B(n_325),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_195),
.B(n_313),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_204),
.B(n_290),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_302),
.C(n_327),
.Y(n_332)
);


endmodule