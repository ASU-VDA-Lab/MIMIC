module fake_jpeg_6887_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

OR2x2_ASAP7_75t_SL g11 ( 
.A(n_10),
.B(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_1),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_14),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_34),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_38),
.B1(n_20),
.B2(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_26),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_12),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_22),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_19),
.B(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_33),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_30),
.A3(n_31),
.B1(n_25),
.B2(n_16),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_37),
.C(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_63),
.B1(n_65),
.B2(n_46),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_40),
.B1(n_30),
.B2(n_23),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_23),
.B1(n_40),
.B2(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_72),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_45),
.B1(n_50),
.B2(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_0),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_67),
.B(n_66),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_54),
.C(n_5),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_64),
.C(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_66),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_84),
.CI(n_77),
.CON(n_86),
.SN(n_86)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_72),
.B(n_69),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_90),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_91),
.B1(n_81),
.B2(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_87),
.B(n_73),
.C(n_6),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_63),
.B1(n_79),
.B2(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_86),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_73),
.B(n_74),
.Y(n_98)
);

AOI31xp67_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_94),
.A3(n_92),
.B(n_8),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.A3(n_2),
.B1(n_3),
.B2(n_59),
.C1(n_75),
.C2(n_99),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_92),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_75),
.C(n_59),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_103),
.Y(n_106)
);


endmodule