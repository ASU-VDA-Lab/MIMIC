module fake_jpeg_8423_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_SL g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_4),
.Y(n_15)
);

AOI21xp33_ASAP7_75t_L g16 ( 
.A1(n_0),
.A2(n_6),
.B(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_23),
.B1(n_25),
.B2(n_17),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_24),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_10),
.Y(n_32)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_2),
.B1(n_6),
.B2(n_11),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_13),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_16),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_10),
.C(n_12),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_30),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_22),
.C(n_20),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_14),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_26),
.B1(n_23),
.B2(n_27),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_34),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.C(n_26),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_26),
.B(n_12),
.C(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_46),
.B(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_9),
.B1(n_19),
.B2(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_9),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_53),
.B(n_21),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_53),
.B(n_19),
.Y(n_56)
);


endmodule