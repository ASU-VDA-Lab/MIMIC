module fake_jpeg_11669_n_62 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_56;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_5),
.B1(n_7),
.B2(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_42),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.C(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_41),
.C(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_46),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_48),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_45),
.C(n_23),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_56),
.A3(n_20),
.B1(n_31),
.B2(n_30),
.C(n_25),
.Y(n_58)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_38),
.A3(n_32),
.B1(n_27),
.B2(n_26),
.C1(n_28),
.C2(n_20),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_34),
.B(n_21),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_30),
.C(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_43),
.Y(n_62)
);


endmodule