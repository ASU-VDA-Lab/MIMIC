module fake_jpeg_2368_n_59 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_20),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_15),
.C(n_14),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_16),
.B(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_18),
.B(n_19),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_21),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_19),
.B(n_18),
.C(n_24),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_29),
.B(n_30),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_28),
.B1(n_29),
.B2(n_21),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_1),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_38),
.B(n_19),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_4),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_13),
.B(n_10),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_5),
.C(n_6),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_49),
.B1(n_7),
.B2(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_46),
.B(n_11),
.C(n_12),
.D(n_9),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_54),
.C(n_11),
.Y(n_57)
);

AOI211xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_56),
.B(n_55),
.C(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule