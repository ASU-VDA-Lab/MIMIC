module fake_jpeg_21076_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_38),
.Y(n_44)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_31),
.B1(n_16),
.B2(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_55),
.B1(n_36),
.B2(n_38),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_31),
.B1(n_16),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_39),
.B1(n_24),
.B2(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_31),
.B1(n_16),
.B2(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_86),
.B1(n_55),
.B2(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_21),
.B1(n_33),
.B2(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_19),
.B1(n_44),
.B2(n_57),
.Y(n_87)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_66),
.B1(n_69),
.B2(n_23),
.Y(n_100)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_57),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_71),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_18),
.B(n_25),
.C(n_24),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_23),
.A3(n_29),
.B1(n_44),
.B2(n_26),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_81),
.B1(n_73),
.B2(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_28),
.B(n_21),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_0),
.B(n_1),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_18),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_29),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_96),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_82),
.B1(n_65),
.B2(n_60),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_96),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_105),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_57),
.B1(n_44),
.B2(n_29),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_111),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_61),
.C(n_63),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_8),
.C(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_5),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_66),
.B1(n_62),
.B2(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_83),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_135),
.C(n_101),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_122),
.B1(n_132),
.B2(n_133),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_111),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_15),
.Y(n_121)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_124),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_130),
.B1(n_102),
.B2(n_106),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_106),
.B1(n_102),
.B2(n_111),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_99),
.B(n_108),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_139),
.B(n_154),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_87),
.B(n_105),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_96),
.B(n_98),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_88),
.B(n_90),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_116),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_122),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_95),
.B(n_111),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_161),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_126),
.B(n_104),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_163),
.B(n_174),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_119),
.B(n_133),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_144),
.C(n_139),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_132),
.B1(n_123),
.B2(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_171),
.B1(n_173),
.B2(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_115),
.B1(n_134),
.B2(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_156),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_94),
.B(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_184),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_166),
.A2(n_141),
.B1(n_157),
.B2(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_153),
.C(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_138),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_161),
.A2(n_150),
.B1(n_107),
.B2(n_13),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_160),
.Y(n_202)
);

XOR2x2_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_199),
.B(n_177),
.Y(n_207)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_172),
.C(n_173),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_179),
.C(n_187),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_164),
.B(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_188),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_181),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_186),
.CI(n_184),
.CON(n_206),
.SN(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_192),
.B1(n_201),
.B2(n_199),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_160),
.C(n_176),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_170),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_214),
.B(n_211),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_200),
.B(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_208),
.B1(n_205),
.B2(n_209),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_221),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_175),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_222),
.A3(n_218),
.B1(n_174),
.B2(n_206),
.C1(n_191),
.C2(n_160),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B1(n_223),
.B2(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_12),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_13),
.Y(n_231)
);


endmodule