module fake_jpeg_15249_n_330 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_23),
.Y(n_87)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_23),
.B1(n_29),
.B2(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_28),
.B1(n_14),
.B2(n_30),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_56),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_38),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_11),
.Y(n_104)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_37),
.B1(n_38),
.B2(n_26),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_89),
.B(n_0),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_79),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_33),
.C(n_29),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_80),
.A2(n_32),
.B(n_36),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_88),
.Y(n_145)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_20),
.C(n_21),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_87),
.B(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_28),
.B1(n_33),
.B2(n_14),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_117),
.B1(n_69),
.B2(n_59),
.Y(n_128)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_36),
.B1(n_2),
.B2(n_4),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_104),
.A2(n_113),
.B1(n_2),
.B2(n_4),
.Y(n_155)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_112),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_22),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_22),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_21),
.B1(n_15),
.B2(n_31),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_133),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_65),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_152),
.C(n_158),
.Y(n_200)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_160),
.B(n_151),
.Y(n_193)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_161),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_64),
.B1(n_66),
.B2(n_52),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_6),
.B1(n_136),
.B2(n_139),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_54),
.B1(n_32),
.B2(n_31),
.Y(n_131)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_22),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_50),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_144),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_43),
.B1(n_67),
.B2(n_63),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_73),
.B1(n_103),
.B2(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_15),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_114),
.B1(n_109),
.B2(n_103),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_2),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_32),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_4),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_109),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_70),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_73),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_180),
.B(n_186),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_200),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_188),
.B1(n_195),
.B2(n_147),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_100),
.B1(n_114),
.B2(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_178),
.B1(n_187),
.B2(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_94),
.B1(n_82),
.B2(n_99),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_185),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_77),
.B(n_101),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_77),
.C(n_101),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_165),
.C(n_174),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_146),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_85),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_124),
.A2(n_99),
.B1(n_5),
.B2(n_6),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_5),
.B1(n_6),
.B2(n_159),
.Y(n_188)
);

XOR2x1_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_160),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_193),
.B(n_194),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_122),
.A2(n_149),
.B(n_134),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_139),
.A2(n_126),
.B1(n_130),
.B2(n_145),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_139),
.B1(n_126),
.B2(n_145),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_163),
.B(n_140),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_121),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_211),
.B1(n_218),
.B2(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_214),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_123),
.B1(n_153),
.B2(n_125),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_219),
.B1(n_228),
.B2(n_171),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_215),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_156),
.B1(n_157),
.B2(n_121),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_133),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_225),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_190),
.B(n_164),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_188),
.A3(n_195),
.B1(n_174),
.B2(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_176),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_184),
.C(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_181),
.A2(n_168),
.B1(n_171),
.B2(n_177),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_182),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_194),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_183),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_173),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

A2O1A1O1Ixp25_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_183),
.B(n_164),
.C(n_184),
.D(n_187),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_235),
.A2(n_217),
.B(n_208),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_207),
.B1(n_212),
.B2(n_223),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_248),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_201),
.A2(n_178),
.B1(n_173),
.B2(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_250),
.B1(n_251),
.B2(n_213),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_169),
.C(n_199),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_169),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_186),
.C(n_166),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_186),
.C(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_219),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_224),
.B1(n_228),
.B2(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_259),
.B(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_270),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_209),
.B(n_211),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_267),
.B(n_271),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_209),
.B(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_278),
.C(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_231),
.B(n_202),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_203),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_275),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_243),
.A2(n_245),
.B1(n_242),
.B2(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_204),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_206),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_278),
.B(n_253),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_206),
.Y(n_278)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_238),
.A3(n_235),
.B1(n_247),
.B2(n_240),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.C(n_291),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_236),
.C(n_248),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_273),
.B(n_275),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_236),
.C(n_244),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_276),
.A3(n_269),
.B1(n_266),
.B2(n_267),
.C1(n_277),
.C2(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_265),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_305),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_280),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_251),
.B(n_274),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_302),
.B(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_233),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_261),
.B(n_268),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_291),
.C(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_306),
.C(n_292),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_260),
.B(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_237),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_284),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_270),
.B1(n_288),
.B2(n_290),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_280),
.C(n_283),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_300),
.A3(n_304),
.B1(n_302),
.B2(n_296),
.C1(n_305),
.C2(n_288),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_255),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_264),
.A3(n_286),
.B1(n_297),
.B2(n_298),
.C1(n_299),
.C2(n_303),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_257),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_321),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_308),
.B(n_314),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_321),
.B(n_316),
.C(n_313),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_206),
.Y(n_330)
);


endmodule