module fake_aes_4224_n_554 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_554);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_554;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_67;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g66 ( .A(n_39), .Y(n_66) );
CKINVDCx16_ASAP7_75t_R g67 ( .A(n_12), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_24), .Y(n_68) );
CKINVDCx5p33_ASAP7_75t_R g69 ( .A(n_29), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_38), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_40), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_63), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_48), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_46), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_23), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_2), .Y(n_76) );
BUFx6f_ASAP7_75t_L g77 ( .A(n_61), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_5), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_52), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_50), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
CKINVDCx14_ASAP7_75t_R g82 ( .A(n_49), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVx3_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_43), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_15), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_56), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_31), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_41), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_6), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_44), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_26), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_25), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_45), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_51), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_47), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_32), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_30), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_79), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_77), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_81), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_86), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_86), .B(n_0), .Y(n_112) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_84), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_88), .B(n_0), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_98), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_88), .B(n_1), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_67), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_86), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
AND2x6_ASAP7_75t_L g122 ( .A(n_104), .B(n_37), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_78), .B(n_1), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_77), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_92), .B(n_3), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_92), .B(n_3), .Y(n_127) );
BUFx8_ASAP7_75t_L g128 ( .A(n_75), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_76), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_129) );
INVx8_ASAP7_75t_L g130 ( .A(n_122), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g131 ( .A(n_128), .B(n_85), .C(n_99), .Y(n_131) );
BUFx8_ASAP7_75t_SL g132 ( .A(n_118), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_126), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
BUFx10_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_111), .B(n_87), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_111), .B(n_66), .Y(n_141) );
AO22x2_ASAP7_75t_L g142 ( .A1(n_112), .A2(n_104), .B1(n_75), .B2(n_76), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_125), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_109), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_126), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_111), .B(n_69), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_106), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_110), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_113), .B(n_68), .Y(n_154) );
NAND3xp33_ASAP7_75t_L g155 ( .A(n_128), .B(n_94), .C(n_102), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_125), .B(n_103), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_113), .B(n_94), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_142), .A2(n_127), .B1(n_128), .B2(n_129), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_140), .B(n_128), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_147), .B(n_107), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_141), .B(n_120), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_131), .B(n_109), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_157), .B(n_120), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_145), .B(n_121), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_134), .A2(n_122), .B(n_121), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_157), .B(n_119), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_133), .B(n_123), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_157), .B(n_122), .Y(n_175) );
NOR2xp67_ASAP7_75t_SL g176 ( .A(n_138), .B(n_69), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_142), .B(n_127), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_157), .B(n_119), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_157), .B(n_127), .Y(n_181) );
OAI221xp5_ASAP7_75t_L g182 ( .A1(n_154), .A2(n_129), .B1(n_114), .B2(n_117), .C(n_89), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_157), .B(n_127), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_158), .A2(n_105), .B1(n_116), .B2(n_94), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_136), .B(n_122), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_142), .B(n_82), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_142), .A2(n_122), .B1(n_71), .B2(n_90), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_143), .A2(n_122), .B1(n_94), .B2(n_70), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_138), .B(n_71), .Y(n_190) );
NOR2x1_ASAP7_75t_R g191 ( .A(n_133), .B(n_102), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_148), .B(n_90), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_138), .B(n_91), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_151), .B(n_91), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
BUFx8_ASAP7_75t_L g197 ( .A(n_193), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_182), .A2(n_158), .B(n_155), .C(n_72), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_196), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
OAI22x1_ASAP7_75t_L g202 ( .A1(n_159), .A2(n_188), .B1(n_193), .B2(n_187), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_146), .B1(n_158), .B2(n_130), .Y(n_204) );
INVx6_ASAP7_75t_L g205 ( .A(n_177), .Y(n_205) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_171), .A2(n_73), .B(n_80), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_163), .B(n_137), .Y(n_207) );
AO22x1_ASAP7_75t_L g208 ( .A1(n_187), .A2(n_132), .B1(n_97), .B2(n_100), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_177), .B(n_137), .Y(n_209) );
AOI21xp33_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_146), .B(n_100), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_161), .B(n_137), .Y(n_211) );
OR2x6_ASAP7_75t_SL g212 ( .A(n_191), .B(n_132), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_188), .B(n_97), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_171), .A2(n_83), .B(n_95), .C(n_96), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g215 ( .A1(n_186), .A2(n_101), .B(n_124), .C(n_115), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_164), .B(n_94), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_192), .B(n_4), .Y(n_217) );
AOI22x1_ASAP7_75t_L g218 ( .A1(n_196), .A2(n_110), .B1(n_115), .B2(n_124), .Y(n_218) );
NOR2x1_ASAP7_75t_L g219 ( .A(n_185), .B(n_156), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_195), .B(n_7), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_186), .A2(n_156), .B(n_153), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_SL g222 ( .A1(n_175), .A2(n_124), .B(n_115), .C(n_153), .Y(n_222) );
AO22x1_ASAP7_75t_L g223 ( .A1(n_191), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_175), .A2(n_150), .B(n_149), .Y(n_224) );
O2A1O1Ixp5_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_150), .B(n_106), .C(n_149), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_179), .B(n_169), .Y(n_226) );
AO21x1_ASAP7_75t_L g227 ( .A1(n_179), .A2(n_106), .B(n_9), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_183), .A2(n_106), .B1(n_11), .B2(n_12), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_169), .A2(n_152), .B(n_149), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_168), .A2(n_106), .B(n_152), .C(n_149), .Y(n_230) );
AO21x1_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_8), .B(n_11), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
NOR2x1_ASAP7_75t_L g234 ( .A(n_217), .B(n_168), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_214), .A2(n_189), .B(n_160), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_214), .A2(n_160), .B(n_184), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_198), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_225), .A2(n_165), .B(n_184), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_220), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_225), .A2(n_226), .B(n_206), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_229), .A2(n_194), .B(n_190), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_201), .A2(n_184), .B(n_165), .C(n_166), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_203), .B(n_176), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_227), .A2(n_165), .A3(n_166), .B(n_174), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_230), .A2(n_166), .B(n_176), .C(n_42), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_209), .B(n_174), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_213), .B(n_174), .Y(n_252) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_152), .B(n_149), .Y(n_253) );
AO32x2_ASAP7_75t_L g254 ( .A1(n_228), .A2(n_13), .A3(n_14), .B1(n_16), .B2(n_17), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_197), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_211), .A2(n_180), .B(n_167), .C(n_196), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_196), .B(n_180), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_221), .A2(n_196), .B(n_180), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_208), .B(n_13), .Y(n_260) );
OAI22x1_ASAP7_75t_L g261 ( .A1(n_212), .A2(n_14), .B1(n_17), .B2(n_18), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_253), .A2(n_218), .B(n_219), .Y(n_262) );
CKINVDCx8_ASAP7_75t_R g263 ( .A(n_236), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_238), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_240), .A2(n_207), .B(n_199), .C(n_204), .Y(n_265) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_230), .B(n_231), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_260), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_239), .A2(n_233), .B(n_211), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_244), .B(n_202), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_222), .A3(n_215), .B(n_223), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_259), .A2(n_222), .B(n_215), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_246), .Y(n_274) );
OAI21x1_ASAP7_75t_SL g275 ( .A1(n_237), .A2(n_210), .B(n_197), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_250), .Y(n_276) );
OR2x6_ASAP7_75t_L g277 ( .A(n_251), .B(n_167), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_243), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_249), .A2(n_196), .B(n_152), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_252), .A2(n_19), .B1(n_152), .B2(n_21), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_245), .A2(n_19), .B(n_20), .C(n_22), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_250), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_257), .B(n_65), .Y(n_283) );
AOI21x1_ASAP7_75t_L g284 ( .A1(n_234), .A2(n_33), .B(n_34), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_249), .A2(n_35), .B(n_36), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
INVx8_ASAP7_75t_L g287 ( .A(n_277), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_274), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_275), .B(n_250), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_273), .A2(n_235), .B(n_242), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_274), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_278), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_282), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_275), .B(n_250), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_267), .B(n_248), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_285), .A2(n_256), .B(n_258), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_279), .A2(n_256), .B(n_247), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_266), .B(n_248), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_266), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_248), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_303), .B(n_277), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_254), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_292), .B(n_248), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_309), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_287), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_309), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_307), .B(n_254), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_254), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_288), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_296), .B(n_265), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_254), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_294), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_296), .B(n_272), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_307), .B(n_269), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_293), .B(n_272), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_290), .Y(n_337) );
NOR2xp67_ASAP7_75t_L g338 ( .A(n_308), .B(n_284), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_290), .B(n_284), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_293), .B(n_272), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_316), .B(n_302), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_335), .B(n_301), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_319), .B(n_308), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_333), .B(n_308), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_333), .B(n_308), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_335), .B(n_298), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_321), .B(n_308), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_311), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_311), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_335), .B(n_298), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_340), .B(n_298), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_340), .B(n_299), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_314), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_340), .B(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_318), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_330), .B(n_300), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_341), .B(n_299), .Y(n_365) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_330), .B(n_290), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_341), .B(n_301), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_341), .B(n_297), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_318), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_321), .B(n_287), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_323), .B(n_297), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_321), .B(n_287), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_339), .B(n_290), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_313), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_324), .B(n_287), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_315), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_326), .B(n_291), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_326), .B(n_291), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_329), .B(n_291), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_336), .B(n_291), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_388), .B(n_329), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_388), .B(n_329), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_381), .B(n_268), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_359), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_382), .A2(n_261), .B1(n_312), .B2(n_324), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_380), .B(n_322), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_352), .B(n_342), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_386), .B(n_337), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_386), .B(n_337), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_359), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_375), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_383), .B(n_312), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_354), .B(n_312), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_387), .B(n_342), .Y(n_404) );
NOR2x1_ASAP7_75t_L g405 ( .A(n_366), .B(n_305), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_387), .B(n_385), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_361), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_336), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_346), .Y(n_409) );
NAND2xp33_ASAP7_75t_L g410 ( .A(n_354), .B(n_287), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_344), .B(n_328), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_353), .A2(n_303), .B(n_281), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_349), .B(n_318), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_384), .B(n_322), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_384), .B(n_328), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_364), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_345), .B(n_317), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_350), .B(n_334), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_363), .A2(n_287), .B1(n_303), .B2(n_313), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_355), .B(n_320), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_362), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_367), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_346), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_369), .B(n_339), .C(n_338), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_367), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_344), .B(n_334), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_356), .B(n_320), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_356), .B(n_334), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_372), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_357), .B(n_339), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_357), .B(n_291), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_343), .B(n_319), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_366), .B(n_286), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_351), .B(n_319), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_389), .B(n_306), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_389), .B(n_306), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_379), .B(n_290), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_358), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_395), .A2(n_363), .B(n_370), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_410), .A2(n_303), .B(n_379), .C(n_286), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_409), .B(n_303), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_409), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_401), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_406), .B(n_374), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_428), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_404), .B(n_378), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_390), .B(n_374), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_404), .B(n_368), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_390), .B(n_347), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_416), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_443), .B(n_425), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_391), .B(n_348), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_417), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_408), .B(n_368), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_425), .Y(n_464) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_403), .B(n_286), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_391), .B(n_376), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_444), .Y(n_467) );
HB1xp67_ASAP7_75t_SL g468 ( .A(n_402), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_397), .B(n_373), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_443), .B(n_363), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_398), .B(n_370), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_408), .B(n_365), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_398), .B(n_370), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_414), .B(n_365), .Y(n_479) );
NOR2xp67_ASAP7_75t_SL g480 ( .A(n_403), .B(n_286), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_396), .B(n_360), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_399), .B(n_360), .Y(n_482) );
OR2x6_ASAP7_75t_L g483 ( .A(n_443), .B(n_290), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_434), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_411), .B(n_371), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_393), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_300), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_415), .B(n_306), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_442), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
OAI32xp33_ASAP7_75t_L g491 ( .A1(n_467), .A2(n_392), .A3(n_436), .B1(n_426), .B2(n_439), .Y(n_491) );
NOR4xp25_ASAP7_75t_SL g492 ( .A(n_445), .B(n_410), .C(n_405), .D(n_437), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_446), .A2(n_438), .B(n_420), .Y(n_493) );
AOI32xp33_ASAP7_75t_L g494 ( .A1(n_465), .A2(n_421), .A3(n_430), .B1(n_429), .B2(n_413), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_449), .A2(n_440), .B(n_439), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_454), .A2(n_419), .B1(n_412), .B2(n_435), .C(n_430), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_473), .B(n_440), .Y(n_499) );
AOI211xp5_ASAP7_75t_L g500 ( .A1(n_480), .A2(n_305), .B(n_338), .C(n_422), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_451), .B(n_432), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_460), .A2(n_305), .B1(n_300), .B2(n_423), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_448), .B(n_441), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_462), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_472), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_463), .B(n_306), .Y(n_509) );
OAI221xp5_ASAP7_75t_SL g510 ( .A1(n_483), .A2(n_464), .B1(n_469), .B2(n_455), .C(n_487), .Y(n_510) );
OAI32xp33_ASAP7_75t_L g511 ( .A1(n_463), .A2(n_280), .A3(n_300), .B1(n_283), .B2(n_251), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_470), .A2(n_269), .B(n_236), .C(n_262), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_474), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
NOR4xp25_ASAP7_75t_SL g515 ( .A(n_510), .B(n_489), .C(n_478), .D(n_484), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_497), .A2(n_483), .B1(n_470), .B2(n_488), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_491), .B(n_479), .C(n_481), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_494), .A2(n_447), .B1(n_485), .B2(n_479), .C(n_466), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_496), .A2(n_481), .B1(n_456), .B2(n_471), .C(n_476), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_501), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_490), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_500), .A2(n_482), .B(n_452), .C(n_475), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_498), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_502), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_495), .A2(n_461), .B1(n_458), .B2(n_486), .C(n_304), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_499), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_504), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_505), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_500), .A2(n_54), .B1(n_55), .B2(n_57), .C(n_58), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_506), .A2(n_60), .B1(n_62), .B2(n_64), .C(n_514), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_507), .A2(n_513), .B1(n_508), .B2(n_509), .C(n_493), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_492), .B(n_503), .Y(n_532) );
AOI211xp5_ASAP7_75t_SL g533 ( .A1(n_512), .A2(n_497), .B(n_510), .C(n_445), .Y(n_533) );
AOI211xp5_ASAP7_75t_SL g534 ( .A1(n_511), .A2(n_497), .B(n_510), .C(n_445), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_497), .A2(n_492), .B(n_445), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_528), .B(n_535), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_527), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_523), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_529), .B(n_532), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_518), .B1(n_516), .B2(n_519), .Y(n_540) );
AND4x2_ASAP7_75t_L g541 ( .A(n_525), .B(n_534), .C(n_531), .D(n_533), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_539), .B(n_528), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_537), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_540), .B(n_516), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_544), .B(n_536), .Y(n_545) );
NOR2x1p5_ASAP7_75t_L g546 ( .A(n_543), .B(n_541), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_546), .B(n_542), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_545), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_548), .A2(n_538), .B(n_517), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_549), .B(n_547), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_550), .A2(n_547), .B1(n_515), .B2(n_526), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_551), .B(n_524), .Y(n_552) );
OR2x6_ASAP7_75t_L g553 ( .A(n_552), .B(n_520), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_553), .A2(n_521), .B1(n_522), .B2(n_530), .Y(n_554) );
endmodule