module real_jpeg_9897_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_312, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_312;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_2),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_2),
.A2(n_38),
.B1(n_60),
.B2(n_61),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_46),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_46),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_83),
.B1(n_86),
.B2(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_32),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_3),
.B(n_32),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_3),
.A2(n_29),
.B(n_33),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_3),
.A2(n_27),
.B1(n_35),
.B2(n_165),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_93),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_93),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_93),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_11),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_127),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_127),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_12),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_154),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_27),
.B1(n_35),
.B2(n_51),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_14),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_16),
.A2(n_60),
.B1(n_61),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_16),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_145),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_145),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_17),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_17),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_94),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.C(n_79),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_23),
.A2(n_66),
.B1(n_67),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_23),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_24),
.A2(n_25),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_54),
.C(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_26),
.A2(n_31),
.B1(n_37),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_26),
.A2(n_31),
.B1(n_92),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_31),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_26),
.A2(n_31),
.B1(n_126),
.B2(n_261),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_27),
.A2(n_28),
.B(n_165),
.C(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_31),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_45),
.B1(n_52),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_42),
.A2(n_45),
.B1(n_71),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_42),
.A2(n_45),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_42),
.A2(n_45),
.B1(n_190),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_42),
.A2(n_45),
.B1(n_206),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_42),
.A2(n_45),
.B1(n_245),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_42),
.A2(n_45),
.B1(n_130),
.B2(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_45),
.B(n_165),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_46),
.B(n_48),
.Y(n_194)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_47),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_55),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_59),
.B1(n_75),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_56),
.A2(n_59),
.B1(n_89),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_56),
.A2(n_59),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_56),
.A2(n_59),
.B1(n_153),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_56),
.A2(n_59),
.B1(n_178),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_56),
.A2(n_59),
.B1(n_186),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_56),
.A2(n_59),
.B1(n_123),
.B2(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_59),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_60),
.B(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_60),
.B(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_61),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_68),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_76),
.A2(n_78),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_81),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_292),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_83),
.A2(n_86),
.B1(n_144),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_83),
.A2(n_86),
.B1(n_147),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_83),
.A2(n_86),
.B1(n_180),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_83),
.A2(n_86),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_83),
.A2(n_86),
.B1(n_121),
.B2(n_233),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_84),
.A2(n_85),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_84),
.A2(n_85),
.B1(n_198),
.B2(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_86),
.B(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_134),
.B(n_310),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_131),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_110),
.B(n_131),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_111),
.Y(n_297)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_117),
.A2(n_118),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_128),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_119),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_120),
.B(n_122),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_286),
.A3(n_298),
.B1(n_304),
.B2(n_309),
.C(n_312),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_251),
.C(n_282),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_222),
.B(n_250),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_200),
.B(n_221),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_182),
.B(n_199),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_172),
.B(n_181),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_160),
.B(n_171),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_159),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_170),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_174),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.CI(n_191),
.CON(n_184),
.SN(n_184)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_196),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_214),
.B2(n_215),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_217),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_213),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_205),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_211),
.C(n_213),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_224),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_237),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_226),
.B(n_236),
.C(n_237),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_231),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_242),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_269),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_253),
.B(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.C(n_268),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_263),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_268),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_280),
.B2(n_281),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_273),
.C(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_276),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_287),
.B(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.C(n_293),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);


endmodule