module fake_jpeg_29699_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_3),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_72),
.Y(n_76)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_64),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_56),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_66),
.B(n_46),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_58),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_57),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_65),
.B1(n_50),
.B2(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_50),
.B1(n_48),
.B2(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_98),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_52),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_63),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_55),
.B1(n_61),
.B2(n_59),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_58),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_41),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_108),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_62),
.B1(n_53),
.B2(n_51),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_1),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_122),
.B1(n_128),
.B2(n_18),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_100),
.B1(n_108),
.B2(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_124),
.B1(n_21),
.B2(n_22),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_8),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_9),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_13),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_139),
.B1(n_120),
.B2(n_121),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_141),
.Y(n_148)
);

XNOR2x2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_20),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_142),
.B(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_152),
.B1(n_132),
.B2(n_145),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_111),
.B(n_118),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_151),
.A2(n_132),
.B(n_144),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_136),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_156),
.C(n_149),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_148),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_155),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_157),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_150),
.B(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_131),
.Y(n_164)
);


endmodule